magic
tech sky130A
magscale 1 2
timestamp 1626450099
<< checkpaint >>
rect -1260 -1260 13444 11004
<< viali >>
rect 8145 6385 8179 6419
rect 3545 6181 3579 6215
rect 4189 6181 4223 6215
rect 7961 6181 7995 6215
rect 3729 6045 3763 6079
rect 6673 5705 6707 5739
rect 8053 5705 8087 5739
rect 6949 5637 6983 5671
rect 6765 5569 6799 5603
rect 7869 5569 7903 5603
rect 6857 5501 6891 5535
rect 7593 5297 7627 5331
rect 3545 5093 3579 5127
rect 4189 5093 4223 5127
rect 6397 5093 6431 5127
rect 6489 5093 6523 5127
rect 6627 5093 6661 5127
rect 6765 5093 6799 5127
rect 6857 5093 6891 5127
rect 7409 5093 7443 5127
rect 7501 5093 7535 5127
rect 7685 5025 7719 5059
rect 8237 5025 8271 5059
rect 3729 4957 3763 4991
rect 5477 4957 5511 4991
rect 6581 4957 6615 4991
rect 5707 4753 5741 4787
rect 7501 4685 7535 4719
rect 5604 4617 5638 4651
rect 6213 4617 6247 4651
rect 6397 4617 6431 4651
rect 6489 4617 6523 4651
rect 6765 4617 6799 4651
rect 7225 4617 7259 4651
rect 7317 4617 7351 4651
rect 7593 4617 7627 4651
rect 7685 4617 7719 4651
rect 6673 4481 6707 4515
rect 7225 4481 7259 4515
rect 5109 4413 5143 4447
rect 6581 4413 6615 4447
rect 6857 4209 6891 4243
rect 7547 4209 7581 4243
rect 6765 4141 6799 4175
rect 6397 4005 6431 4039
rect 6581 4005 6615 4039
rect 6673 4005 6707 4039
rect 6949 4005 6983 4039
rect 7444 4005 7478 4039
rect 5385 3869 5419 3903
rect 6627 3665 6661 3699
rect 7961 3665 7995 3699
rect 6524 3529 6558 3563
rect 7501 3529 7535 3563
rect 8145 3529 8179 3563
<< metal1 >>
rect 3240 6530 8944 6552
rect 3240 6478 4019 6530
rect 4071 6478 4083 6530
rect 4135 6478 4147 6530
rect 4199 6478 4211 6530
rect 4263 6478 4275 6530
rect 4327 6478 4339 6530
rect 4391 6478 5950 6530
rect 6002 6478 6014 6530
rect 6066 6478 6078 6530
rect 6130 6478 6142 6530
rect 6194 6478 6206 6530
rect 6258 6478 6270 6530
rect 6322 6478 7880 6530
rect 7932 6478 7944 6530
rect 7996 6478 8008 6530
rect 8060 6478 8072 6530
rect 8124 6478 8136 6530
rect 8188 6478 8200 6530
rect 8252 6478 8944 6530
rect 3240 6456 8944 6478
rect 8133 6419 8191 6425
rect 8133 6385 8145 6419
rect 8179 6416 8191 6419
rect 9142 6416 9148 6428
rect 8179 6388 9148 6416
rect 8179 6385 8191 6388
rect 8133 6379 8191 6385
rect 9142 6376 9148 6388
rect 9200 6376 9206 6428
rect 3162 6172 3168 6224
rect 3220 6212 3226 6224
rect 3533 6215 3591 6221
rect 3533 6212 3545 6215
rect 3220 6184 3545 6212
rect 3220 6172 3226 6184
rect 3533 6181 3545 6184
rect 3579 6212 3591 6215
rect 4177 6215 4235 6221
rect 4177 6212 4189 6215
rect 3579 6184 4189 6212
rect 3579 6181 3591 6184
rect 3533 6175 3591 6181
rect 4177 6181 4189 6184
rect 4223 6181 4235 6215
rect 4177 6175 4235 6181
rect 7578 6172 7584 6224
rect 7636 6212 7642 6224
rect 7949 6215 8007 6221
rect 7949 6212 7961 6215
rect 7636 6184 7961 6212
rect 7636 6172 7642 6184
rect 7949 6181 7961 6184
rect 7995 6181 8007 6215
rect 7949 6175 8007 6181
rect 3717 6079 3775 6085
rect 3717 6045 3729 6079
rect 3763 6076 3775 6079
rect 6658 6076 6664 6088
rect 3763 6048 6664 6076
rect 3763 6045 3775 6048
rect 3717 6039 3775 6045
rect 6658 6036 6664 6048
rect 6716 6036 6722 6088
rect 3240 5986 8944 6008
rect 3240 5934 4984 5986
rect 5036 5934 5048 5986
rect 5100 5934 5112 5986
rect 5164 5934 5176 5986
rect 5228 5934 5240 5986
rect 5292 5934 5304 5986
rect 5356 5934 6915 5986
rect 6967 5934 6979 5986
rect 7031 5934 7043 5986
rect 7095 5934 7107 5986
rect 7159 5934 7171 5986
rect 7223 5934 7235 5986
rect 7287 5934 8944 5986
rect 3240 5912 8944 5934
rect 6566 5696 6572 5748
rect 6624 5736 6630 5748
rect 6661 5739 6719 5745
rect 6661 5736 6673 5739
rect 6624 5708 6673 5736
rect 6624 5696 6630 5708
rect 6661 5705 6673 5708
rect 6707 5705 6719 5739
rect 6661 5699 6719 5705
rect 8041 5739 8099 5745
rect 8041 5705 8053 5739
rect 8087 5736 8099 5739
rect 8314 5736 8320 5748
rect 8087 5708 8320 5736
rect 8087 5705 8099 5708
rect 8041 5699 8099 5705
rect 8314 5696 8320 5708
rect 8372 5696 8378 5748
rect 6937 5671 6995 5677
rect 6937 5637 6949 5671
rect 6983 5668 6995 5671
rect 7578 5668 7584 5680
rect 6983 5640 7584 5668
rect 6983 5637 6995 5640
rect 6937 5631 6995 5637
rect 7578 5628 7584 5640
rect 7636 5628 7642 5680
rect 6750 5600 6756 5612
rect 6711 5572 6756 5600
rect 6750 5560 6756 5572
rect 6808 5560 6814 5612
rect 7026 5560 7032 5612
rect 7084 5600 7090 5612
rect 7857 5603 7915 5609
rect 7857 5600 7869 5603
rect 7084 5572 7869 5600
rect 7084 5560 7090 5572
rect 7857 5569 7869 5572
rect 7903 5569 7915 5603
rect 7857 5563 7915 5569
rect 6845 5535 6903 5541
rect 6845 5501 6857 5535
rect 6891 5532 6903 5535
rect 7394 5532 7400 5544
rect 6891 5504 7400 5532
rect 6891 5501 6903 5504
rect 6845 5495 6903 5501
rect 7394 5492 7400 5504
rect 7452 5492 7458 5544
rect 3240 5442 8944 5464
rect 3240 5390 4019 5442
rect 4071 5390 4083 5442
rect 4135 5390 4147 5442
rect 4199 5390 4211 5442
rect 4263 5390 4275 5442
rect 4327 5390 4339 5442
rect 4391 5390 5950 5442
rect 6002 5390 6014 5442
rect 6066 5390 6078 5442
rect 6130 5390 6142 5442
rect 6194 5390 6206 5442
rect 6258 5390 6270 5442
rect 6322 5390 7880 5442
rect 7932 5390 7944 5442
rect 7996 5390 8008 5442
rect 8060 5390 8072 5442
rect 8124 5390 8136 5442
rect 8188 5390 8200 5442
rect 8252 5390 8944 5442
rect 3240 5368 8944 5390
rect 7578 5328 7584 5340
rect 6400 5300 6796 5328
rect 7539 5300 7584 5328
rect 3162 5084 3168 5136
rect 3220 5124 3226 5136
rect 6400 5133 6428 5300
rect 6658 5260 6664 5272
rect 6492 5232 6664 5260
rect 6492 5133 6520 5232
rect 6658 5220 6664 5232
rect 6716 5220 6722 5272
rect 6768 5192 6796 5300
rect 7578 5288 7584 5300
rect 7636 5288 7642 5340
rect 6768 5164 7532 5192
rect 7504 5136 7532 5164
rect 3533 5127 3591 5133
rect 3533 5124 3545 5127
rect 3220 5096 3545 5124
rect 3220 5084 3226 5096
rect 3533 5093 3545 5096
rect 3579 5124 3591 5127
rect 4177 5127 4235 5133
rect 4177 5124 4189 5127
rect 3579 5096 4189 5124
rect 3579 5093 3591 5096
rect 3533 5087 3591 5093
rect 4177 5093 4189 5096
rect 4223 5093 4235 5127
rect 4177 5087 4235 5093
rect 6385 5127 6443 5133
rect 6385 5093 6397 5127
rect 6431 5093 6443 5127
rect 6385 5087 6443 5093
rect 6477 5127 6535 5133
rect 6477 5093 6489 5127
rect 6523 5093 6535 5127
rect 6477 5087 6535 5093
rect 6615 5127 6673 5133
rect 6615 5093 6627 5127
rect 6661 5093 6673 5127
rect 6615 5087 6673 5093
rect 6753 5127 6811 5133
rect 6753 5093 6765 5127
rect 6799 5124 6811 5127
rect 6845 5127 6903 5133
rect 6845 5124 6857 5127
rect 6799 5096 6857 5124
rect 6799 5093 6811 5096
rect 6753 5087 6811 5093
rect 6845 5093 6857 5096
rect 6891 5124 6903 5127
rect 7026 5124 7032 5136
rect 6891 5096 7032 5124
rect 6891 5093 6903 5096
rect 6845 5087 6903 5093
rect 6630 5056 6658 5087
rect 7026 5084 7032 5096
rect 7084 5084 7090 5136
rect 7394 5124 7400 5136
rect 7355 5096 7400 5124
rect 7394 5084 7400 5096
rect 7452 5084 7458 5136
rect 7486 5084 7492 5136
rect 7544 5124 7550 5136
rect 7544 5096 7589 5124
rect 7544 5084 7550 5096
rect 6400 5028 6658 5056
rect 7044 5056 7072 5084
rect 7302 5056 7308 5068
rect 7044 5028 7308 5056
rect 6400 5000 6428 5028
rect 7302 5016 7308 5028
rect 7360 5016 7366 5068
rect 7670 5056 7676 5068
rect 7631 5028 7676 5056
rect 7670 5016 7676 5028
rect 7728 5016 7734 5068
rect 8225 5059 8283 5065
rect 8225 5025 8237 5059
rect 8271 5056 8283 5059
rect 8314 5056 8320 5068
rect 8271 5028 8320 5056
rect 8271 5025 8283 5028
rect 8225 5019 8283 5025
rect 8314 5016 8320 5028
rect 8372 5056 8378 5068
rect 9142 5056 9148 5068
rect 8372 5028 9148 5056
rect 8372 5016 8378 5028
rect 9142 5016 9148 5028
rect 9200 5016 9206 5068
rect 3714 4988 3720 5000
rect 3675 4960 3720 4988
rect 3714 4948 3720 4960
rect 3772 4948 3778 5000
rect 5462 4988 5468 5000
rect 5423 4960 5468 4988
rect 5462 4948 5468 4960
rect 5520 4948 5526 5000
rect 6382 4948 6388 5000
rect 6440 4948 6446 5000
rect 6566 4988 6572 5000
rect 6527 4960 6572 4988
rect 6566 4948 6572 4960
rect 6624 4948 6630 5000
rect 6658 4948 6664 5000
rect 6716 4988 6722 5000
rect 7394 4988 7400 5000
rect 6716 4960 7400 4988
rect 6716 4948 6722 4960
rect 7394 4948 7400 4960
rect 7452 4948 7458 5000
rect 3240 4898 8944 4920
rect 3240 4846 4984 4898
rect 5036 4846 5048 4898
rect 5100 4846 5112 4898
rect 5164 4846 5176 4898
rect 5228 4846 5240 4898
rect 5292 4846 5304 4898
rect 5356 4846 6915 4898
rect 6967 4846 6979 4898
rect 7031 4846 7043 4898
rect 7095 4846 7107 4898
rect 7159 4846 7171 4898
rect 7223 4846 7235 4898
rect 7287 4846 8944 4898
rect 3240 4824 8944 4846
rect 5695 4787 5753 4793
rect 5695 4753 5707 4787
rect 5741 4784 5753 4787
rect 6382 4784 6388 4796
rect 5741 4756 6388 4784
rect 5741 4753 5753 4756
rect 5695 4747 5753 4753
rect 6382 4744 6388 4756
rect 6440 4784 6446 4796
rect 6440 4756 7532 4784
rect 6440 4744 6446 4756
rect 3714 4676 3720 4728
rect 3772 4716 3778 4728
rect 3772 4688 6520 4716
rect 3772 4676 3778 4688
rect 5462 4648 5468 4660
rect 5112 4620 5468 4648
rect 5112 4456 5140 4620
rect 5462 4608 5468 4620
rect 5520 4648 5526 4660
rect 5592 4651 5650 4657
rect 5592 4648 5604 4651
rect 5520 4620 5604 4648
rect 5520 4608 5526 4620
rect 5592 4617 5604 4620
rect 5638 4648 5650 4651
rect 6201 4651 6259 4657
rect 5638 4620 6152 4648
rect 5638 4617 5650 4620
rect 5592 4611 5650 4617
rect 6124 4580 6152 4620
rect 6201 4617 6213 4651
rect 6247 4648 6259 4651
rect 6290 4648 6296 4660
rect 6247 4620 6296 4648
rect 6247 4617 6259 4620
rect 6201 4611 6259 4617
rect 6290 4608 6296 4620
rect 6348 4608 6354 4660
rect 6492 4657 6520 4688
rect 6566 4676 6572 4728
rect 6624 4716 6630 4728
rect 7504 4725 7532 4756
rect 7489 4719 7547 4725
rect 6624 4688 7256 4716
rect 6624 4676 6630 4688
rect 6385 4651 6443 4657
rect 6385 4617 6397 4651
rect 6431 4617 6443 4651
rect 6385 4611 6443 4617
rect 6477 4651 6535 4657
rect 6477 4617 6489 4651
rect 6523 4648 6535 4651
rect 6658 4648 6664 4660
rect 6523 4620 6664 4648
rect 6523 4617 6535 4620
rect 6477 4611 6535 4617
rect 6400 4580 6428 4611
rect 6658 4608 6664 4620
rect 6716 4608 6722 4660
rect 7228 4657 7256 4688
rect 7489 4685 7501 4719
rect 7535 4685 7547 4719
rect 7489 4679 7547 4685
rect 6753 4651 6811 4657
rect 6753 4617 6765 4651
rect 6799 4617 6811 4651
rect 6753 4611 6811 4617
rect 7213 4651 7271 4657
rect 7213 4617 7225 4651
rect 7259 4617 7271 4651
rect 7213 4611 7271 4617
rect 7305 4651 7363 4657
rect 7305 4617 7317 4651
rect 7351 4648 7363 4651
rect 7394 4648 7400 4660
rect 7351 4620 7400 4648
rect 7351 4617 7363 4620
rect 7305 4611 7363 4617
rect 6124 4552 6428 4580
rect 6768 4580 6796 4611
rect 7394 4608 7400 4620
rect 7452 4608 7458 4660
rect 7581 4651 7639 4657
rect 7581 4617 7593 4651
rect 7627 4648 7639 4651
rect 7673 4651 7731 4657
rect 7673 4648 7685 4651
rect 7627 4620 7685 4648
rect 7627 4617 7639 4620
rect 7581 4611 7639 4617
rect 7673 4617 7685 4620
rect 7719 4648 7731 4651
rect 7762 4648 7768 4660
rect 7719 4620 7768 4648
rect 7719 4617 7731 4620
rect 7673 4611 7731 4617
rect 7596 4580 7624 4611
rect 7762 4608 7768 4620
rect 7820 4608 7826 4660
rect 6768 4552 7624 4580
rect 6661 4515 6719 4521
rect 6661 4481 6673 4515
rect 6707 4512 6719 4515
rect 6768 4512 6796 4552
rect 6707 4484 6796 4512
rect 7213 4515 7271 4521
rect 6707 4481 6719 4484
rect 6661 4475 6719 4481
rect 7213 4481 7225 4515
rect 7259 4512 7271 4515
rect 7486 4512 7492 4524
rect 7259 4484 7492 4512
rect 7259 4481 7271 4484
rect 7213 4475 7271 4481
rect 7486 4472 7492 4484
rect 7544 4472 7550 4524
rect 5094 4444 5100 4456
rect 5055 4416 5100 4444
rect 5094 4404 5100 4416
rect 5152 4404 5158 4456
rect 6382 4404 6388 4456
rect 6440 4444 6446 4456
rect 6569 4447 6627 4453
rect 6569 4444 6581 4447
rect 6440 4416 6581 4444
rect 6440 4404 6446 4416
rect 6569 4413 6581 4416
rect 6615 4413 6627 4447
rect 6569 4407 6627 4413
rect 3240 4354 8944 4376
rect 3240 4302 4019 4354
rect 4071 4302 4083 4354
rect 4135 4302 4147 4354
rect 4199 4302 4211 4354
rect 4263 4302 4275 4354
rect 4327 4302 4339 4354
rect 4391 4302 5950 4354
rect 6002 4302 6014 4354
rect 6066 4302 6078 4354
rect 6130 4302 6142 4354
rect 6194 4302 6206 4354
rect 6258 4302 6270 4354
rect 6322 4302 7880 4354
rect 7932 4302 7944 4354
rect 7996 4302 8008 4354
rect 8060 4302 8072 4354
rect 8124 4302 8136 4354
rect 8188 4302 8200 4354
rect 8252 4302 8944 4354
rect 3240 4280 8944 4302
rect 6845 4243 6903 4249
rect 6845 4209 6857 4243
rect 6891 4240 6903 4243
rect 6934 4240 6940 4252
rect 6891 4212 6940 4240
rect 6891 4209 6903 4212
rect 6845 4203 6903 4209
rect 6934 4200 6940 4212
rect 6992 4240 6998 4252
rect 7302 4240 7308 4252
rect 6992 4212 7308 4240
rect 6992 4200 6998 4212
rect 7302 4200 7308 4212
rect 7360 4200 7366 4252
rect 7535 4243 7593 4249
rect 7535 4209 7547 4243
rect 7581 4240 7593 4243
rect 7670 4240 7676 4252
rect 7581 4212 7676 4240
rect 7581 4209 7593 4212
rect 7535 4203 7593 4209
rect 7670 4200 7676 4212
rect 7728 4200 7734 4252
rect 6474 4132 6480 4184
rect 6532 4172 6538 4184
rect 6753 4175 6811 4181
rect 6753 4172 6765 4175
rect 6532 4144 6765 4172
rect 6532 4132 6538 4144
rect 6753 4141 6765 4144
rect 6799 4172 6811 4175
rect 6799 4144 7072 4172
rect 6799 4141 6811 4144
rect 6753 4135 6811 4141
rect 6382 4036 6388 4048
rect 6343 4008 6388 4036
rect 6382 3996 6388 4008
rect 6440 3996 6446 4048
rect 6569 4039 6627 4045
rect 6569 4005 6581 4039
rect 6615 4005 6627 4039
rect 6569 3999 6627 4005
rect 5094 3928 5100 3980
rect 5152 3928 5158 3980
rect 6584 3968 6612 3999
rect 6658 3996 6664 4048
rect 6716 4036 6722 4048
rect 6934 4036 6940 4048
rect 6716 4008 6761 4036
rect 6895 4008 6940 4036
rect 6716 3996 6722 4008
rect 6934 3996 6940 4008
rect 6992 3996 6998 4048
rect 7044 4036 7072 4144
rect 7432 4039 7490 4045
rect 7432 4036 7444 4039
rect 7044 4008 7444 4036
rect 7432 4005 7444 4008
rect 7478 4005 7490 4039
rect 7432 3999 7490 4005
rect 5388 3940 6612 3968
rect 3162 3860 3168 3912
rect 3220 3900 3226 3912
rect 5112 3900 5140 3928
rect 5388 3909 5416 3940
rect 5373 3903 5431 3909
rect 5373 3900 5385 3903
rect 3220 3872 5385 3900
rect 3220 3860 3226 3872
rect 5373 3869 5385 3872
rect 5419 3869 5431 3903
rect 5373 3863 5431 3869
rect 3240 3810 8944 3832
rect 3240 3758 4984 3810
rect 5036 3758 5048 3810
rect 5100 3758 5112 3810
rect 5164 3758 5176 3810
rect 5228 3758 5240 3810
rect 5292 3758 5304 3810
rect 5356 3758 6915 3810
rect 6967 3758 6979 3810
rect 7031 3758 7043 3810
rect 7095 3758 7107 3810
rect 7159 3758 7171 3810
rect 7223 3758 7235 3810
rect 7287 3758 8944 3810
rect 3240 3736 8944 3758
rect 6615 3699 6673 3705
rect 6615 3665 6627 3699
rect 6661 3696 6673 3699
rect 6750 3696 6756 3708
rect 6661 3668 6756 3696
rect 6661 3665 6673 3668
rect 6615 3659 6673 3665
rect 6750 3656 6756 3668
rect 6808 3656 6814 3708
rect 7762 3656 7768 3708
rect 7820 3696 7826 3708
rect 7949 3699 8007 3705
rect 7949 3696 7961 3699
rect 7820 3668 7961 3696
rect 7820 3656 7826 3668
rect 7949 3665 7961 3668
rect 7995 3665 8007 3699
rect 7949 3659 8007 3665
rect 6382 3520 6388 3572
rect 6440 3560 6446 3572
rect 6512 3563 6570 3569
rect 6512 3560 6524 3563
rect 6440 3532 6524 3560
rect 6440 3520 6446 3532
rect 6512 3529 6524 3532
rect 6558 3529 6570 3563
rect 6512 3523 6570 3529
rect 7489 3563 7547 3569
rect 7489 3529 7501 3563
rect 7535 3560 7547 3563
rect 8133 3563 8191 3569
rect 8133 3560 8145 3563
rect 7535 3532 8145 3560
rect 7535 3529 7547 3532
rect 7489 3523 7547 3529
rect 8133 3529 8145 3532
rect 8179 3560 8191 3563
rect 9142 3560 9148 3572
rect 8179 3532 9148 3560
rect 8179 3529 8191 3532
rect 8133 3523 8191 3529
rect 9142 3520 9148 3532
rect 9200 3520 9206 3572
rect 3240 3266 8944 3288
rect 3240 3214 4019 3266
rect 4071 3214 4083 3266
rect 4135 3214 4147 3266
rect 4199 3214 4211 3266
rect 4263 3214 4275 3266
rect 4327 3214 4339 3266
rect 4391 3214 5950 3266
rect 6002 3214 6014 3266
rect 6066 3214 6078 3266
rect 6130 3214 6142 3266
rect 6194 3214 6206 3266
rect 6258 3214 6270 3266
rect 6322 3214 7880 3266
rect 7932 3214 7944 3266
rect 7996 3214 8008 3266
rect 8060 3214 8072 3266
rect 8124 3214 8136 3266
rect 8188 3214 8200 3266
rect 8252 3214 8944 3266
rect 3240 3192 8944 3214
<< via1 >>
rect 4019 6478 4071 6530
rect 4083 6478 4135 6530
rect 4147 6478 4199 6530
rect 4211 6478 4263 6530
rect 4275 6478 4327 6530
rect 4339 6478 4391 6530
rect 5950 6478 6002 6530
rect 6014 6478 6066 6530
rect 6078 6478 6130 6530
rect 6142 6478 6194 6530
rect 6206 6478 6258 6530
rect 6270 6478 6322 6530
rect 7880 6478 7932 6530
rect 7944 6478 7996 6530
rect 8008 6478 8060 6530
rect 8072 6478 8124 6530
rect 8136 6478 8188 6530
rect 8200 6478 8252 6530
rect 9148 6376 9200 6428
rect 3168 6172 3220 6224
rect 7584 6172 7636 6224
rect 6664 6036 6716 6088
rect 4984 5934 5036 5986
rect 5048 5934 5100 5986
rect 5112 5934 5164 5986
rect 5176 5934 5228 5986
rect 5240 5934 5292 5986
rect 5304 5934 5356 5986
rect 6915 5934 6967 5986
rect 6979 5934 7031 5986
rect 7043 5934 7095 5986
rect 7107 5934 7159 5986
rect 7171 5934 7223 5986
rect 7235 5934 7287 5986
rect 6572 5696 6624 5748
rect 8320 5696 8372 5748
rect 7584 5628 7636 5680
rect 6756 5603 6808 5612
rect 6756 5569 6765 5603
rect 6765 5569 6799 5603
rect 6799 5569 6808 5603
rect 6756 5560 6808 5569
rect 7032 5560 7084 5612
rect 7400 5492 7452 5544
rect 4019 5390 4071 5442
rect 4083 5390 4135 5442
rect 4147 5390 4199 5442
rect 4211 5390 4263 5442
rect 4275 5390 4327 5442
rect 4339 5390 4391 5442
rect 5950 5390 6002 5442
rect 6014 5390 6066 5442
rect 6078 5390 6130 5442
rect 6142 5390 6194 5442
rect 6206 5390 6258 5442
rect 6270 5390 6322 5442
rect 7880 5390 7932 5442
rect 7944 5390 7996 5442
rect 8008 5390 8060 5442
rect 8072 5390 8124 5442
rect 8136 5390 8188 5442
rect 8200 5390 8252 5442
rect 7584 5331 7636 5340
rect 3168 5084 3220 5136
rect 6664 5220 6716 5272
rect 7584 5297 7593 5331
rect 7593 5297 7627 5331
rect 7627 5297 7636 5331
rect 7584 5288 7636 5297
rect 7032 5084 7084 5136
rect 7400 5127 7452 5136
rect 7400 5093 7409 5127
rect 7409 5093 7443 5127
rect 7443 5093 7452 5127
rect 7400 5084 7452 5093
rect 7492 5127 7544 5136
rect 7492 5093 7501 5127
rect 7501 5093 7535 5127
rect 7535 5093 7544 5127
rect 7492 5084 7544 5093
rect 7308 5016 7360 5068
rect 7676 5059 7728 5068
rect 7676 5025 7685 5059
rect 7685 5025 7719 5059
rect 7719 5025 7728 5059
rect 7676 5016 7728 5025
rect 8320 5016 8372 5068
rect 9148 5016 9200 5068
rect 3720 4991 3772 5000
rect 3720 4957 3729 4991
rect 3729 4957 3763 4991
rect 3763 4957 3772 4991
rect 3720 4948 3772 4957
rect 5468 4991 5520 5000
rect 5468 4957 5477 4991
rect 5477 4957 5511 4991
rect 5511 4957 5520 4991
rect 5468 4948 5520 4957
rect 6388 4948 6440 5000
rect 6572 4991 6624 5000
rect 6572 4957 6581 4991
rect 6581 4957 6615 4991
rect 6615 4957 6624 4991
rect 6572 4948 6624 4957
rect 6664 4948 6716 5000
rect 7400 4948 7452 5000
rect 4984 4846 5036 4898
rect 5048 4846 5100 4898
rect 5112 4846 5164 4898
rect 5176 4846 5228 4898
rect 5240 4846 5292 4898
rect 5304 4846 5356 4898
rect 6915 4846 6967 4898
rect 6979 4846 7031 4898
rect 7043 4846 7095 4898
rect 7107 4846 7159 4898
rect 7171 4846 7223 4898
rect 7235 4846 7287 4898
rect 6388 4744 6440 4796
rect 3720 4676 3772 4728
rect 5468 4608 5520 4660
rect 6296 4608 6348 4660
rect 6572 4676 6624 4728
rect 6664 4608 6716 4660
rect 7400 4608 7452 4660
rect 7768 4608 7820 4660
rect 7492 4472 7544 4524
rect 5100 4447 5152 4456
rect 5100 4413 5109 4447
rect 5109 4413 5143 4447
rect 5143 4413 5152 4447
rect 5100 4404 5152 4413
rect 6388 4404 6440 4456
rect 4019 4302 4071 4354
rect 4083 4302 4135 4354
rect 4147 4302 4199 4354
rect 4211 4302 4263 4354
rect 4275 4302 4327 4354
rect 4339 4302 4391 4354
rect 5950 4302 6002 4354
rect 6014 4302 6066 4354
rect 6078 4302 6130 4354
rect 6142 4302 6194 4354
rect 6206 4302 6258 4354
rect 6270 4302 6322 4354
rect 7880 4302 7932 4354
rect 7944 4302 7996 4354
rect 8008 4302 8060 4354
rect 8072 4302 8124 4354
rect 8136 4302 8188 4354
rect 8200 4302 8252 4354
rect 6940 4200 6992 4252
rect 7308 4200 7360 4252
rect 7676 4200 7728 4252
rect 6480 4132 6532 4184
rect 6388 4039 6440 4048
rect 6388 4005 6397 4039
rect 6397 4005 6431 4039
rect 6431 4005 6440 4039
rect 6388 3996 6440 4005
rect 5100 3928 5152 3980
rect 6664 4039 6716 4048
rect 6664 4005 6673 4039
rect 6673 4005 6707 4039
rect 6707 4005 6716 4039
rect 6940 4039 6992 4048
rect 6664 3996 6716 4005
rect 6940 4005 6949 4039
rect 6949 4005 6983 4039
rect 6983 4005 6992 4039
rect 6940 3996 6992 4005
rect 3168 3860 3220 3912
rect 4984 3758 5036 3810
rect 5048 3758 5100 3810
rect 5112 3758 5164 3810
rect 5176 3758 5228 3810
rect 5240 3758 5292 3810
rect 5304 3758 5356 3810
rect 6915 3758 6967 3810
rect 6979 3758 7031 3810
rect 7043 3758 7095 3810
rect 7107 3758 7159 3810
rect 7171 3758 7223 3810
rect 7235 3758 7287 3810
rect 6756 3656 6808 3708
rect 7768 3656 7820 3708
rect 6388 3520 6440 3572
rect 9148 3520 9200 3572
rect 4019 3214 4071 3266
rect 4083 3214 4135 3266
rect 4147 3214 4199 3266
rect 4211 3214 4263 3266
rect 4275 3214 4327 3266
rect 4339 3214 4391 3266
rect 5950 3214 6002 3266
rect 6014 3214 6066 3266
rect 6078 3214 6130 3266
rect 6142 3214 6194 3266
rect 6206 3214 6258 3266
rect 6270 3214 6322 3266
rect 7880 3214 7932 3266
rect 7944 3214 7996 3266
rect 8008 3214 8060 3266
rect 8072 3214 8124 3266
rect 8136 3214 8188 3266
rect 8200 3214 8252 3266
<< metal2 >>
rect 2136 7748 2936 8560
rect 9336 7748 10136 7846
rect 2136 7720 3208 7748
rect 2136 7622 2936 7720
rect 3180 6230 3208 7720
rect 9160 7720 10136 7748
rect 4017 6532 4393 6552
rect 4073 6530 4097 6532
rect 4153 6530 4177 6532
rect 4233 6530 4257 6532
rect 4313 6530 4337 6532
rect 4073 6478 4083 6530
rect 4327 6478 4337 6530
rect 4073 6476 4097 6478
rect 4153 6476 4177 6478
rect 4233 6476 4257 6478
rect 4313 6476 4337 6478
rect 4017 6456 4393 6476
rect 5948 6532 6324 6552
rect 6004 6530 6028 6532
rect 6084 6530 6108 6532
rect 6164 6530 6188 6532
rect 6244 6530 6268 6532
rect 6004 6478 6014 6530
rect 6258 6478 6268 6530
rect 6004 6476 6028 6478
rect 6084 6476 6108 6478
rect 6164 6476 6188 6478
rect 6244 6476 6268 6478
rect 5948 6456 6324 6476
rect 7878 6532 8254 6552
rect 7934 6530 7958 6532
rect 8014 6530 8038 6532
rect 8094 6530 8118 6532
rect 8174 6530 8198 6532
rect 7934 6478 7944 6530
rect 8188 6478 8198 6530
rect 7934 6476 7958 6478
rect 8014 6476 8038 6478
rect 8094 6476 8118 6478
rect 8174 6476 8198 6478
rect 7878 6456 8254 6476
rect 9160 6434 9188 7720
rect 9336 7622 10136 7720
rect 9148 6428 9200 6434
rect 9148 6370 9200 6376
rect 3168 6224 3220 6230
rect 3168 6166 3220 6172
rect 7584 6224 7636 6230
rect 7584 6166 7636 6172
rect 6664 6088 6716 6094
rect 6664 6030 6716 6036
rect 4982 5988 5358 6008
rect 5038 5986 5062 5988
rect 5118 5986 5142 5988
rect 5198 5986 5222 5988
rect 5278 5986 5302 5988
rect 5038 5934 5048 5986
rect 5292 5934 5302 5986
rect 5038 5932 5062 5934
rect 5118 5932 5142 5934
rect 5198 5932 5222 5934
rect 5278 5932 5302 5934
rect 4982 5912 5358 5932
rect 6572 5748 6624 5754
rect 6572 5690 6624 5696
rect 4017 5444 4393 5464
rect 4073 5442 4097 5444
rect 4153 5442 4177 5444
rect 4233 5442 4257 5444
rect 4313 5442 4337 5444
rect 4073 5390 4083 5442
rect 4327 5390 4337 5442
rect 4073 5388 4097 5390
rect 4153 5388 4177 5390
rect 4233 5388 4257 5390
rect 4313 5388 4337 5390
rect 4017 5368 4393 5388
rect 5948 5444 6324 5464
rect 6004 5442 6028 5444
rect 6084 5442 6108 5444
rect 6164 5442 6188 5444
rect 6244 5442 6268 5444
rect 6004 5390 6014 5442
rect 6258 5390 6268 5442
rect 6004 5388 6028 5390
rect 6084 5388 6108 5390
rect 6164 5388 6188 5390
rect 6244 5388 6268 5390
rect 5948 5368 6324 5388
rect 20 5080 2936 5178
rect 3168 5136 3220 5142
rect 3168 5080 3220 5084
rect 20 5078 3220 5080
rect 20 5052 3208 5078
rect 20 4954 2936 5052
rect 6584 5006 6612 5690
rect 6676 5278 6704 6030
rect 6913 5988 7289 6008
rect 6969 5986 6993 5988
rect 7049 5986 7073 5988
rect 7129 5986 7153 5988
rect 7209 5986 7233 5988
rect 6969 5934 6979 5986
rect 7223 5934 7233 5986
rect 6969 5932 6993 5934
rect 7049 5932 7073 5934
rect 7129 5932 7153 5934
rect 7209 5932 7233 5934
rect 6913 5912 7289 5932
rect 7596 5686 7624 6166
rect 8320 5748 8372 5754
rect 8320 5690 8372 5696
rect 7584 5680 7636 5686
rect 7584 5622 7636 5628
rect 6756 5612 6808 5618
rect 6756 5554 6808 5560
rect 7032 5612 7084 5618
rect 7032 5554 7084 5560
rect 6664 5272 6716 5278
rect 6664 5214 6716 5220
rect 6676 5006 6704 5214
rect 3720 5000 3772 5006
rect 3720 4942 3772 4948
rect 5468 5000 5520 5006
rect 5468 4942 5520 4948
rect 6388 5000 6440 5006
rect 6388 4942 6440 4948
rect 6572 5000 6624 5006
rect 6572 4942 6624 4948
rect 6664 5000 6716 5006
rect 6664 4942 6716 4948
rect 3732 4734 3760 4942
rect 4982 4900 5358 4920
rect 5038 4898 5062 4900
rect 5118 4898 5142 4900
rect 5198 4898 5222 4900
rect 5278 4898 5302 4900
rect 5038 4846 5048 4898
rect 5292 4846 5302 4898
rect 5038 4844 5062 4846
rect 5118 4844 5142 4846
rect 5198 4844 5222 4846
rect 5278 4844 5302 4846
rect 4982 4824 5358 4844
rect 3720 4728 3772 4734
rect 3720 4670 3772 4676
rect 5480 4666 5508 4942
rect 6400 4802 6428 4942
rect 6388 4796 6440 4802
rect 6388 4738 6440 4744
rect 6584 4734 6612 4942
rect 6572 4728 6624 4734
rect 6572 4670 6624 4676
rect 5468 4660 5520 4666
rect 5468 4602 5520 4608
rect 6296 4660 6348 4666
rect 6296 4602 6348 4608
rect 6664 4660 6716 4666
rect 6664 4602 6716 4608
rect 6308 4546 6336 4602
rect 6308 4518 6520 4546
rect 5100 4456 5152 4462
rect 5100 4398 5152 4404
rect 6388 4456 6440 4462
rect 6388 4398 6440 4404
rect 4017 4356 4393 4376
rect 4073 4354 4097 4356
rect 4153 4354 4177 4356
rect 4233 4354 4257 4356
rect 4313 4354 4337 4356
rect 4073 4302 4083 4354
rect 4327 4302 4337 4354
rect 4073 4300 4097 4302
rect 4153 4300 4177 4302
rect 4233 4300 4257 4302
rect 4313 4300 4337 4302
rect 4017 4280 4393 4300
rect 5112 3986 5140 4398
rect 5948 4356 6324 4376
rect 6004 4354 6028 4356
rect 6084 4354 6108 4356
rect 6164 4354 6188 4356
rect 6244 4354 6268 4356
rect 6004 4302 6014 4354
rect 6258 4302 6268 4354
rect 6004 4300 6028 4302
rect 6084 4300 6108 4302
rect 6164 4300 6188 4302
rect 6244 4300 6268 4302
rect 5948 4280 6324 4300
rect 6400 4054 6428 4398
rect 6492 4190 6520 4518
rect 6480 4184 6532 4190
rect 6480 4126 6532 4132
rect 6676 4054 6704 4602
rect 6388 4048 6440 4054
rect 6388 3990 6440 3996
rect 6664 4048 6716 4054
rect 6664 3990 6716 3996
rect 5100 3980 5152 3986
rect 5100 3922 5152 3928
rect 3168 3912 3220 3918
rect 3168 3854 3220 3860
rect 2136 2412 2936 2510
rect 3180 2412 3208 3854
rect 4982 3812 5358 3832
rect 5038 3810 5062 3812
rect 5118 3810 5142 3812
rect 5198 3810 5222 3812
rect 5278 3810 5302 3812
rect 5038 3758 5048 3810
rect 5292 3758 5302 3810
rect 5038 3756 5062 3758
rect 5118 3756 5142 3758
rect 5198 3756 5222 3758
rect 5278 3756 5302 3758
rect 4982 3736 5358 3756
rect 6400 3578 6428 3990
rect 6768 3714 6796 5554
rect 7044 5142 7072 5554
rect 7400 5544 7452 5550
rect 7400 5486 7452 5492
rect 7412 5142 7440 5486
rect 7596 5346 7624 5622
rect 7878 5444 8254 5464
rect 7934 5442 7958 5444
rect 8014 5442 8038 5444
rect 8094 5442 8118 5444
rect 8174 5442 8198 5444
rect 7934 5390 7944 5442
rect 8188 5390 8198 5442
rect 7934 5388 7958 5390
rect 8014 5388 8038 5390
rect 8094 5388 8118 5390
rect 8174 5388 8198 5390
rect 7878 5368 8254 5388
rect 7584 5340 7636 5346
rect 7584 5282 7636 5288
rect 7032 5136 7084 5142
rect 7032 5078 7084 5084
rect 7400 5136 7452 5142
rect 7400 5078 7452 5084
rect 7492 5136 7544 5142
rect 7492 5078 7544 5084
rect 7308 5068 7360 5074
rect 7308 5010 7360 5016
rect 6913 4900 7289 4920
rect 6969 4898 6993 4900
rect 7049 4898 7073 4900
rect 7129 4898 7153 4900
rect 7209 4898 7233 4900
rect 6969 4846 6979 4898
rect 7223 4846 7233 4898
rect 6969 4844 6993 4846
rect 7049 4844 7073 4846
rect 7129 4844 7153 4846
rect 7209 4844 7233 4846
rect 6913 4824 7289 4844
rect 7320 4258 7348 5010
rect 7400 5000 7452 5006
rect 7400 4942 7452 4948
rect 7412 4666 7440 4942
rect 7400 4660 7452 4666
rect 7400 4602 7452 4608
rect 7504 4530 7532 5078
rect 8332 5074 8360 5690
rect 9336 5080 10136 5178
rect 9160 5074 10136 5080
rect 7676 5068 7728 5074
rect 7676 5010 7728 5016
rect 8320 5068 8372 5074
rect 8320 5010 8372 5016
rect 9148 5068 10136 5074
rect 9200 5052 10136 5068
rect 9148 5010 9200 5016
rect 7492 4524 7544 4530
rect 7492 4466 7544 4472
rect 7688 4258 7716 5010
rect 9336 4954 10136 5052
rect 7768 4660 7820 4666
rect 7768 4602 7820 4608
rect 6940 4252 6992 4258
rect 6940 4194 6992 4200
rect 7308 4252 7360 4258
rect 7308 4194 7360 4200
rect 7676 4252 7728 4258
rect 7676 4194 7728 4200
rect 6952 4054 6980 4194
rect 6940 4048 6992 4054
rect 6940 3990 6992 3996
rect 6913 3812 7289 3832
rect 6969 3810 6993 3812
rect 7049 3810 7073 3812
rect 7129 3810 7153 3812
rect 7209 3810 7233 3812
rect 6969 3758 6979 3810
rect 7223 3758 7233 3810
rect 6969 3756 6993 3758
rect 7049 3756 7073 3758
rect 7129 3756 7153 3758
rect 7209 3756 7233 3758
rect 6913 3736 7289 3756
rect 7780 3714 7808 4602
rect 7878 4356 8254 4376
rect 7934 4354 7958 4356
rect 8014 4354 8038 4356
rect 8094 4354 8118 4356
rect 8174 4354 8198 4356
rect 7934 4302 7944 4354
rect 8188 4302 8198 4354
rect 7934 4300 7958 4302
rect 8014 4300 8038 4302
rect 8094 4300 8118 4302
rect 8174 4300 8198 4302
rect 7878 4280 8254 4300
rect 6756 3708 6808 3714
rect 6756 3650 6808 3656
rect 7768 3708 7820 3714
rect 7768 3650 7820 3656
rect 6388 3572 6440 3578
rect 6388 3514 6440 3520
rect 9148 3572 9200 3578
rect 9148 3514 9200 3520
rect 4017 3268 4393 3288
rect 4073 3266 4097 3268
rect 4153 3266 4177 3268
rect 4233 3266 4257 3268
rect 4313 3266 4337 3268
rect 4073 3214 4083 3266
rect 4327 3214 4337 3266
rect 4073 3212 4097 3214
rect 4153 3212 4177 3214
rect 4233 3212 4257 3214
rect 4313 3212 4337 3214
rect 4017 3192 4393 3212
rect 5948 3268 6324 3288
rect 6004 3266 6028 3268
rect 6084 3266 6108 3268
rect 6164 3266 6188 3268
rect 6244 3266 6268 3268
rect 6004 3214 6014 3266
rect 6258 3214 6268 3266
rect 6004 3212 6028 3214
rect 6084 3212 6108 3214
rect 6164 3212 6188 3214
rect 6244 3212 6268 3214
rect 5948 3192 6324 3212
rect 7878 3268 8254 3288
rect 7934 3266 7958 3268
rect 8014 3266 8038 3268
rect 8094 3266 8118 3268
rect 8174 3266 8198 3268
rect 7934 3214 7944 3266
rect 8188 3214 8198 3266
rect 7934 3212 7958 3214
rect 8014 3212 8038 3214
rect 8094 3212 8118 3214
rect 8174 3212 8198 3214
rect 7878 3192 8254 3212
rect 2136 2384 3208 2412
rect 9160 2412 9188 3514
rect 9336 2412 10136 2510
rect 9160 2384 10136 2412
rect 2136 2286 2936 2384
rect 9336 2286 10136 2384
<< via2 >>
rect 4017 6530 4073 6532
rect 4097 6530 4153 6532
rect 4177 6530 4233 6532
rect 4257 6530 4313 6532
rect 4337 6530 4393 6532
rect 4017 6478 4019 6530
rect 4019 6478 4071 6530
rect 4071 6478 4073 6530
rect 4097 6478 4135 6530
rect 4135 6478 4147 6530
rect 4147 6478 4153 6530
rect 4177 6478 4199 6530
rect 4199 6478 4211 6530
rect 4211 6478 4233 6530
rect 4257 6478 4263 6530
rect 4263 6478 4275 6530
rect 4275 6478 4313 6530
rect 4337 6478 4339 6530
rect 4339 6478 4391 6530
rect 4391 6478 4393 6530
rect 4017 6476 4073 6478
rect 4097 6476 4153 6478
rect 4177 6476 4233 6478
rect 4257 6476 4313 6478
rect 4337 6476 4393 6478
rect 5948 6530 6004 6532
rect 6028 6530 6084 6532
rect 6108 6530 6164 6532
rect 6188 6530 6244 6532
rect 6268 6530 6324 6532
rect 5948 6478 5950 6530
rect 5950 6478 6002 6530
rect 6002 6478 6004 6530
rect 6028 6478 6066 6530
rect 6066 6478 6078 6530
rect 6078 6478 6084 6530
rect 6108 6478 6130 6530
rect 6130 6478 6142 6530
rect 6142 6478 6164 6530
rect 6188 6478 6194 6530
rect 6194 6478 6206 6530
rect 6206 6478 6244 6530
rect 6268 6478 6270 6530
rect 6270 6478 6322 6530
rect 6322 6478 6324 6530
rect 5948 6476 6004 6478
rect 6028 6476 6084 6478
rect 6108 6476 6164 6478
rect 6188 6476 6244 6478
rect 6268 6476 6324 6478
rect 7878 6530 7934 6532
rect 7958 6530 8014 6532
rect 8038 6530 8094 6532
rect 8118 6530 8174 6532
rect 8198 6530 8254 6532
rect 7878 6478 7880 6530
rect 7880 6478 7932 6530
rect 7932 6478 7934 6530
rect 7958 6478 7996 6530
rect 7996 6478 8008 6530
rect 8008 6478 8014 6530
rect 8038 6478 8060 6530
rect 8060 6478 8072 6530
rect 8072 6478 8094 6530
rect 8118 6478 8124 6530
rect 8124 6478 8136 6530
rect 8136 6478 8174 6530
rect 8198 6478 8200 6530
rect 8200 6478 8252 6530
rect 8252 6478 8254 6530
rect 7878 6476 7934 6478
rect 7958 6476 8014 6478
rect 8038 6476 8094 6478
rect 8118 6476 8174 6478
rect 8198 6476 8254 6478
rect 4982 5986 5038 5988
rect 5062 5986 5118 5988
rect 5142 5986 5198 5988
rect 5222 5986 5278 5988
rect 5302 5986 5358 5988
rect 4982 5934 4984 5986
rect 4984 5934 5036 5986
rect 5036 5934 5038 5986
rect 5062 5934 5100 5986
rect 5100 5934 5112 5986
rect 5112 5934 5118 5986
rect 5142 5934 5164 5986
rect 5164 5934 5176 5986
rect 5176 5934 5198 5986
rect 5222 5934 5228 5986
rect 5228 5934 5240 5986
rect 5240 5934 5278 5986
rect 5302 5934 5304 5986
rect 5304 5934 5356 5986
rect 5356 5934 5358 5986
rect 4982 5932 5038 5934
rect 5062 5932 5118 5934
rect 5142 5932 5198 5934
rect 5222 5932 5278 5934
rect 5302 5932 5358 5934
rect 4017 5442 4073 5444
rect 4097 5442 4153 5444
rect 4177 5442 4233 5444
rect 4257 5442 4313 5444
rect 4337 5442 4393 5444
rect 4017 5390 4019 5442
rect 4019 5390 4071 5442
rect 4071 5390 4073 5442
rect 4097 5390 4135 5442
rect 4135 5390 4147 5442
rect 4147 5390 4153 5442
rect 4177 5390 4199 5442
rect 4199 5390 4211 5442
rect 4211 5390 4233 5442
rect 4257 5390 4263 5442
rect 4263 5390 4275 5442
rect 4275 5390 4313 5442
rect 4337 5390 4339 5442
rect 4339 5390 4391 5442
rect 4391 5390 4393 5442
rect 4017 5388 4073 5390
rect 4097 5388 4153 5390
rect 4177 5388 4233 5390
rect 4257 5388 4313 5390
rect 4337 5388 4393 5390
rect 5948 5442 6004 5444
rect 6028 5442 6084 5444
rect 6108 5442 6164 5444
rect 6188 5442 6244 5444
rect 6268 5442 6324 5444
rect 5948 5390 5950 5442
rect 5950 5390 6002 5442
rect 6002 5390 6004 5442
rect 6028 5390 6066 5442
rect 6066 5390 6078 5442
rect 6078 5390 6084 5442
rect 6108 5390 6130 5442
rect 6130 5390 6142 5442
rect 6142 5390 6164 5442
rect 6188 5390 6194 5442
rect 6194 5390 6206 5442
rect 6206 5390 6244 5442
rect 6268 5390 6270 5442
rect 6270 5390 6322 5442
rect 6322 5390 6324 5442
rect 5948 5388 6004 5390
rect 6028 5388 6084 5390
rect 6108 5388 6164 5390
rect 6188 5388 6244 5390
rect 6268 5388 6324 5390
rect 6913 5986 6969 5988
rect 6993 5986 7049 5988
rect 7073 5986 7129 5988
rect 7153 5986 7209 5988
rect 7233 5986 7289 5988
rect 6913 5934 6915 5986
rect 6915 5934 6967 5986
rect 6967 5934 6969 5986
rect 6993 5934 7031 5986
rect 7031 5934 7043 5986
rect 7043 5934 7049 5986
rect 7073 5934 7095 5986
rect 7095 5934 7107 5986
rect 7107 5934 7129 5986
rect 7153 5934 7159 5986
rect 7159 5934 7171 5986
rect 7171 5934 7209 5986
rect 7233 5934 7235 5986
rect 7235 5934 7287 5986
rect 7287 5934 7289 5986
rect 6913 5932 6969 5934
rect 6993 5932 7049 5934
rect 7073 5932 7129 5934
rect 7153 5932 7209 5934
rect 7233 5932 7289 5934
rect 4982 4898 5038 4900
rect 5062 4898 5118 4900
rect 5142 4898 5198 4900
rect 5222 4898 5278 4900
rect 5302 4898 5358 4900
rect 4982 4846 4984 4898
rect 4984 4846 5036 4898
rect 5036 4846 5038 4898
rect 5062 4846 5100 4898
rect 5100 4846 5112 4898
rect 5112 4846 5118 4898
rect 5142 4846 5164 4898
rect 5164 4846 5176 4898
rect 5176 4846 5198 4898
rect 5222 4846 5228 4898
rect 5228 4846 5240 4898
rect 5240 4846 5278 4898
rect 5302 4846 5304 4898
rect 5304 4846 5356 4898
rect 5356 4846 5358 4898
rect 4982 4844 5038 4846
rect 5062 4844 5118 4846
rect 5142 4844 5198 4846
rect 5222 4844 5278 4846
rect 5302 4844 5358 4846
rect 4017 4354 4073 4356
rect 4097 4354 4153 4356
rect 4177 4354 4233 4356
rect 4257 4354 4313 4356
rect 4337 4354 4393 4356
rect 4017 4302 4019 4354
rect 4019 4302 4071 4354
rect 4071 4302 4073 4354
rect 4097 4302 4135 4354
rect 4135 4302 4147 4354
rect 4147 4302 4153 4354
rect 4177 4302 4199 4354
rect 4199 4302 4211 4354
rect 4211 4302 4233 4354
rect 4257 4302 4263 4354
rect 4263 4302 4275 4354
rect 4275 4302 4313 4354
rect 4337 4302 4339 4354
rect 4339 4302 4391 4354
rect 4391 4302 4393 4354
rect 4017 4300 4073 4302
rect 4097 4300 4153 4302
rect 4177 4300 4233 4302
rect 4257 4300 4313 4302
rect 4337 4300 4393 4302
rect 5948 4354 6004 4356
rect 6028 4354 6084 4356
rect 6108 4354 6164 4356
rect 6188 4354 6244 4356
rect 6268 4354 6324 4356
rect 5948 4302 5950 4354
rect 5950 4302 6002 4354
rect 6002 4302 6004 4354
rect 6028 4302 6066 4354
rect 6066 4302 6078 4354
rect 6078 4302 6084 4354
rect 6108 4302 6130 4354
rect 6130 4302 6142 4354
rect 6142 4302 6164 4354
rect 6188 4302 6194 4354
rect 6194 4302 6206 4354
rect 6206 4302 6244 4354
rect 6268 4302 6270 4354
rect 6270 4302 6322 4354
rect 6322 4302 6324 4354
rect 5948 4300 6004 4302
rect 6028 4300 6084 4302
rect 6108 4300 6164 4302
rect 6188 4300 6244 4302
rect 6268 4300 6324 4302
rect 4982 3810 5038 3812
rect 5062 3810 5118 3812
rect 5142 3810 5198 3812
rect 5222 3810 5278 3812
rect 5302 3810 5358 3812
rect 4982 3758 4984 3810
rect 4984 3758 5036 3810
rect 5036 3758 5038 3810
rect 5062 3758 5100 3810
rect 5100 3758 5112 3810
rect 5112 3758 5118 3810
rect 5142 3758 5164 3810
rect 5164 3758 5176 3810
rect 5176 3758 5198 3810
rect 5222 3758 5228 3810
rect 5228 3758 5240 3810
rect 5240 3758 5278 3810
rect 5302 3758 5304 3810
rect 5304 3758 5356 3810
rect 5356 3758 5358 3810
rect 4982 3756 5038 3758
rect 5062 3756 5118 3758
rect 5142 3756 5198 3758
rect 5222 3756 5278 3758
rect 5302 3756 5358 3758
rect 7878 5442 7934 5444
rect 7958 5442 8014 5444
rect 8038 5442 8094 5444
rect 8118 5442 8174 5444
rect 8198 5442 8254 5444
rect 7878 5390 7880 5442
rect 7880 5390 7932 5442
rect 7932 5390 7934 5442
rect 7958 5390 7996 5442
rect 7996 5390 8008 5442
rect 8008 5390 8014 5442
rect 8038 5390 8060 5442
rect 8060 5390 8072 5442
rect 8072 5390 8094 5442
rect 8118 5390 8124 5442
rect 8124 5390 8136 5442
rect 8136 5390 8174 5442
rect 8198 5390 8200 5442
rect 8200 5390 8252 5442
rect 8252 5390 8254 5442
rect 7878 5388 7934 5390
rect 7958 5388 8014 5390
rect 8038 5388 8094 5390
rect 8118 5388 8174 5390
rect 8198 5388 8254 5390
rect 6913 4898 6969 4900
rect 6993 4898 7049 4900
rect 7073 4898 7129 4900
rect 7153 4898 7209 4900
rect 7233 4898 7289 4900
rect 6913 4846 6915 4898
rect 6915 4846 6967 4898
rect 6967 4846 6969 4898
rect 6993 4846 7031 4898
rect 7031 4846 7043 4898
rect 7043 4846 7049 4898
rect 7073 4846 7095 4898
rect 7095 4846 7107 4898
rect 7107 4846 7129 4898
rect 7153 4846 7159 4898
rect 7159 4846 7171 4898
rect 7171 4846 7209 4898
rect 7233 4846 7235 4898
rect 7235 4846 7287 4898
rect 7287 4846 7289 4898
rect 6913 4844 6969 4846
rect 6993 4844 7049 4846
rect 7073 4844 7129 4846
rect 7153 4844 7209 4846
rect 7233 4844 7289 4846
rect 6913 3810 6969 3812
rect 6993 3810 7049 3812
rect 7073 3810 7129 3812
rect 7153 3810 7209 3812
rect 7233 3810 7289 3812
rect 6913 3758 6915 3810
rect 6915 3758 6967 3810
rect 6967 3758 6969 3810
rect 6993 3758 7031 3810
rect 7031 3758 7043 3810
rect 7043 3758 7049 3810
rect 7073 3758 7095 3810
rect 7095 3758 7107 3810
rect 7107 3758 7129 3810
rect 7153 3758 7159 3810
rect 7159 3758 7171 3810
rect 7171 3758 7209 3810
rect 7233 3758 7235 3810
rect 7235 3758 7287 3810
rect 7287 3758 7289 3810
rect 6913 3756 6969 3758
rect 6993 3756 7049 3758
rect 7073 3756 7129 3758
rect 7153 3756 7209 3758
rect 7233 3756 7289 3758
rect 7878 4354 7934 4356
rect 7958 4354 8014 4356
rect 8038 4354 8094 4356
rect 8118 4354 8174 4356
rect 8198 4354 8254 4356
rect 7878 4302 7880 4354
rect 7880 4302 7932 4354
rect 7932 4302 7934 4354
rect 7958 4302 7996 4354
rect 7996 4302 8008 4354
rect 8008 4302 8014 4354
rect 8038 4302 8060 4354
rect 8060 4302 8072 4354
rect 8072 4302 8094 4354
rect 8118 4302 8124 4354
rect 8124 4302 8136 4354
rect 8136 4302 8174 4354
rect 8198 4302 8200 4354
rect 8200 4302 8252 4354
rect 8252 4302 8254 4354
rect 7878 4300 7934 4302
rect 7958 4300 8014 4302
rect 8038 4300 8094 4302
rect 8118 4300 8174 4302
rect 8198 4300 8254 4302
rect 4017 3266 4073 3268
rect 4097 3266 4153 3268
rect 4177 3266 4233 3268
rect 4257 3266 4313 3268
rect 4337 3266 4393 3268
rect 4017 3214 4019 3266
rect 4019 3214 4071 3266
rect 4071 3214 4073 3266
rect 4097 3214 4135 3266
rect 4135 3214 4147 3266
rect 4147 3214 4153 3266
rect 4177 3214 4199 3266
rect 4199 3214 4211 3266
rect 4211 3214 4233 3266
rect 4257 3214 4263 3266
rect 4263 3214 4275 3266
rect 4275 3214 4313 3266
rect 4337 3214 4339 3266
rect 4339 3214 4391 3266
rect 4391 3214 4393 3266
rect 4017 3212 4073 3214
rect 4097 3212 4153 3214
rect 4177 3212 4233 3214
rect 4257 3212 4313 3214
rect 4337 3212 4393 3214
rect 5948 3266 6004 3268
rect 6028 3266 6084 3268
rect 6108 3266 6164 3268
rect 6188 3266 6244 3268
rect 6268 3266 6324 3268
rect 5948 3214 5950 3266
rect 5950 3214 6002 3266
rect 6002 3214 6004 3266
rect 6028 3214 6066 3266
rect 6066 3214 6078 3266
rect 6078 3214 6084 3266
rect 6108 3214 6130 3266
rect 6130 3214 6142 3266
rect 6142 3214 6164 3266
rect 6188 3214 6194 3266
rect 6194 3214 6206 3266
rect 6206 3214 6244 3266
rect 6268 3214 6270 3266
rect 6270 3214 6322 3266
rect 6322 3214 6324 3266
rect 5948 3212 6004 3214
rect 6028 3212 6084 3214
rect 6108 3212 6164 3214
rect 6188 3212 6244 3214
rect 6268 3212 6324 3214
rect 7878 3266 7934 3268
rect 7958 3266 8014 3268
rect 8038 3266 8094 3268
rect 8118 3266 8174 3268
rect 8198 3266 8254 3268
rect 7878 3214 7880 3266
rect 7880 3214 7932 3266
rect 7932 3214 7934 3266
rect 7958 3214 7996 3266
rect 7996 3214 8008 3266
rect 8008 3214 8014 3266
rect 8038 3214 8060 3266
rect 8060 3214 8072 3266
rect 8072 3214 8094 3266
rect 8118 3214 8124 3266
rect 8124 3214 8136 3266
rect 8136 3214 8174 3266
rect 8198 3214 8200 3266
rect 8200 3214 8252 3266
rect 8252 3214 8254 3266
rect 7878 3212 7934 3214
rect 7958 3212 8014 3214
rect 8038 3212 8094 3214
rect 8118 3212 8174 3214
rect 8198 3212 8254 3214
<< metal3 >>
rect 0 9736 12184 9744
rect 0 8952 8 9736
rect 792 8952 4978 9736
rect 5362 8952 6909 9736
rect 7293 8952 11392 9736
rect 12176 8952 12184 9736
rect 0 8944 12184 8952
rect 1140 8596 11044 8604
rect 1140 7812 1148 8596
rect 1932 7812 4013 8596
rect 4397 7812 5944 8596
rect 6328 7812 7874 8596
rect 8258 7812 10252 8596
rect 11036 7812 11044 8596
rect 1140 7804 11044 7812
rect 3995 6536 4415 6537
rect 3995 6472 4013 6536
rect 4077 6472 4093 6536
rect 4157 6472 4173 6536
rect 4237 6472 4253 6536
rect 4317 6472 4333 6536
rect 4397 6472 4415 6536
rect 3995 6471 4415 6472
rect 5926 6536 6346 6537
rect 5926 6472 5944 6536
rect 6008 6472 6024 6536
rect 6088 6472 6104 6536
rect 6168 6472 6184 6536
rect 6248 6472 6264 6536
rect 6328 6472 6346 6536
rect 5926 6471 6346 6472
rect 7856 6536 8276 6537
rect 7856 6472 7874 6536
rect 7938 6472 7954 6536
rect 8018 6472 8034 6536
rect 8098 6472 8114 6536
rect 8178 6472 8194 6536
rect 8258 6472 8276 6536
rect 7856 6471 8276 6472
rect 4960 5992 5380 5993
rect 4960 5928 4978 5992
rect 5042 5928 5058 5992
rect 5122 5928 5138 5992
rect 5202 5928 5218 5992
rect 5282 5928 5298 5992
rect 5362 5928 5380 5992
rect 4960 5927 5380 5928
rect 6891 5992 7311 5993
rect 6891 5928 6909 5992
rect 6973 5928 6989 5992
rect 7053 5928 7069 5992
rect 7133 5928 7149 5992
rect 7213 5928 7229 5992
rect 7293 5928 7311 5992
rect 6891 5927 7311 5928
rect 3995 5448 4415 5449
rect 3995 5384 4013 5448
rect 4077 5384 4093 5448
rect 4157 5384 4173 5448
rect 4237 5384 4253 5448
rect 4317 5384 4333 5448
rect 4397 5384 4415 5448
rect 3995 5383 4415 5384
rect 5926 5448 6346 5449
rect 5926 5384 5944 5448
rect 6008 5384 6024 5448
rect 6088 5384 6104 5448
rect 6168 5384 6184 5448
rect 6248 5384 6264 5448
rect 6328 5384 6346 5448
rect 5926 5383 6346 5384
rect 7856 5448 8276 5449
rect 7856 5384 7874 5448
rect 7938 5384 7954 5448
rect 8018 5384 8034 5448
rect 8098 5384 8114 5448
rect 8178 5384 8194 5448
rect 8258 5384 8276 5448
rect 7856 5383 8276 5384
rect 4960 4904 5380 4905
rect 4960 4840 4978 4904
rect 5042 4840 5058 4904
rect 5122 4840 5138 4904
rect 5202 4840 5218 4904
rect 5282 4840 5298 4904
rect 5362 4840 5380 4904
rect 4960 4839 5380 4840
rect 6891 4904 7311 4905
rect 6891 4840 6909 4904
rect 6973 4840 6989 4904
rect 7053 4840 7069 4904
rect 7133 4840 7149 4904
rect 7213 4840 7229 4904
rect 7293 4840 7311 4904
rect 6891 4839 7311 4840
rect 3995 4360 4415 4361
rect 3995 4296 4013 4360
rect 4077 4296 4093 4360
rect 4157 4296 4173 4360
rect 4237 4296 4253 4360
rect 4317 4296 4333 4360
rect 4397 4296 4415 4360
rect 3995 4295 4415 4296
rect 5926 4360 6346 4361
rect 5926 4296 5944 4360
rect 6008 4296 6024 4360
rect 6088 4296 6104 4360
rect 6168 4296 6184 4360
rect 6248 4296 6264 4360
rect 6328 4296 6346 4360
rect 5926 4295 6346 4296
rect 7856 4360 8276 4361
rect 7856 4296 7874 4360
rect 7938 4296 7954 4360
rect 8018 4296 8034 4360
rect 8098 4296 8114 4360
rect 8178 4296 8194 4360
rect 8258 4296 8276 4360
rect 7856 4295 8276 4296
rect 4960 3816 5380 3817
rect 4960 3752 4978 3816
rect 5042 3752 5058 3816
rect 5122 3752 5138 3816
rect 5202 3752 5218 3816
rect 5282 3752 5298 3816
rect 5362 3752 5380 3816
rect 4960 3751 5380 3752
rect 6891 3816 7311 3817
rect 6891 3752 6909 3816
rect 6973 3752 6989 3816
rect 7053 3752 7069 3816
rect 7133 3752 7149 3816
rect 7213 3752 7229 3816
rect 7293 3752 7311 3816
rect 6891 3751 7311 3752
rect 3995 3272 4415 3273
rect 3995 3208 4013 3272
rect 4077 3208 4093 3272
rect 4157 3208 4173 3272
rect 4237 3208 4253 3272
rect 4317 3208 4333 3272
rect 4397 3208 4415 3272
rect 3995 3207 4415 3208
rect 5926 3272 6346 3273
rect 5926 3208 5944 3272
rect 6008 3208 6024 3272
rect 6088 3208 6104 3272
rect 6168 3208 6184 3272
rect 6248 3208 6264 3272
rect 6328 3208 6346 3272
rect 5926 3207 6346 3208
rect 7856 3272 8276 3273
rect 7856 3208 7874 3272
rect 7938 3208 7954 3272
rect 8018 3208 8034 3272
rect 8098 3208 8114 3272
rect 8178 3208 8194 3272
rect 8258 3208 8276 3272
rect 7856 3207 8276 3208
rect 1140 1932 11044 1940
rect 1140 1148 1148 1932
rect 1932 1148 4013 1932
rect 4397 1148 5944 1932
rect 6328 1148 7874 1932
rect 8258 1148 10252 1932
rect 11036 1148 11044 1932
rect 1140 1140 11044 1148
rect 0 792 12184 800
rect 0 8 8 792
rect 792 8 4978 792
rect 5362 8 6909 792
rect 7293 8 11392 792
rect 12176 8 12184 792
rect 0 0 12184 8
<< via3 >>
rect 8 8952 792 9736
rect 4978 8952 5362 9736
rect 6909 8952 7293 9736
rect 11392 8952 12176 9736
rect 1148 7812 1932 8596
rect 4013 7812 4397 8596
rect 5944 7812 6328 8596
rect 7874 7812 8258 8596
rect 10252 7812 11036 8596
rect 4013 6532 4077 6536
rect 4013 6476 4017 6532
rect 4017 6476 4073 6532
rect 4073 6476 4077 6532
rect 4013 6472 4077 6476
rect 4093 6532 4157 6536
rect 4093 6476 4097 6532
rect 4097 6476 4153 6532
rect 4153 6476 4157 6532
rect 4093 6472 4157 6476
rect 4173 6532 4237 6536
rect 4173 6476 4177 6532
rect 4177 6476 4233 6532
rect 4233 6476 4237 6532
rect 4173 6472 4237 6476
rect 4253 6532 4317 6536
rect 4253 6476 4257 6532
rect 4257 6476 4313 6532
rect 4313 6476 4317 6532
rect 4253 6472 4317 6476
rect 4333 6532 4397 6536
rect 4333 6476 4337 6532
rect 4337 6476 4393 6532
rect 4393 6476 4397 6532
rect 4333 6472 4397 6476
rect 5944 6532 6008 6536
rect 5944 6476 5948 6532
rect 5948 6476 6004 6532
rect 6004 6476 6008 6532
rect 5944 6472 6008 6476
rect 6024 6532 6088 6536
rect 6024 6476 6028 6532
rect 6028 6476 6084 6532
rect 6084 6476 6088 6532
rect 6024 6472 6088 6476
rect 6104 6532 6168 6536
rect 6104 6476 6108 6532
rect 6108 6476 6164 6532
rect 6164 6476 6168 6532
rect 6104 6472 6168 6476
rect 6184 6532 6248 6536
rect 6184 6476 6188 6532
rect 6188 6476 6244 6532
rect 6244 6476 6248 6532
rect 6184 6472 6248 6476
rect 6264 6532 6328 6536
rect 6264 6476 6268 6532
rect 6268 6476 6324 6532
rect 6324 6476 6328 6532
rect 6264 6472 6328 6476
rect 7874 6532 7938 6536
rect 7874 6476 7878 6532
rect 7878 6476 7934 6532
rect 7934 6476 7938 6532
rect 7874 6472 7938 6476
rect 7954 6532 8018 6536
rect 7954 6476 7958 6532
rect 7958 6476 8014 6532
rect 8014 6476 8018 6532
rect 7954 6472 8018 6476
rect 8034 6532 8098 6536
rect 8034 6476 8038 6532
rect 8038 6476 8094 6532
rect 8094 6476 8098 6532
rect 8034 6472 8098 6476
rect 8114 6532 8178 6536
rect 8114 6476 8118 6532
rect 8118 6476 8174 6532
rect 8174 6476 8178 6532
rect 8114 6472 8178 6476
rect 8194 6532 8258 6536
rect 8194 6476 8198 6532
rect 8198 6476 8254 6532
rect 8254 6476 8258 6532
rect 8194 6472 8258 6476
rect 4978 5988 5042 5992
rect 4978 5932 4982 5988
rect 4982 5932 5038 5988
rect 5038 5932 5042 5988
rect 4978 5928 5042 5932
rect 5058 5988 5122 5992
rect 5058 5932 5062 5988
rect 5062 5932 5118 5988
rect 5118 5932 5122 5988
rect 5058 5928 5122 5932
rect 5138 5988 5202 5992
rect 5138 5932 5142 5988
rect 5142 5932 5198 5988
rect 5198 5932 5202 5988
rect 5138 5928 5202 5932
rect 5218 5988 5282 5992
rect 5218 5932 5222 5988
rect 5222 5932 5278 5988
rect 5278 5932 5282 5988
rect 5218 5928 5282 5932
rect 5298 5988 5362 5992
rect 5298 5932 5302 5988
rect 5302 5932 5358 5988
rect 5358 5932 5362 5988
rect 5298 5928 5362 5932
rect 6909 5988 6973 5992
rect 6909 5932 6913 5988
rect 6913 5932 6969 5988
rect 6969 5932 6973 5988
rect 6909 5928 6973 5932
rect 6989 5988 7053 5992
rect 6989 5932 6993 5988
rect 6993 5932 7049 5988
rect 7049 5932 7053 5988
rect 6989 5928 7053 5932
rect 7069 5988 7133 5992
rect 7069 5932 7073 5988
rect 7073 5932 7129 5988
rect 7129 5932 7133 5988
rect 7069 5928 7133 5932
rect 7149 5988 7213 5992
rect 7149 5932 7153 5988
rect 7153 5932 7209 5988
rect 7209 5932 7213 5988
rect 7149 5928 7213 5932
rect 7229 5988 7293 5992
rect 7229 5932 7233 5988
rect 7233 5932 7289 5988
rect 7289 5932 7293 5988
rect 7229 5928 7293 5932
rect 4013 5444 4077 5448
rect 4013 5388 4017 5444
rect 4017 5388 4073 5444
rect 4073 5388 4077 5444
rect 4013 5384 4077 5388
rect 4093 5444 4157 5448
rect 4093 5388 4097 5444
rect 4097 5388 4153 5444
rect 4153 5388 4157 5444
rect 4093 5384 4157 5388
rect 4173 5444 4237 5448
rect 4173 5388 4177 5444
rect 4177 5388 4233 5444
rect 4233 5388 4237 5444
rect 4173 5384 4237 5388
rect 4253 5444 4317 5448
rect 4253 5388 4257 5444
rect 4257 5388 4313 5444
rect 4313 5388 4317 5444
rect 4253 5384 4317 5388
rect 4333 5444 4397 5448
rect 4333 5388 4337 5444
rect 4337 5388 4393 5444
rect 4393 5388 4397 5444
rect 4333 5384 4397 5388
rect 5944 5444 6008 5448
rect 5944 5388 5948 5444
rect 5948 5388 6004 5444
rect 6004 5388 6008 5444
rect 5944 5384 6008 5388
rect 6024 5444 6088 5448
rect 6024 5388 6028 5444
rect 6028 5388 6084 5444
rect 6084 5388 6088 5444
rect 6024 5384 6088 5388
rect 6104 5444 6168 5448
rect 6104 5388 6108 5444
rect 6108 5388 6164 5444
rect 6164 5388 6168 5444
rect 6104 5384 6168 5388
rect 6184 5444 6248 5448
rect 6184 5388 6188 5444
rect 6188 5388 6244 5444
rect 6244 5388 6248 5444
rect 6184 5384 6248 5388
rect 6264 5444 6328 5448
rect 6264 5388 6268 5444
rect 6268 5388 6324 5444
rect 6324 5388 6328 5444
rect 6264 5384 6328 5388
rect 7874 5444 7938 5448
rect 7874 5388 7878 5444
rect 7878 5388 7934 5444
rect 7934 5388 7938 5444
rect 7874 5384 7938 5388
rect 7954 5444 8018 5448
rect 7954 5388 7958 5444
rect 7958 5388 8014 5444
rect 8014 5388 8018 5444
rect 7954 5384 8018 5388
rect 8034 5444 8098 5448
rect 8034 5388 8038 5444
rect 8038 5388 8094 5444
rect 8094 5388 8098 5444
rect 8034 5384 8098 5388
rect 8114 5444 8178 5448
rect 8114 5388 8118 5444
rect 8118 5388 8174 5444
rect 8174 5388 8178 5444
rect 8114 5384 8178 5388
rect 8194 5444 8258 5448
rect 8194 5388 8198 5444
rect 8198 5388 8254 5444
rect 8254 5388 8258 5444
rect 8194 5384 8258 5388
rect 4978 4900 5042 4904
rect 4978 4844 4982 4900
rect 4982 4844 5038 4900
rect 5038 4844 5042 4900
rect 4978 4840 5042 4844
rect 5058 4900 5122 4904
rect 5058 4844 5062 4900
rect 5062 4844 5118 4900
rect 5118 4844 5122 4900
rect 5058 4840 5122 4844
rect 5138 4900 5202 4904
rect 5138 4844 5142 4900
rect 5142 4844 5198 4900
rect 5198 4844 5202 4900
rect 5138 4840 5202 4844
rect 5218 4900 5282 4904
rect 5218 4844 5222 4900
rect 5222 4844 5278 4900
rect 5278 4844 5282 4900
rect 5218 4840 5282 4844
rect 5298 4900 5362 4904
rect 5298 4844 5302 4900
rect 5302 4844 5358 4900
rect 5358 4844 5362 4900
rect 5298 4840 5362 4844
rect 6909 4900 6973 4904
rect 6909 4844 6913 4900
rect 6913 4844 6969 4900
rect 6969 4844 6973 4900
rect 6909 4840 6973 4844
rect 6989 4900 7053 4904
rect 6989 4844 6993 4900
rect 6993 4844 7049 4900
rect 7049 4844 7053 4900
rect 6989 4840 7053 4844
rect 7069 4900 7133 4904
rect 7069 4844 7073 4900
rect 7073 4844 7129 4900
rect 7129 4844 7133 4900
rect 7069 4840 7133 4844
rect 7149 4900 7213 4904
rect 7149 4844 7153 4900
rect 7153 4844 7209 4900
rect 7209 4844 7213 4900
rect 7149 4840 7213 4844
rect 7229 4900 7293 4904
rect 7229 4844 7233 4900
rect 7233 4844 7289 4900
rect 7289 4844 7293 4900
rect 7229 4840 7293 4844
rect 4013 4356 4077 4360
rect 4013 4300 4017 4356
rect 4017 4300 4073 4356
rect 4073 4300 4077 4356
rect 4013 4296 4077 4300
rect 4093 4356 4157 4360
rect 4093 4300 4097 4356
rect 4097 4300 4153 4356
rect 4153 4300 4157 4356
rect 4093 4296 4157 4300
rect 4173 4356 4237 4360
rect 4173 4300 4177 4356
rect 4177 4300 4233 4356
rect 4233 4300 4237 4356
rect 4173 4296 4237 4300
rect 4253 4356 4317 4360
rect 4253 4300 4257 4356
rect 4257 4300 4313 4356
rect 4313 4300 4317 4356
rect 4253 4296 4317 4300
rect 4333 4356 4397 4360
rect 4333 4300 4337 4356
rect 4337 4300 4393 4356
rect 4393 4300 4397 4356
rect 4333 4296 4397 4300
rect 5944 4356 6008 4360
rect 5944 4300 5948 4356
rect 5948 4300 6004 4356
rect 6004 4300 6008 4356
rect 5944 4296 6008 4300
rect 6024 4356 6088 4360
rect 6024 4300 6028 4356
rect 6028 4300 6084 4356
rect 6084 4300 6088 4356
rect 6024 4296 6088 4300
rect 6104 4356 6168 4360
rect 6104 4300 6108 4356
rect 6108 4300 6164 4356
rect 6164 4300 6168 4356
rect 6104 4296 6168 4300
rect 6184 4356 6248 4360
rect 6184 4300 6188 4356
rect 6188 4300 6244 4356
rect 6244 4300 6248 4356
rect 6184 4296 6248 4300
rect 6264 4356 6328 4360
rect 6264 4300 6268 4356
rect 6268 4300 6324 4356
rect 6324 4300 6328 4356
rect 6264 4296 6328 4300
rect 7874 4356 7938 4360
rect 7874 4300 7878 4356
rect 7878 4300 7934 4356
rect 7934 4300 7938 4356
rect 7874 4296 7938 4300
rect 7954 4356 8018 4360
rect 7954 4300 7958 4356
rect 7958 4300 8014 4356
rect 8014 4300 8018 4356
rect 7954 4296 8018 4300
rect 8034 4356 8098 4360
rect 8034 4300 8038 4356
rect 8038 4300 8094 4356
rect 8094 4300 8098 4356
rect 8034 4296 8098 4300
rect 8114 4356 8178 4360
rect 8114 4300 8118 4356
rect 8118 4300 8174 4356
rect 8174 4300 8178 4356
rect 8114 4296 8178 4300
rect 8194 4356 8258 4360
rect 8194 4300 8198 4356
rect 8198 4300 8254 4356
rect 8254 4300 8258 4356
rect 8194 4296 8258 4300
rect 4978 3812 5042 3816
rect 4978 3756 4982 3812
rect 4982 3756 5038 3812
rect 5038 3756 5042 3812
rect 4978 3752 5042 3756
rect 5058 3812 5122 3816
rect 5058 3756 5062 3812
rect 5062 3756 5118 3812
rect 5118 3756 5122 3812
rect 5058 3752 5122 3756
rect 5138 3812 5202 3816
rect 5138 3756 5142 3812
rect 5142 3756 5198 3812
rect 5198 3756 5202 3812
rect 5138 3752 5202 3756
rect 5218 3812 5282 3816
rect 5218 3756 5222 3812
rect 5222 3756 5278 3812
rect 5278 3756 5282 3812
rect 5218 3752 5282 3756
rect 5298 3812 5362 3816
rect 5298 3756 5302 3812
rect 5302 3756 5358 3812
rect 5358 3756 5362 3812
rect 5298 3752 5362 3756
rect 6909 3812 6973 3816
rect 6909 3756 6913 3812
rect 6913 3756 6969 3812
rect 6969 3756 6973 3812
rect 6909 3752 6973 3756
rect 6989 3812 7053 3816
rect 6989 3756 6993 3812
rect 6993 3756 7049 3812
rect 7049 3756 7053 3812
rect 6989 3752 7053 3756
rect 7069 3812 7133 3816
rect 7069 3756 7073 3812
rect 7073 3756 7129 3812
rect 7129 3756 7133 3812
rect 7069 3752 7133 3756
rect 7149 3812 7213 3816
rect 7149 3756 7153 3812
rect 7153 3756 7209 3812
rect 7209 3756 7213 3812
rect 7149 3752 7213 3756
rect 7229 3812 7293 3816
rect 7229 3756 7233 3812
rect 7233 3756 7289 3812
rect 7289 3756 7293 3812
rect 7229 3752 7293 3756
rect 4013 3268 4077 3272
rect 4013 3212 4017 3268
rect 4017 3212 4073 3268
rect 4073 3212 4077 3268
rect 4013 3208 4077 3212
rect 4093 3268 4157 3272
rect 4093 3212 4097 3268
rect 4097 3212 4153 3268
rect 4153 3212 4157 3268
rect 4093 3208 4157 3212
rect 4173 3268 4237 3272
rect 4173 3212 4177 3268
rect 4177 3212 4233 3268
rect 4233 3212 4237 3268
rect 4173 3208 4237 3212
rect 4253 3268 4317 3272
rect 4253 3212 4257 3268
rect 4257 3212 4313 3268
rect 4313 3212 4317 3268
rect 4253 3208 4317 3212
rect 4333 3268 4397 3272
rect 4333 3212 4337 3268
rect 4337 3212 4393 3268
rect 4393 3212 4397 3268
rect 4333 3208 4397 3212
rect 5944 3268 6008 3272
rect 5944 3212 5948 3268
rect 5948 3212 6004 3268
rect 6004 3212 6008 3268
rect 5944 3208 6008 3212
rect 6024 3268 6088 3272
rect 6024 3212 6028 3268
rect 6028 3212 6084 3268
rect 6084 3212 6088 3268
rect 6024 3208 6088 3212
rect 6104 3268 6168 3272
rect 6104 3212 6108 3268
rect 6108 3212 6164 3268
rect 6164 3212 6168 3268
rect 6104 3208 6168 3212
rect 6184 3268 6248 3272
rect 6184 3212 6188 3268
rect 6188 3212 6244 3268
rect 6244 3212 6248 3268
rect 6184 3208 6248 3212
rect 6264 3268 6328 3272
rect 6264 3212 6268 3268
rect 6268 3212 6324 3268
rect 6324 3212 6328 3268
rect 6264 3208 6328 3212
rect 7874 3268 7938 3272
rect 7874 3212 7878 3268
rect 7878 3212 7934 3268
rect 7934 3212 7938 3268
rect 7874 3208 7938 3212
rect 7954 3268 8018 3272
rect 7954 3212 7958 3268
rect 7958 3212 8014 3268
rect 8014 3212 8018 3268
rect 7954 3208 8018 3212
rect 8034 3268 8098 3272
rect 8034 3212 8038 3268
rect 8038 3212 8094 3268
rect 8094 3212 8098 3268
rect 8034 3208 8098 3212
rect 8114 3268 8178 3272
rect 8114 3212 8118 3268
rect 8118 3212 8174 3268
rect 8174 3212 8178 3268
rect 8114 3208 8178 3212
rect 8194 3268 8258 3272
rect 8194 3212 8198 3268
rect 8198 3212 8254 3268
rect 8254 3212 8258 3268
rect 8194 3208 8258 3212
rect 1148 1148 1932 1932
rect 4013 1148 4397 1932
rect 5944 1148 6328 1932
rect 7874 1148 8258 1932
rect 10252 1148 11036 1932
rect 8 8 792 792
rect 4978 8 5362 792
rect 6909 8 7293 792
rect 11392 8 12176 792
<< metal4 >>
rect 0 9736 800 9744
rect 0 8952 8 9736
rect 792 8952 800 9736
rect 0 792 800 8952
rect 1140 8596 1940 8604
rect 1140 7812 1148 8596
rect 1932 7812 1940 8596
rect 1140 1932 1940 7812
rect 1140 1148 1148 1932
rect 1932 1148 1940 1932
rect 1140 1140 1940 1148
rect 3995 8596 4415 9744
rect 3995 7812 4013 8596
rect 4397 7812 4415 8596
rect 3995 6536 4415 7812
rect 3995 6472 4013 6536
rect 4077 6472 4093 6536
rect 4157 6472 4173 6536
rect 4237 6472 4253 6536
rect 4317 6472 4333 6536
rect 4397 6472 4415 6536
rect 3995 5448 4415 6472
rect 3995 5384 4013 5448
rect 4077 5384 4093 5448
rect 4157 5384 4173 5448
rect 4237 5384 4253 5448
rect 4317 5384 4333 5448
rect 4397 5384 4415 5448
rect 3995 4360 4415 5384
rect 3995 4296 4013 4360
rect 4077 4296 4093 4360
rect 4157 4296 4173 4360
rect 4237 4296 4253 4360
rect 4317 4296 4333 4360
rect 4397 4296 4415 4360
rect 3995 3272 4415 4296
rect 3995 3208 4013 3272
rect 4077 3208 4093 3272
rect 4157 3208 4173 3272
rect 4237 3208 4253 3272
rect 4317 3208 4333 3272
rect 4397 3208 4415 3272
rect 3995 1932 4415 3208
rect 3995 1148 4013 1932
rect 4397 1148 4415 1932
rect 0 8 8 792
rect 792 8 800 792
rect 0 0 800 8
rect 3995 0 4415 1148
rect 4960 9736 5381 9744
rect 4960 8952 4978 9736
rect 5362 8952 5381 9736
rect 4960 5992 5381 8952
rect 4960 5928 4978 5992
rect 5042 5928 5058 5992
rect 5122 5928 5138 5992
rect 5202 5928 5218 5992
rect 5282 5928 5298 5992
rect 5362 5928 5381 5992
rect 4960 4904 5381 5928
rect 4960 4840 4978 4904
rect 5042 4840 5058 4904
rect 5122 4840 5138 4904
rect 5202 4840 5218 4904
rect 5282 4840 5298 4904
rect 5362 4840 5381 4904
rect 4960 3816 5381 4840
rect 4960 3752 4978 3816
rect 5042 3752 5058 3816
rect 5122 3752 5138 3816
rect 5202 3752 5218 3816
rect 5282 3752 5298 3816
rect 5362 3752 5381 3816
rect 4960 792 5381 3752
rect 4960 8 4978 792
rect 5362 8 5381 792
rect 4960 0 5381 8
rect 5926 8596 6346 9744
rect 5926 7812 5944 8596
rect 6328 7812 6346 8596
rect 5926 6536 6346 7812
rect 5926 6472 5944 6536
rect 6008 6472 6024 6536
rect 6088 6472 6104 6536
rect 6168 6472 6184 6536
rect 6248 6472 6264 6536
rect 6328 6472 6346 6536
rect 5926 5448 6346 6472
rect 5926 5384 5944 5448
rect 6008 5384 6024 5448
rect 6088 5384 6104 5448
rect 6168 5384 6184 5448
rect 6248 5384 6264 5448
rect 6328 5384 6346 5448
rect 5926 4360 6346 5384
rect 5926 4296 5944 4360
rect 6008 4296 6024 4360
rect 6088 4296 6104 4360
rect 6168 4296 6184 4360
rect 6248 4296 6264 4360
rect 6328 4296 6346 4360
rect 5926 3272 6346 4296
rect 5926 3208 5944 3272
rect 6008 3208 6024 3272
rect 6088 3208 6104 3272
rect 6168 3208 6184 3272
rect 6248 3208 6264 3272
rect 6328 3208 6346 3272
rect 5926 1932 6346 3208
rect 5926 1148 5944 1932
rect 6328 1148 6346 1932
rect 5926 0 6346 1148
rect 6891 9736 7311 9744
rect 6891 8952 6909 9736
rect 7293 8952 7311 9736
rect 6891 5992 7311 8952
rect 6891 5928 6909 5992
rect 6973 5928 6989 5992
rect 7053 5928 7069 5992
rect 7133 5928 7149 5992
rect 7213 5928 7229 5992
rect 7293 5928 7311 5992
rect 6891 4904 7311 5928
rect 6891 4840 6909 4904
rect 6973 4840 6989 4904
rect 7053 4840 7069 4904
rect 7133 4840 7149 4904
rect 7213 4840 7229 4904
rect 7293 4840 7311 4904
rect 6891 3816 7311 4840
rect 6891 3752 6909 3816
rect 6973 3752 6989 3816
rect 7053 3752 7069 3816
rect 7133 3752 7149 3816
rect 7213 3752 7229 3816
rect 7293 3752 7311 3816
rect 6891 792 7311 3752
rect 6891 8 6909 792
rect 7293 8 7311 792
rect 6891 0 7311 8
rect 7856 8596 8277 9744
rect 11384 9736 12184 9744
rect 11384 8952 11392 9736
rect 12176 8952 12184 9736
rect 7856 7812 7874 8596
rect 8258 7812 8277 8596
rect 7856 6536 8277 7812
rect 7856 6472 7874 6536
rect 7938 6472 7954 6536
rect 8018 6472 8034 6536
rect 8098 6472 8114 6536
rect 8178 6472 8194 6536
rect 8258 6472 8277 6536
rect 7856 5448 8277 6472
rect 7856 5384 7874 5448
rect 7938 5384 7954 5448
rect 8018 5384 8034 5448
rect 8098 5384 8114 5448
rect 8178 5384 8194 5448
rect 8258 5384 8277 5448
rect 7856 4360 8277 5384
rect 7856 4296 7874 4360
rect 7938 4296 7954 4360
rect 8018 4296 8034 4360
rect 8098 4296 8114 4360
rect 8178 4296 8194 4360
rect 8258 4296 8277 4360
rect 7856 3272 8277 4296
rect 7856 3208 7874 3272
rect 7938 3208 7954 3272
rect 8018 3208 8034 3272
rect 8098 3208 8114 3272
rect 8178 3208 8194 3272
rect 8258 3208 8277 3272
rect 7856 1932 8277 3208
rect 7856 1148 7874 1932
rect 8258 1148 8277 1932
rect 7856 0 8277 1148
rect 10244 8596 11044 8604
rect 10244 7812 10252 8596
rect 11036 7812 11044 8596
rect 10244 1932 11044 7812
rect 10244 1148 10252 1932
rect 11036 1148 11044 1932
rect 10244 1140 11044 1148
rect 11384 792 12184 8952
rect 11384 8 11392 792
rect 12176 8 12184 792
rect 11384 0 12184 8
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1626450099
transform -1 0 8944 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1626450099
transform 1 0 8576 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_54
timestamp 1626450099
transform 1 0 8208 0 1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1626450099
transform 1 0 7932 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_42
timestamp 1626450099
transform 1 0 7104 0 1 5960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_50
timestamp 1626450099
transform 1 0 7840 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18
timestamp 1626450099
transform 1 0 5908 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_28
timestamp 1626450099
transform 1 0 5816 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1626450099
transform 1 0 6000 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1626450099
transform 1 0 5448 0 1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1626450099
transform 1 0 3240 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1626450099
transform 1 0 3516 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1626450099
transform -1 0 4344 0 1 5960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1626450099
transform 1 0 3792 0 1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_12
timestamp 1626450099
transform 1 0 4344 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1626450099
transform -1 0 8944 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1626450099
transform 1 0 8484 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1626450099
transform 1 0 8116 0 -1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1626450099
transform 1 0 8576 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1626450099
transform -1 0 8116 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1626450099
transform 1 0 7012 0 -1 5960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp 1626450099
transform 1 0 7748 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  x11
timestamp 1626450099
transform 1 0 6644 0 -1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_27
timestamp 1626450099
transform 1 0 5724 0 -1 5960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1626450099
transform 1 0 6460 0 -1 5960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1626450099
transform 1 0 4620 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1626450099
transform 1 0 3240 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1626450099
transform 1 0 3516 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1626450099
transform -1 0 8944 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1626450099
transform 1 0 8116 0 1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_55
timestamp 1626450099
transform 1 0 8300 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  x10
timestamp 1626450099
transform 1 0 7380 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_41
timestamp 1626450099
transform 1 0 7012 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_49
timestamp 1626450099
transform 1 0 7748 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_1  x8
timestamp 1626450099
transform 1 0 6368 0 1 4872
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16
timestamp 1626450099
transform 1 0 5908 0 1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1626450099
transform 1 0 6000 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x15_A
timestamp 1626450099
transform -1 0 5540 0 1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_20
timestamp 1626450099
transform 1 0 5080 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1626450099
transform 1 0 5540 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1626450099
transform 1 0 3240 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1626450099
transform -1 0 3792 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1626450099
transform -1 0 4344 0 1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1626450099
transform 1 0 3792 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_12
timestamp 1626450099
transform 1 0 4344 0 1 4872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1626450099
transform -1 0 8944 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1626450099
transform 1 0 8484 0 -1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1626450099
transform 1 0 8392 0 -1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_58
timestamp 1626450099
transform 1 0 8576 0 -1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__a221oi_1  x7
timestamp 1626450099
transform 1 0 7196 0 -1 4872
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1626450099
transform 1 0 6828 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_50
timestamp 1626450099
transform 1 0 7840 0 -1 4872
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_1  x6
timestamp 1626450099
transform 1 0 6184 0 -1 4872
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_28
timestamp 1626450099
transform 1 0 5816 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  x15
timestamp 1626450099
transform 1 0 5540 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x6_B1
timestamp 1626450099
transform 1 0 4988 0 -1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1626450099
transform 1 0 4620 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_21
timestamp 1626450099
transform 1 0 5172 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1626450099
transform 1 0 3240 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1626450099
transform 1 0 3516 0 -1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1626450099
transform -1 0 8944 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1626450099
transform -1 0 8944 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1626450099
transform 1 0 8576 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1626450099
transform 1 0 8208 0 -1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_56
timestamp 1626450099
transform 1 0 8392 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1626450099
transform 1 0 7380 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1626450099
transform -1 0 8208 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1626450099
transform -1 0 7564 0 -1 3784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44
timestamp 1626450099
transform 1 0 7288 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1626450099
transform 1 0 7564 0 -1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1626450099
transform 1 0 7012 0 1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1626450099
transform 1 0 7656 0 1 3784
box -38 -48 774 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1626450099
transform 1 0 6460 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  x9
timestamp 1626450099
transform 1 0 6368 0 1 3784
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12
timestamp 1626450099
transform 1 0 5908 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14
timestamp 1626450099
transform 1 0 5908 0 1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1626450099
transform 1 0 5724 0 -1 3784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1626450099
transform 1 0 6000 0 -1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34
timestamp 1626450099
transform 1 0 6368 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38
timestamp 1626450099
transform 1 0 6736 0 -1 3784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1626450099
transform 1 0 6000 0 1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x9_B1
timestamp 1626450099
transform 1 0 5356 0 1 3784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1626450099
transform 1 0 4620 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1626450099
transform 1 0 4620 0 1 3784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_25
timestamp 1626450099
transform 1 0 5540 0 1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1626450099
transform 1 0 3240 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1626450099
transform 1 0 3240 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1626450099
transform 1 0 3516 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1626450099
transform 1 0 3516 0 1 3784
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 9336 4954 10136 5178 4 INN
port 1 nsew
rlabel metal2 s 9336 2286 10136 2510 4 INP
port 2 nsew
rlabel metal2 s 9336 7622 10136 7846 4 Q
port 3 nsew
rlabel metal2 s 2136 7622 2936 8560 4 VDD
port 4 nsew
rlabel metal2 s 20 4954 2936 5178 4 VSS
port 5 nsew
rlabel metal2 s 2136 2286 2936 2510 4 clk
port 6 nsew
rlabel metal3 s 1140 7804 11044 8604 4 vccd2
port 7 nsew
rlabel metal3 s 1140 1140 11044 1940 4 vccd2
port 7 nsew
rlabel metal3 s 0 8944 12184 9744 4 vssd2
port 8 nsew
rlabel metal3 s 0 0 12184 800 4 vssd2
port 8 nsew
rlabel metal4 s 7857 0 8277 9744 4 vccd2
port 7 nsew
rlabel metal4 s 5926 0 6346 9744 4 vccd2
port 7 nsew
rlabel metal4 s 3995 0 4415 9744 4 vccd2
port 7 nsew
rlabel metal4 s 10244 1140 11044 8604 4 vccd2
port 7 nsew
rlabel metal4 s 1140 1140 1940 8604 4 vccd2
port 7 nsew
rlabel metal4 s 11384 0 12184 9744 4 vssd2
port 8 nsew
rlabel metal4 s 6891 0 7311 9744 4 vssd2
port 8 nsew
rlabel metal4 s 4961 0 5381 9744 4 vssd2
port 8 nsew
rlabel metal4 s 0 0 800 9744 4 vssd2
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 12184 9744
string GDS_FILE gds/adc_wrapper.gds
string GDS_END 507114
string GDS_START 360724
<< end >>
