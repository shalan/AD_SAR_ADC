magic
tech sky130A
magscale 1 2
timestamp 1626378698
<< viali >>
rect 8145 6385 8179 6419
rect 3545 6181 3579 6215
rect 4189 6181 4223 6215
rect 7961 6181 7995 6215
rect 3729 6045 3763 6079
rect 6673 5705 6707 5739
rect 8053 5705 8087 5739
rect 6949 5637 6983 5671
rect 6765 5569 6799 5603
rect 7869 5569 7903 5603
rect 6857 5501 6891 5535
rect 7593 5297 7627 5331
rect 3545 5093 3579 5127
rect 4189 5093 4223 5127
rect 6397 5093 6431 5127
rect 6489 5093 6523 5127
rect 6627 5093 6661 5127
rect 6765 5093 6799 5127
rect 6857 5093 6891 5127
rect 7409 5093 7443 5127
rect 7501 5093 7535 5127
rect 7685 5025 7719 5059
rect 8237 5025 8271 5059
rect 3729 4957 3763 4991
rect 5477 4957 5511 4991
rect 6581 4957 6615 4991
rect 5707 4753 5741 4787
rect 7501 4685 7535 4719
rect 5604 4617 5638 4651
rect 6213 4617 6247 4651
rect 6397 4617 6431 4651
rect 6489 4617 6523 4651
rect 6765 4617 6799 4651
rect 7225 4617 7259 4651
rect 7317 4617 7351 4651
rect 7593 4617 7627 4651
rect 7685 4617 7719 4651
rect 6673 4481 6707 4515
rect 7225 4481 7259 4515
rect 5109 4413 5143 4447
rect 6581 4413 6615 4447
rect 6857 4209 6891 4243
rect 7547 4209 7581 4243
rect 6765 4141 6799 4175
rect 6397 4005 6431 4039
rect 6581 4005 6615 4039
rect 6673 4005 6707 4039
rect 6949 4005 6983 4039
rect 7444 4005 7478 4039
rect 5385 3869 5419 3903
rect 6627 3665 6661 3699
rect 7961 3665 7995 3699
rect 6524 3529 6558 3563
rect 7501 3529 7535 3563
rect 8145 3529 8179 3563
<< metal1 >>
rect 3240 6530 8944 6552
rect 3240 6478 4019 6530
rect 4071 6478 4083 6530
rect 4135 6478 4147 6530
rect 4199 6478 4211 6530
rect 4263 6478 4275 6530
rect 4327 6478 4339 6530
rect 4391 6478 5950 6530
rect 6002 6478 6014 6530
rect 6066 6478 6078 6530
rect 6130 6478 6142 6530
rect 6194 6478 6206 6530
rect 6258 6478 6270 6530
rect 6322 6478 7880 6530
rect 7932 6478 7944 6530
rect 7996 6478 8008 6530
rect 8060 6478 8072 6530
rect 8124 6478 8136 6530
rect 8188 6478 8200 6530
rect 8252 6478 8944 6530
rect 3240 6456 8944 6478
rect 8133 6419 8191 6425
rect 8133 6385 8145 6419
rect 8179 6416 8191 6419
rect 9142 6416 9148 6428
rect 8179 6388 9148 6416
rect 8179 6385 8191 6388
rect 8133 6379 8191 6385
rect 9142 6376 9148 6388
rect 9200 6376 9206 6428
rect 3162 6172 3168 6224
rect 3220 6212 3226 6224
rect 3533 6215 3591 6221
rect 3533 6212 3545 6215
rect 3220 6184 3545 6212
rect 3220 6172 3226 6184
rect 3533 6181 3545 6184
rect 3579 6212 3591 6215
rect 4177 6215 4235 6221
rect 4177 6212 4189 6215
rect 3579 6184 4189 6212
rect 3579 6181 3591 6184
rect 3533 6175 3591 6181
rect 4177 6181 4189 6184
rect 4223 6181 4235 6215
rect 4177 6175 4235 6181
rect 7578 6172 7584 6224
rect 7636 6212 7642 6224
rect 7949 6215 8007 6221
rect 7949 6212 7961 6215
rect 7636 6184 7961 6212
rect 7636 6172 7642 6184
rect 7949 6181 7961 6184
rect 7995 6181 8007 6215
rect 7949 6175 8007 6181
rect 3717 6079 3775 6085
rect 3717 6045 3729 6079
rect 3763 6076 3775 6079
rect 6658 6076 6664 6088
rect 3763 6048 6664 6076
rect 3763 6045 3775 6048
rect 3717 6039 3775 6045
rect 6658 6036 6664 6048
rect 6716 6036 6722 6088
rect 3240 5986 8944 6008
rect 3240 5934 4984 5986
rect 5036 5934 5048 5986
rect 5100 5934 5112 5986
rect 5164 5934 5176 5986
rect 5228 5934 5240 5986
rect 5292 5934 5304 5986
rect 5356 5934 6915 5986
rect 6967 5934 6979 5986
rect 7031 5934 7043 5986
rect 7095 5934 7107 5986
rect 7159 5934 7171 5986
rect 7223 5934 7235 5986
rect 7287 5934 8944 5986
rect 3240 5912 8944 5934
rect 6566 5696 6572 5748
rect 6624 5736 6630 5748
rect 6661 5739 6719 5745
rect 6661 5736 6673 5739
rect 6624 5708 6673 5736
rect 6624 5696 6630 5708
rect 6661 5705 6673 5708
rect 6707 5705 6719 5739
rect 6661 5699 6719 5705
rect 8041 5739 8099 5745
rect 8041 5705 8053 5739
rect 8087 5736 8099 5739
rect 8314 5736 8320 5748
rect 8087 5708 8320 5736
rect 8087 5705 8099 5708
rect 8041 5699 8099 5705
rect 8314 5696 8320 5708
rect 8372 5696 8378 5748
rect 6937 5671 6995 5677
rect 6937 5637 6949 5671
rect 6983 5668 6995 5671
rect 7578 5668 7584 5680
rect 6983 5640 7584 5668
rect 6983 5637 6995 5640
rect 6937 5631 6995 5637
rect 7578 5628 7584 5640
rect 7636 5628 7642 5680
rect 6750 5600 6756 5612
rect 6711 5572 6756 5600
rect 6750 5560 6756 5572
rect 6808 5560 6814 5612
rect 7026 5560 7032 5612
rect 7084 5600 7090 5612
rect 7857 5603 7915 5609
rect 7857 5600 7869 5603
rect 7084 5572 7869 5600
rect 7084 5560 7090 5572
rect 7857 5569 7869 5572
rect 7903 5569 7915 5603
rect 7857 5563 7915 5569
rect 6845 5535 6903 5541
rect 6845 5501 6857 5535
rect 6891 5532 6903 5535
rect 7394 5532 7400 5544
rect 6891 5504 7400 5532
rect 6891 5501 6903 5504
rect 6845 5495 6903 5501
rect 7394 5492 7400 5504
rect 7452 5492 7458 5544
rect 3240 5442 8944 5464
rect 3240 5390 4019 5442
rect 4071 5390 4083 5442
rect 4135 5390 4147 5442
rect 4199 5390 4211 5442
rect 4263 5390 4275 5442
rect 4327 5390 4339 5442
rect 4391 5390 5950 5442
rect 6002 5390 6014 5442
rect 6066 5390 6078 5442
rect 6130 5390 6142 5442
rect 6194 5390 6206 5442
rect 6258 5390 6270 5442
rect 6322 5390 7880 5442
rect 7932 5390 7944 5442
rect 7996 5390 8008 5442
rect 8060 5390 8072 5442
rect 8124 5390 8136 5442
rect 8188 5390 8200 5442
rect 8252 5390 8944 5442
rect 3240 5368 8944 5390
rect 7578 5328 7584 5340
rect 6400 5300 6796 5328
rect 7539 5300 7584 5328
rect 3162 5084 3168 5136
rect 3220 5124 3226 5136
rect 6400 5133 6428 5300
rect 6658 5260 6664 5272
rect 6492 5232 6664 5260
rect 6492 5133 6520 5232
rect 6658 5220 6664 5232
rect 6716 5220 6722 5272
rect 6768 5192 6796 5300
rect 7578 5288 7584 5300
rect 7636 5288 7642 5340
rect 6768 5164 7532 5192
rect 7504 5136 7532 5164
rect 3533 5127 3591 5133
rect 3533 5124 3545 5127
rect 3220 5096 3545 5124
rect 3220 5084 3226 5096
rect 3533 5093 3545 5096
rect 3579 5124 3591 5127
rect 4177 5127 4235 5133
rect 4177 5124 4189 5127
rect 3579 5096 4189 5124
rect 3579 5093 3591 5096
rect 3533 5087 3591 5093
rect 4177 5093 4189 5096
rect 4223 5093 4235 5127
rect 4177 5087 4235 5093
rect 6385 5127 6443 5133
rect 6385 5093 6397 5127
rect 6431 5093 6443 5127
rect 6385 5087 6443 5093
rect 6477 5127 6535 5133
rect 6477 5093 6489 5127
rect 6523 5093 6535 5127
rect 6477 5087 6535 5093
rect 6615 5127 6673 5133
rect 6615 5093 6627 5127
rect 6661 5093 6673 5127
rect 6615 5087 6673 5093
rect 6753 5127 6811 5133
rect 6753 5093 6765 5127
rect 6799 5124 6811 5127
rect 6845 5127 6903 5133
rect 6845 5124 6857 5127
rect 6799 5096 6857 5124
rect 6799 5093 6811 5096
rect 6753 5087 6811 5093
rect 6845 5093 6857 5096
rect 6891 5124 6903 5127
rect 7026 5124 7032 5136
rect 6891 5096 7032 5124
rect 6891 5093 6903 5096
rect 6845 5087 6903 5093
rect 6630 5056 6658 5087
rect 7026 5084 7032 5096
rect 7084 5084 7090 5136
rect 7394 5124 7400 5136
rect 7355 5096 7400 5124
rect 7394 5084 7400 5096
rect 7452 5084 7458 5136
rect 7486 5084 7492 5136
rect 7544 5124 7550 5136
rect 7544 5096 7589 5124
rect 7544 5084 7550 5096
rect 6400 5028 6658 5056
rect 7044 5056 7072 5084
rect 7302 5056 7308 5068
rect 7044 5028 7308 5056
rect 6400 5000 6428 5028
rect 7302 5016 7308 5028
rect 7360 5016 7366 5068
rect 7670 5056 7676 5068
rect 7631 5028 7676 5056
rect 7670 5016 7676 5028
rect 7728 5016 7734 5068
rect 8225 5059 8283 5065
rect 8225 5025 8237 5059
rect 8271 5056 8283 5059
rect 8314 5056 8320 5068
rect 8271 5028 8320 5056
rect 8271 5025 8283 5028
rect 8225 5019 8283 5025
rect 8314 5016 8320 5028
rect 8372 5056 8378 5068
rect 9142 5056 9148 5068
rect 8372 5028 9148 5056
rect 8372 5016 8378 5028
rect 9142 5016 9148 5028
rect 9200 5016 9206 5068
rect 3714 4988 3720 5000
rect 3675 4960 3720 4988
rect 3714 4948 3720 4960
rect 3772 4948 3778 5000
rect 5462 4988 5468 5000
rect 5423 4960 5468 4988
rect 5462 4948 5468 4960
rect 5520 4948 5526 5000
rect 6382 4948 6388 5000
rect 6440 4948 6446 5000
rect 6566 4988 6572 5000
rect 6527 4960 6572 4988
rect 6566 4948 6572 4960
rect 6624 4948 6630 5000
rect 6658 4948 6664 5000
rect 6716 4988 6722 5000
rect 7394 4988 7400 5000
rect 6716 4960 7400 4988
rect 6716 4948 6722 4960
rect 7394 4948 7400 4960
rect 7452 4948 7458 5000
rect 3240 4898 8944 4920
rect 3240 4846 4984 4898
rect 5036 4846 5048 4898
rect 5100 4846 5112 4898
rect 5164 4846 5176 4898
rect 5228 4846 5240 4898
rect 5292 4846 5304 4898
rect 5356 4846 6915 4898
rect 6967 4846 6979 4898
rect 7031 4846 7043 4898
rect 7095 4846 7107 4898
rect 7159 4846 7171 4898
rect 7223 4846 7235 4898
rect 7287 4846 8944 4898
rect 3240 4824 8944 4846
rect 5695 4787 5753 4793
rect 5695 4753 5707 4787
rect 5741 4784 5753 4787
rect 6382 4784 6388 4796
rect 5741 4756 6388 4784
rect 5741 4753 5753 4756
rect 5695 4747 5753 4753
rect 6382 4744 6388 4756
rect 6440 4784 6446 4796
rect 6440 4756 7532 4784
rect 6440 4744 6446 4756
rect 3714 4676 3720 4728
rect 3772 4716 3778 4728
rect 3772 4688 6520 4716
rect 3772 4676 3778 4688
rect 5462 4648 5468 4660
rect 5112 4620 5468 4648
rect 5112 4456 5140 4620
rect 5462 4608 5468 4620
rect 5520 4648 5526 4660
rect 5592 4651 5650 4657
rect 5592 4648 5604 4651
rect 5520 4620 5604 4648
rect 5520 4608 5526 4620
rect 5592 4617 5604 4620
rect 5638 4648 5650 4651
rect 6201 4651 6259 4657
rect 5638 4620 6152 4648
rect 5638 4617 5650 4620
rect 5592 4611 5650 4617
rect 6124 4580 6152 4620
rect 6201 4617 6213 4651
rect 6247 4648 6259 4651
rect 6290 4648 6296 4660
rect 6247 4620 6296 4648
rect 6247 4617 6259 4620
rect 6201 4611 6259 4617
rect 6290 4608 6296 4620
rect 6348 4608 6354 4660
rect 6492 4657 6520 4688
rect 6566 4676 6572 4728
rect 6624 4716 6630 4728
rect 7504 4725 7532 4756
rect 7489 4719 7547 4725
rect 6624 4688 7256 4716
rect 6624 4676 6630 4688
rect 6385 4651 6443 4657
rect 6385 4617 6397 4651
rect 6431 4617 6443 4651
rect 6385 4611 6443 4617
rect 6477 4651 6535 4657
rect 6477 4617 6489 4651
rect 6523 4648 6535 4651
rect 6658 4648 6664 4660
rect 6523 4620 6664 4648
rect 6523 4617 6535 4620
rect 6477 4611 6535 4617
rect 6400 4580 6428 4611
rect 6658 4608 6664 4620
rect 6716 4608 6722 4660
rect 7228 4657 7256 4688
rect 7489 4685 7501 4719
rect 7535 4685 7547 4719
rect 7489 4679 7547 4685
rect 6753 4651 6811 4657
rect 6753 4617 6765 4651
rect 6799 4617 6811 4651
rect 6753 4611 6811 4617
rect 7213 4651 7271 4657
rect 7213 4617 7225 4651
rect 7259 4617 7271 4651
rect 7213 4611 7271 4617
rect 7305 4651 7363 4657
rect 7305 4617 7317 4651
rect 7351 4648 7363 4651
rect 7394 4648 7400 4660
rect 7351 4620 7400 4648
rect 7351 4617 7363 4620
rect 7305 4611 7363 4617
rect 6124 4552 6428 4580
rect 6768 4580 6796 4611
rect 7394 4608 7400 4620
rect 7452 4608 7458 4660
rect 7581 4651 7639 4657
rect 7581 4617 7593 4651
rect 7627 4648 7639 4651
rect 7673 4651 7731 4657
rect 7673 4648 7685 4651
rect 7627 4620 7685 4648
rect 7627 4617 7639 4620
rect 7581 4611 7639 4617
rect 7673 4617 7685 4620
rect 7719 4648 7731 4651
rect 7762 4648 7768 4660
rect 7719 4620 7768 4648
rect 7719 4617 7731 4620
rect 7673 4611 7731 4617
rect 7596 4580 7624 4611
rect 7762 4608 7768 4620
rect 7820 4608 7826 4660
rect 6768 4552 7624 4580
rect 6661 4515 6719 4521
rect 6661 4481 6673 4515
rect 6707 4512 6719 4515
rect 6768 4512 6796 4552
rect 6707 4484 6796 4512
rect 7213 4515 7271 4521
rect 6707 4481 6719 4484
rect 6661 4475 6719 4481
rect 7213 4481 7225 4515
rect 7259 4512 7271 4515
rect 7486 4512 7492 4524
rect 7259 4484 7492 4512
rect 7259 4481 7271 4484
rect 7213 4475 7271 4481
rect 7486 4472 7492 4484
rect 7544 4472 7550 4524
rect 5094 4444 5100 4456
rect 5055 4416 5100 4444
rect 5094 4404 5100 4416
rect 5152 4404 5158 4456
rect 6382 4404 6388 4456
rect 6440 4444 6446 4456
rect 6569 4447 6627 4453
rect 6569 4444 6581 4447
rect 6440 4416 6581 4444
rect 6440 4404 6446 4416
rect 6569 4413 6581 4416
rect 6615 4413 6627 4447
rect 6569 4407 6627 4413
rect 3240 4354 8944 4376
rect 3240 4302 4019 4354
rect 4071 4302 4083 4354
rect 4135 4302 4147 4354
rect 4199 4302 4211 4354
rect 4263 4302 4275 4354
rect 4327 4302 4339 4354
rect 4391 4302 5950 4354
rect 6002 4302 6014 4354
rect 6066 4302 6078 4354
rect 6130 4302 6142 4354
rect 6194 4302 6206 4354
rect 6258 4302 6270 4354
rect 6322 4302 7880 4354
rect 7932 4302 7944 4354
rect 7996 4302 8008 4354
rect 8060 4302 8072 4354
rect 8124 4302 8136 4354
rect 8188 4302 8200 4354
rect 8252 4302 8944 4354
rect 3240 4280 8944 4302
rect 6845 4243 6903 4249
rect 6845 4209 6857 4243
rect 6891 4240 6903 4243
rect 6934 4240 6940 4252
rect 6891 4212 6940 4240
rect 6891 4209 6903 4212
rect 6845 4203 6903 4209
rect 6934 4200 6940 4212
rect 6992 4240 6998 4252
rect 7302 4240 7308 4252
rect 6992 4212 7308 4240
rect 6992 4200 6998 4212
rect 7302 4200 7308 4212
rect 7360 4200 7366 4252
rect 7535 4243 7593 4249
rect 7535 4209 7547 4243
rect 7581 4240 7593 4243
rect 7670 4240 7676 4252
rect 7581 4212 7676 4240
rect 7581 4209 7593 4212
rect 7535 4203 7593 4209
rect 7670 4200 7676 4212
rect 7728 4200 7734 4252
rect 6474 4132 6480 4184
rect 6532 4172 6538 4184
rect 6753 4175 6811 4181
rect 6753 4172 6765 4175
rect 6532 4144 6765 4172
rect 6532 4132 6538 4144
rect 6753 4141 6765 4144
rect 6799 4172 6811 4175
rect 6799 4144 7072 4172
rect 6799 4141 6811 4144
rect 6753 4135 6811 4141
rect 6382 4036 6388 4048
rect 6343 4008 6388 4036
rect 6382 3996 6388 4008
rect 6440 3996 6446 4048
rect 6569 4039 6627 4045
rect 6569 4005 6581 4039
rect 6615 4005 6627 4039
rect 6569 3999 6627 4005
rect 5094 3928 5100 3980
rect 5152 3928 5158 3980
rect 6584 3968 6612 3999
rect 6658 3996 6664 4048
rect 6716 4036 6722 4048
rect 6934 4036 6940 4048
rect 6716 4008 6761 4036
rect 6895 4008 6940 4036
rect 6716 3996 6722 4008
rect 6934 3996 6940 4008
rect 6992 3996 6998 4048
rect 7044 4036 7072 4144
rect 7432 4039 7490 4045
rect 7432 4036 7444 4039
rect 7044 4008 7444 4036
rect 7432 4005 7444 4008
rect 7478 4005 7490 4039
rect 7432 3999 7490 4005
rect 5388 3940 6612 3968
rect 3162 3860 3168 3912
rect 3220 3900 3226 3912
rect 5112 3900 5140 3928
rect 5388 3909 5416 3940
rect 5373 3903 5431 3909
rect 5373 3900 5385 3903
rect 3220 3872 5385 3900
rect 3220 3860 3226 3872
rect 5373 3869 5385 3872
rect 5419 3869 5431 3903
rect 5373 3863 5431 3869
rect 3240 3810 8944 3832
rect 3240 3758 4984 3810
rect 5036 3758 5048 3810
rect 5100 3758 5112 3810
rect 5164 3758 5176 3810
rect 5228 3758 5240 3810
rect 5292 3758 5304 3810
rect 5356 3758 6915 3810
rect 6967 3758 6979 3810
rect 7031 3758 7043 3810
rect 7095 3758 7107 3810
rect 7159 3758 7171 3810
rect 7223 3758 7235 3810
rect 7287 3758 8944 3810
rect 3240 3736 8944 3758
rect 6615 3699 6673 3705
rect 6615 3665 6627 3699
rect 6661 3696 6673 3699
rect 6750 3696 6756 3708
rect 6661 3668 6756 3696
rect 6661 3665 6673 3668
rect 6615 3659 6673 3665
rect 6750 3656 6756 3668
rect 6808 3656 6814 3708
rect 7762 3656 7768 3708
rect 7820 3696 7826 3708
rect 7949 3699 8007 3705
rect 7949 3696 7961 3699
rect 7820 3668 7961 3696
rect 7820 3656 7826 3668
rect 7949 3665 7961 3668
rect 7995 3665 8007 3699
rect 7949 3659 8007 3665
rect 6382 3520 6388 3572
rect 6440 3560 6446 3572
rect 6512 3563 6570 3569
rect 6512 3560 6524 3563
rect 6440 3532 6524 3560
rect 6440 3520 6446 3532
rect 6512 3529 6524 3532
rect 6558 3529 6570 3563
rect 6512 3523 6570 3529
rect 7489 3563 7547 3569
rect 7489 3529 7501 3563
rect 7535 3560 7547 3563
rect 8133 3563 8191 3569
rect 8133 3560 8145 3563
rect 7535 3532 8145 3560
rect 7535 3529 7547 3532
rect 7489 3523 7547 3529
rect 8133 3529 8145 3532
rect 8179 3560 8191 3563
rect 9142 3560 9148 3572
rect 8179 3532 9148 3560
rect 8179 3529 8191 3532
rect 8133 3523 8191 3529
rect 9142 3520 9148 3532
rect 9200 3520 9206 3572
rect 3240 3266 8944 3288
rect 3240 3214 4019 3266
rect 4071 3214 4083 3266
rect 4135 3214 4147 3266
rect 4199 3214 4211 3266
rect 4263 3214 4275 3266
rect 4327 3214 4339 3266
rect 4391 3214 5950 3266
rect 6002 3214 6014 3266
rect 6066 3214 6078 3266
rect 6130 3214 6142 3266
rect 6194 3214 6206 3266
rect 6258 3214 6270 3266
rect 6322 3214 7880 3266
rect 7932 3214 7944 3266
rect 7996 3214 8008 3266
rect 8060 3214 8072 3266
rect 8124 3214 8136 3266
rect 8188 3214 8200 3266
rect 8252 3214 8944 3266
rect 3240 3192 8944 3214
<< via1 >>
rect 4019 6478 4071 6530
rect 4083 6478 4135 6530
rect 4147 6478 4199 6530
rect 4211 6478 4263 6530
rect 4275 6478 4327 6530
rect 4339 6478 4391 6530
rect 5950 6478 6002 6530
rect 6014 6478 6066 6530
rect 6078 6478 6130 6530
rect 6142 6478 6194 6530
rect 6206 6478 6258 6530
rect 6270 6478 6322 6530
rect 7880 6478 7932 6530
rect 7944 6478 7996 6530
rect 8008 6478 8060 6530
rect 8072 6478 8124 6530
rect 8136 6478 8188 6530
rect 8200 6478 8252 6530
rect 9148 6376 9200 6428
rect 3168 6172 3220 6224
rect 7584 6172 7636 6224
rect 6664 6036 6716 6088
rect 4984 5934 5036 5986
rect 5048 5934 5100 5986
rect 5112 5934 5164 5986
rect 5176 5934 5228 5986
rect 5240 5934 5292 5986
rect 5304 5934 5356 5986
rect 6915 5934 6967 5986
rect 6979 5934 7031 5986
rect 7043 5934 7095 5986
rect 7107 5934 7159 5986
rect 7171 5934 7223 5986
rect 7235 5934 7287 5986
rect 6572 5696 6624 5748
rect 8320 5696 8372 5748
rect 7584 5628 7636 5680
rect 6756 5603 6808 5612
rect 6756 5569 6765 5603
rect 6765 5569 6799 5603
rect 6799 5569 6808 5603
rect 6756 5560 6808 5569
rect 7032 5560 7084 5612
rect 7400 5492 7452 5544
rect 4019 5390 4071 5442
rect 4083 5390 4135 5442
rect 4147 5390 4199 5442
rect 4211 5390 4263 5442
rect 4275 5390 4327 5442
rect 4339 5390 4391 5442
rect 5950 5390 6002 5442
rect 6014 5390 6066 5442
rect 6078 5390 6130 5442
rect 6142 5390 6194 5442
rect 6206 5390 6258 5442
rect 6270 5390 6322 5442
rect 7880 5390 7932 5442
rect 7944 5390 7996 5442
rect 8008 5390 8060 5442
rect 8072 5390 8124 5442
rect 8136 5390 8188 5442
rect 8200 5390 8252 5442
rect 7584 5331 7636 5340
rect 3168 5084 3220 5136
rect 6664 5220 6716 5272
rect 7584 5297 7593 5331
rect 7593 5297 7627 5331
rect 7627 5297 7636 5331
rect 7584 5288 7636 5297
rect 7032 5084 7084 5136
rect 7400 5127 7452 5136
rect 7400 5093 7409 5127
rect 7409 5093 7443 5127
rect 7443 5093 7452 5127
rect 7400 5084 7452 5093
rect 7492 5127 7544 5136
rect 7492 5093 7501 5127
rect 7501 5093 7535 5127
rect 7535 5093 7544 5127
rect 7492 5084 7544 5093
rect 7308 5016 7360 5068
rect 7676 5059 7728 5068
rect 7676 5025 7685 5059
rect 7685 5025 7719 5059
rect 7719 5025 7728 5059
rect 7676 5016 7728 5025
rect 8320 5016 8372 5068
rect 9148 5016 9200 5068
rect 3720 4991 3772 5000
rect 3720 4957 3729 4991
rect 3729 4957 3763 4991
rect 3763 4957 3772 4991
rect 3720 4948 3772 4957
rect 5468 4991 5520 5000
rect 5468 4957 5477 4991
rect 5477 4957 5511 4991
rect 5511 4957 5520 4991
rect 5468 4948 5520 4957
rect 6388 4948 6440 5000
rect 6572 4991 6624 5000
rect 6572 4957 6581 4991
rect 6581 4957 6615 4991
rect 6615 4957 6624 4991
rect 6572 4948 6624 4957
rect 6664 4948 6716 5000
rect 7400 4948 7452 5000
rect 4984 4846 5036 4898
rect 5048 4846 5100 4898
rect 5112 4846 5164 4898
rect 5176 4846 5228 4898
rect 5240 4846 5292 4898
rect 5304 4846 5356 4898
rect 6915 4846 6967 4898
rect 6979 4846 7031 4898
rect 7043 4846 7095 4898
rect 7107 4846 7159 4898
rect 7171 4846 7223 4898
rect 7235 4846 7287 4898
rect 6388 4744 6440 4796
rect 3720 4676 3772 4728
rect 5468 4608 5520 4660
rect 6296 4608 6348 4660
rect 6572 4676 6624 4728
rect 6664 4608 6716 4660
rect 7400 4608 7452 4660
rect 7768 4608 7820 4660
rect 7492 4472 7544 4524
rect 5100 4447 5152 4456
rect 5100 4413 5109 4447
rect 5109 4413 5143 4447
rect 5143 4413 5152 4447
rect 5100 4404 5152 4413
rect 6388 4404 6440 4456
rect 4019 4302 4071 4354
rect 4083 4302 4135 4354
rect 4147 4302 4199 4354
rect 4211 4302 4263 4354
rect 4275 4302 4327 4354
rect 4339 4302 4391 4354
rect 5950 4302 6002 4354
rect 6014 4302 6066 4354
rect 6078 4302 6130 4354
rect 6142 4302 6194 4354
rect 6206 4302 6258 4354
rect 6270 4302 6322 4354
rect 7880 4302 7932 4354
rect 7944 4302 7996 4354
rect 8008 4302 8060 4354
rect 8072 4302 8124 4354
rect 8136 4302 8188 4354
rect 8200 4302 8252 4354
rect 6940 4200 6992 4252
rect 7308 4200 7360 4252
rect 7676 4200 7728 4252
rect 6480 4132 6532 4184
rect 6388 4039 6440 4048
rect 6388 4005 6397 4039
rect 6397 4005 6431 4039
rect 6431 4005 6440 4039
rect 6388 3996 6440 4005
rect 5100 3928 5152 3980
rect 6664 4039 6716 4048
rect 6664 4005 6673 4039
rect 6673 4005 6707 4039
rect 6707 4005 6716 4039
rect 6940 4039 6992 4048
rect 6664 3996 6716 4005
rect 6940 4005 6949 4039
rect 6949 4005 6983 4039
rect 6983 4005 6992 4039
rect 6940 3996 6992 4005
rect 3168 3860 3220 3912
rect 4984 3758 5036 3810
rect 5048 3758 5100 3810
rect 5112 3758 5164 3810
rect 5176 3758 5228 3810
rect 5240 3758 5292 3810
rect 5304 3758 5356 3810
rect 6915 3758 6967 3810
rect 6979 3758 7031 3810
rect 7043 3758 7095 3810
rect 7107 3758 7159 3810
rect 7171 3758 7223 3810
rect 7235 3758 7287 3810
rect 6756 3656 6808 3708
rect 7768 3656 7820 3708
rect 6388 3520 6440 3572
rect 9148 3520 9200 3572
rect 4019 3214 4071 3266
rect 4083 3214 4135 3266
rect 4147 3214 4199 3266
rect 4211 3214 4263 3266
rect 4275 3214 4327 3266
rect 4339 3214 4391 3266
rect 5950 3214 6002 3266
rect 6014 3214 6066 3266
rect 6078 3214 6130 3266
rect 6142 3214 6194 3266
rect 6206 3214 6258 3266
rect 6270 3214 6322 3266
rect 7880 3214 7932 3266
rect 7944 3214 7996 3266
rect 8008 3214 8060 3266
rect 8072 3214 8124 3266
rect 8136 3214 8188 3266
rect 8200 3214 8252 3266
<< metal2 >>
rect 2136 7748 2936 7846
rect 9336 7748 10136 7846
rect 2136 7720 3208 7748
rect 2136 7622 2936 7720
rect 3180 6230 3208 7720
rect 9160 7720 10136 7748
rect 4017 6532 4393 6552
rect 4073 6530 4097 6532
rect 4153 6530 4177 6532
rect 4233 6530 4257 6532
rect 4313 6530 4337 6532
rect 4073 6478 4083 6530
rect 4327 6478 4337 6530
rect 4073 6476 4097 6478
rect 4153 6476 4177 6478
rect 4233 6476 4257 6478
rect 4313 6476 4337 6478
rect 4017 6456 4393 6476
rect 5948 6532 6324 6552
rect 6004 6530 6028 6532
rect 6084 6530 6108 6532
rect 6164 6530 6188 6532
rect 6244 6530 6268 6532
rect 6004 6478 6014 6530
rect 6258 6478 6268 6530
rect 6004 6476 6028 6478
rect 6084 6476 6108 6478
rect 6164 6476 6188 6478
rect 6244 6476 6268 6478
rect 5948 6456 6324 6476
rect 7878 6532 8254 6552
rect 7934 6530 7958 6532
rect 8014 6530 8038 6532
rect 8094 6530 8118 6532
rect 8174 6530 8198 6532
rect 7934 6478 7944 6530
rect 8188 6478 8198 6530
rect 7934 6476 7958 6478
rect 8014 6476 8038 6478
rect 8094 6476 8118 6478
rect 8174 6476 8198 6478
rect 7878 6456 8254 6476
rect 9160 6434 9188 7720
rect 9336 7622 10136 7720
rect 9148 6428 9200 6434
rect 9148 6370 9200 6376
rect 3168 6224 3220 6230
rect 3168 6166 3220 6172
rect 7584 6224 7636 6230
rect 7584 6166 7636 6172
rect 6664 6088 6716 6094
rect 6664 6030 6716 6036
rect 4982 5988 5358 6008
rect 5038 5986 5062 5988
rect 5118 5986 5142 5988
rect 5198 5986 5222 5988
rect 5278 5986 5302 5988
rect 5038 5934 5048 5986
rect 5292 5934 5302 5986
rect 5038 5932 5062 5934
rect 5118 5932 5142 5934
rect 5198 5932 5222 5934
rect 5278 5932 5302 5934
rect 4982 5912 5358 5932
rect 6572 5748 6624 5754
rect 6572 5690 6624 5696
rect 4017 5444 4393 5464
rect 4073 5442 4097 5444
rect 4153 5442 4177 5444
rect 4233 5442 4257 5444
rect 4313 5442 4337 5444
rect 4073 5390 4083 5442
rect 4327 5390 4337 5442
rect 4073 5388 4097 5390
rect 4153 5388 4177 5390
rect 4233 5388 4257 5390
rect 4313 5388 4337 5390
rect 4017 5368 4393 5388
rect 5948 5444 6324 5464
rect 6004 5442 6028 5444
rect 6084 5442 6108 5444
rect 6164 5442 6188 5444
rect 6244 5442 6268 5444
rect 6004 5390 6014 5442
rect 6258 5390 6268 5442
rect 6004 5388 6028 5390
rect 6084 5388 6108 5390
rect 6164 5388 6188 5390
rect 6244 5388 6268 5390
rect 5948 5368 6324 5388
rect 2136 5080 2936 5178
rect 3168 5136 3220 5142
rect 3168 5080 3220 5084
rect 2136 5078 3220 5080
rect 2136 5052 3208 5078
rect 2136 4954 2936 5052
rect 6584 5006 6612 5690
rect 6676 5278 6704 6030
rect 6913 5988 7289 6008
rect 6969 5986 6993 5988
rect 7049 5986 7073 5988
rect 7129 5986 7153 5988
rect 7209 5986 7233 5988
rect 6969 5934 6979 5986
rect 7223 5934 7233 5986
rect 6969 5932 6993 5934
rect 7049 5932 7073 5934
rect 7129 5932 7153 5934
rect 7209 5932 7233 5934
rect 6913 5912 7289 5932
rect 7596 5686 7624 6166
rect 8320 5748 8372 5754
rect 8320 5690 8372 5696
rect 7584 5680 7636 5686
rect 7584 5622 7636 5628
rect 6756 5612 6808 5618
rect 6756 5554 6808 5560
rect 7032 5612 7084 5618
rect 7032 5554 7084 5560
rect 6664 5272 6716 5278
rect 6664 5214 6716 5220
rect 6676 5006 6704 5214
rect 3720 5000 3772 5006
rect 3720 4942 3772 4948
rect 5468 5000 5520 5006
rect 5468 4942 5520 4948
rect 6388 5000 6440 5006
rect 6388 4942 6440 4948
rect 6572 5000 6624 5006
rect 6572 4942 6624 4948
rect 6664 5000 6716 5006
rect 6664 4942 6716 4948
rect 3732 4734 3760 4942
rect 4982 4900 5358 4920
rect 5038 4898 5062 4900
rect 5118 4898 5142 4900
rect 5198 4898 5222 4900
rect 5278 4898 5302 4900
rect 5038 4846 5048 4898
rect 5292 4846 5302 4898
rect 5038 4844 5062 4846
rect 5118 4844 5142 4846
rect 5198 4844 5222 4846
rect 5278 4844 5302 4846
rect 4982 4824 5358 4844
rect 3720 4728 3772 4734
rect 3720 4670 3772 4676
rect 5480 4666 5508 4942
rect 6400 4802 6428 4942
rect 6388 4796 6440 4802
rect 6388 4738 6440 4744
rect 6584 4734 6612 4942
rect 6572 4728 6624 4734
rect 6572 4670 6624 4676
rect 5468 4660 5520 4666
rect 5468 4602 5520 4608
rect 6296 4660 6348 4666
rect 6296 4602 6348 4608
rect 6664 4660 6716 4666
rect 6664 4602 6716 4608
rect 6308 4546 6336 4602
rect 6308 4518 6520 4546
rect 5100 4456 5152 4462
rect 5100 4398 5152 4404
rect 6388 4456 6440 4462
rect 6388 4398 6440 4404
rect 4017 4356 4393 4376
rect 4073 4354 4097 4356
rect 4153 4354 4177 4356
rect 4233 4354 4257 4356
rect 4313 4354 4337 4356
rect 4073 4302 4083 4354
rect 4327 4302 4337 4354
rect 4073 4300 4097 4302
rect 4153 4300 4177 4302
rect 4233 4300 4257 4302
rect 4313 4300 4337 4302
rect 4017 4280 4393 4300
rect 5112 3986 5140 4398
rect 5948 4356 6324 4376
rect 6004 4354 6028 4356
rect 6084 4354 6108 4356
rect 6164 4354 6188 4356
rect 6244 4354 6268 4356
rect 6004 4302 6014 4354
rect 6258 4302 6268 4354
rect 6004 4300 6028 4302
rect 6084 4300 6108 4302
rect 6164 4300 6188 4302
rect 6244 4300 6268 4302
rect 5948 4280 6324 4300
rect 6400 4054 6428 4398
rect 6492 4190 6520 4518
rect 6480 4184 6532 4190
rect 6480 4126 6532 4132
rect 6676 4054 6704 4602
rect 6388 4048 6440 4054
rect 6388 3990 6440 3996
rect 6664 4048 6716 4054
rect 6664 3990 6716 3996
rect 5100 3980 5152 3986
rect 5100 3922 5152 3928
rect 3168 3912 3220 3918
rect 3168 3854 3220 3860
rect 2136 2412 2936 2510
rect 3180 2412 3208 3854
rect 4982 3812 5358 3832
rect 5038 3810 5062 3812
rect 5118 3810 5142 3812
rect 5198 3810 5222 3812
rect 5278 3810 5302 3812
rect 5038 3758 5048 3810
rect 5292 3758 5302 3810
rect 5038 3756 5062 3758
rect 5118 3756 5142 3758
rect 5198 3756 5222 3758
rect 5278 3756 5302 3758
rect 4982 3736 5358 3756
rect 6400 3578 6428 3990
rect 6768 3714 6796 5554
rect 7044 5142 7072 5554
rect 7400 5544 7452 5550
rect 7400 5486 7452 5492
rect 7412 5142 7440 5486
rect 7596 5346 7624 5622
rect 7878 5444 8254 5464
rect 7934 5442 7958 5444
rect 8014 5442 8038 5444
rect 8094 5442 8118 5444
rect 8174 5442 8198 5444
rect 7934 5390 7944 5442
rect 8188 5390 8198 5442
rect 7934 5388 7958 5390
rect 8014 5388 8038 5390
rect 8094 5388 8118 5390
rect 8174 5388 8198 5390
rect 7878 5368 8254 5388
rect 7584 5340 7636 5346
rect 7584 5282 7636 5288
rect 7032 5136 7084 5142
rect 7032 5078 7084 5084
rect 7400 5136 7452 5142
rect 7400 5078 7452 5084
rect 7492 5136 7544 5142
rect 7492 5078 7544 5084
rect 7308 5068 7360 5074
rect 7308 5010 7360 5016
rect 6913 4900 7289 4920
rect 6969 4898 6993 4900
rect 7049 4898 7073 4900
rect 7129 4898 7153 4900
rect 7209 4898 7233 4900
rect 6969 4846 6979 4898
rect 7223 4846 7233 4898
rect 6969 4844 6993 4846
rect 7049 4844 7073 4846
rect 7129 4844 7153 4846
rect 7209 4844 7233 4846
rect 6913 4824 7289 4844
rect 7320 4258 7348 5010
rect 7400 5000 7452 5006
rect 7400 4942 7452 4948
rect 7412 4666 7440 4942
rect 7400 4660 7452 4666
rect 7400 4602 7452 4608
rect 7504 4530 7532 5078
rect 8332 5074 8360 5690
rect 9336 5080 10136 5178
rect 9160 5074 10136 5080
rect 7676 5068 7728 5074
rect 7676 5010 7728 5016
rect 8320 5068 8372 5074
rect 8320 5010 8372 5016
rect 9148 5068 10136 5074
rect 9200 5052 10136 5068
rect 9148 5010 9200 5016
rect 7492 4524 7544 4530
rect 7492 4466 7544 4472
rect 7688 4258 7716 5010
rect 9336 4954 10136 5052
rect 7768 4660 7820 4666
rect 7768 4602 7820 4608
rect 6940 4252 6992 4258
rect 6940 4194 6992 4200
rect 7308 4252 7360 4258
rect 7308 4194 7360 4200
rect 7676 4252 7728 4258
rect 7676 4194 7728 4200
rect 6952 4054 6980 4194
rect 6940 4048 6992 4054
rect 6940 3990 6992 3996
rect 6913 3812 7289 3832
rect 6969 3810 6993 3812
rect 7049 3810 7073 3812
rect 7129 3810 7153 3812
rect 7209 3810 7233 3812
rect 6969 3758 6979 3810
rect 7223 3758 7233 3810
rect 6969 3756 6993 3758
rect 7049 3756 7073 3758
rect 7129 3756 7153 3758
rect 7209 3756 7233 3758
rect 6913 3736 7289 3756
rect 7780 3714 7808 4602
rect 7878 4356 8254 4376
rect 7934 4354 7958 4356
rect 8014 4354 8038 4356
rect 8094 4354 8118 4356
rect 8174 4354 8198 4356
rect 7934 4302 7944 4354
rect 8188 4302 8198 4354
rect 7934 4300 7958 4302
rect 8014 4300 8038 4302
rect 8094 4300 8118 4302
rect 8174 4300 8198 4302
rect 7878 4280 8254 4300
rect 6756 3708 6808 3714
rect 6756 3650 6808 3656
rect 7768 3708 7820 3714
rect 7768 3650 7820 3656
rect 6388 3572 6440 3578
rect 6388 3514 6440 3520
rect 9148 3572 9200 3578
rect 9148 3514 9200 3520
rect 4017 3268 4393 3288
rect 4073 3266 4097 3268
rect 4153 3266 4177 3268
rect 4233 3266 4257 3268
rect 4313 3266 4337 3268
rect 4073 3214 4083 3266
rect 4327 3214 4337 3266
rect 4073 3212 4097 3214
rect 4153 3212 4177 3214
rect 4233 3212 4257 3214
rect 4313 3212 4337 3214
rect 4017 3192 4393 3212
rect 5948 3268 6324 3288
rect 6004 3266 6028 3268
rect 6084 3266 6108 3268
rect 6164 3266 6188 3268
rect 6244 3266 6268 3268
rect 6004 3214 6014 3266
rect 6258 3214 6268 3266
rect 6004 3212 6028 3214
rect 6084 3212 6108 3214
rect 6164 3212 6188 3214
rect 6244 3212 6268 3214
rect 5948 3192 6324 3212
rect 7878 3268 8254 3288
rect 7934 3266 7958 3268
rect 8014 3266 8038 3268
rect 8094 3266 8118 3268
rect 8174 3266 8198 3268
rect 7934 3214 7944 3266
rect 8188 3214 8198 3266
rect 7934 3212 7958 3214
rect 8014 3212 8038 3214
rect 8094 3212 8118 3214
rect 8174 3212 8198 3214
rect 7878 3192 8254 3212
rect 2136 2384 3208 2412
rect 9160 2412 9188 3514
rect 9336 2412 10136 2510
rect 9160 2384 10136 2412
rect 2136 2286 2936 2384
rect 9336 2286 10136 2384
<< via2 >>
rect 4017 6530 4073 6532
rect 4097 6530 4153 6532
rect 4177 6530 4233 6532
rect 4257 6530 4313 6532
rect 4337 6530 4393 6532
rect 4017 6478 4019 6530
rect 4019 6478 4071 6530
rect 4071 6478 4073 6530
rect 4097 6478 4135 6530
rect 4135 6478 4147 6530
rect 4147 6478 4153 6530
rect 4177 6478 4199 6530
rect 4199 6478 4211 6530
rect 4211 6478 4233 6530
rect 4257 6478 4263 6530
rect 4263 6478 4275 6530
rect 4275 6478 4313 6530
rect 4337 6478 4339 6530
rect 4339 6478 4391 6530
rect 4391 6478 4393 6530
rect 4017 6476 4073 6478
rect 4097 6476 4153 6478
rect 4177 6476 4233 6478
rect 4257 6476 4313 6478
rect 4337 6476 4393 6478
rect 5948 6530 6004 6532
rect 6028 6530 6084 6532
rect 6108 6530 6164 6532
rect 6188 6530 6244 6532
rect 6268 6530 6324 6532
rect 5948 6478 5950 6530
rect 5950 6478 6002 6530
rect 6002 6478 6004 6530
rect 6028 6478 6066 6530
rect 6066 6478 6078 6530
rect 6078 6478 6084 6530
rect 6108 6478 6130 6530
rect 6130 6478 6142 6530
rect 6142 6478 6164 6530
rect 6188 6478 6194 6530
rect 6194 6478 6206 6530
rect 6206 6478 6244 6530
rect 6268 6478 6270 6530
rect 6270 6478 6322 6530
rect 6322 6478 6324 6530
rect 5948 6476 6004 6478
rect 6028 6476 6084 6478
rect 6108 6476 6164 6478
rect 6188 6476 6244 6478
rect 6268 6476 6324 6478
rect 7878 6530 7934 6532
rect 7958 6530 8014 6532
rect 8038 6530 8094 6532
rect 8118 6530 8174 6532
rect 8198 6530 8254 6532
rect 7878 6478 7880 6530
rect 7880 6478 7932 6530
rect 7932 6478 7934 6530
rect 7958 6478 7996 6530
rect 7996 6478 8008 6530
rect 8008 6478 8014 6530
rect 8038 6478 8060 6530
rect 8060 6478 8072 6530
rect 8072 6478 8094 6530
rect 8118 6478 8124 6530
rect 8124 6478 8136 6530
rect 8136 6478 8174 6530
rect 8198 6478 8200 6530
rect 8200 6478 8252 6530
rect 8252 6478 8254 6530
rect 7878 6476 7934 6478
rect 7958 6476 8014 6478
rect 8038 6476 8094 6478
rect 8118 6476 8174 6478
rect 8198 6476 8254 6478
rect 4982 5986 5038 5988
rect 5062 5986 5118 5988
rect 5142 5986 5198 5988
rect 5222 5986 5278 5988
rect 5302 5986 5358 5988
rect 4982 5934 4984 5986
rect 4984 5934 5036 5986
rect 5036 5934 5038 5986
rect 5062 5934 5100 5986
rect 5100 5934 5112 5986
rect 5112 5934 5118 5986
rect 5142 5934 5164 5986
rect 5164 5934 5176 5986
rect 5176 5934 5198 5986
rect 5222 5934 5228 5986
rect 5228 5934 5240 5986
rect 5240 5934 5278 5986
rect 5302 5934 5304 5986
rect 5304 5934 5356 5986
rect 5356 5934 5358 5986
rect 4982 5932 5038 5934
rect 5062 5932 5118 5934
rect 5142 5932 5198 5934
rect 5222 5932 5278 5934
rect 5302 5932 5358 5934
rect 4017 5442 4073 5444
rect 4097 5442 4153 5444
rect 4177 5442 4233 5444
rect 4257 5442 4313 5444
rect 4337 5442 4393 5444
rect 4017 5390 4019 5442
rect 4019 5390 4071 5442
rect 4071 5390 4073 5442
rect 4097 5390 4135 5442
rect 4135 5390 4147 5442
rect 4147 5390 4153 5442
rect 4177 5390 4199 5442
rect 4199 5390 4211 5442
rect 4211 5390 4233 5442
rect 4257 5390 4263 5442
rect 4263 5390 4275 5442
rect 4275 5390 4313 5442
rect 4337 5390 4339 5442
rect 4339 5390 4391 5442
rect 4391 5390 4393 5442
rect 4017 5388 4073 5390
rect 4097 5388 4153 5390
rect 4177 5388 4233 5390
rect 4257 5388 4313 5390
rect 4337 5388 4393 5390
rect 5948 5442 6004 5444
rect 6028 5442 6084 5444
rect 6108 5442 6164 5444
rect 6188 5442 6244 5444
rect 6268 5442 6324 5444
rect 5948 5390 5950 5442
rect 5950 5390 6002 5442
rect 6002 5390 6004 5442
rect 6028 5390 6066 5442
rect 6066 5390 6078 5442
rect 6078 5390 6084 5442
rect 6108 5390 6130 5442
rect 6130 5390 6142 5442
rect 6142 5390 6164 5442
rect 6188 5390 6194 5442
rect 6194 5390 6206 5442
rect 6206 5390 6244 5442
rect 6268 5390 6270 5442
rect 6270 5390 6322 5442
rect 6322 5390 6324 5442
rect 5948 5388 6004 5390
rect 6028 5388 6084 5390
rect 6108 5388 6164 5390
rect 6188 5388 6244 5390
rect 6268 5388 6324 5390
rect 6913 5986 6969 5988
rect 6993 5986 7049 5988
rect 7073 5986 7129 5988
rect 7153 5986 7209 5988
rect 7233 5986 7289 5988
rect 6913 5934 6915 5986
rect 6915 5934 6967 5986
rect 6967 5934 6969 5986
rect 6993 5934 7031 5986
rect 7031 5934 7043 5986
rect 7043 5934 7049 5986
rect 7073 5934 7095 5986
rect 7095 5934 7107 5986
rect 7107 5934 7129 5986
rect 7153 5934 7159 5986
rect 7159 5934 7171 5986
rect 7171 5934 7209 5986
rect 7233 5934 7235 5986
rect 7235 5934 7287 5986
rect 7287 5934 7289 5986
rect 6913 5932 6969 5934
rect 6993 5932 7049 5934
rect 7073 5932 7129 5934
rect 7153 5932 7209 5934
rect 7233 5932 7289 5934
rect 4982 4898 5038 4900
rect 5062 4898 5118 4900
rect 5142 4898 5198 4900
rect 5222 4898 5278 4900
rect 5302 4898 5358 4900
rect 4982 4846 4984 4898
rect 4984 4846 5036 4898
rect 5036 4846 5038 4898
rect 5062 4846 5100 4898
rect 5100 4846 5112 4898
rect 5112 4846 5118 4898
rect 5142 4846 5164 4898
rect 5164 4846 5176 4898
rect 5176 4846 5198 4898
rect 5222 4846 5228 4898
rect 5228 4846 5240 4898
rect 5240 4846 5278 4898
rect 5302 4846 5304 4898
rect 5304 4846 5356 4898
rect 5356 4846 5358 4898
rect 4982 4844 5038 4846
rect 5062 4844 5118 4846
rect 5142 4844 5198 4846
rect 5222 4844 5278 4846
rect 5302 4844 5358 4846
rect 4017 4354 4073 4356
rect 4097 4354 4153 4356
rect 4177 4354 4233 4356
rect 4257 4354 4313 4356
rect 4337 4354 4393 4356
rect 4017 4302 4019 4354
rect 4019 4302 4071 4354
rect 4071 4302 4073 4354
rect 4097 4302 4135 4354
rect 4135 4302 4147 4354
rect 4147 4302 4153 4354
rect 4177 4302 4199 4354
rect 4199 4302 4211 4354
rect 4211 4302 4233 4354
rect 4257 4302 4263 4354
rect 4263 4302 4275 4354
rect 4275 4302 4313 4354
rect 4337 4302 4339 4354
rect 4339 4302 4391 4354
rect 4391 4302 4393 4354
rect 4017 4300 4073 4302
rect 4097 4300 4153 4302
rect 4177 4300 4233 4302
rect 4257 4300 4313 4302
rect 4337 4300 4393 4302
rect 5948 4354 6004 4356
rect 6028 4354 6084 4356
rect 6108 4354 6164 4356
rect 6188 4354 6244 4356
rect 6268 4354 6324 4356
rect 5948 4302 5950 4354
rect 5950 4302 6002 4354
rect 6002 4302 6004 4354
rect 6028 4302 6066 4354
rect 6066 4302 6078 4354
rect 6078 4302 6084 4354
rect 6108 4302 6130 4354
rect 6130 4302 6142 4354
rect 6142 4302 6164 4354
rect 6188 4302 6194 4354
rect 6194 4302 6206 4354
rect 6206 4302 6244 4354
rect 6268 4302 6270 4354
rect 6270 4302 6322 4354
rect 6322 4302 6324 4354
rect 5948 4300 6004 4302
rect 6028 4300 6084 4302
rect 6108 4300 6164 4302
rect 6188 4300 6244 4302
rect 6268 4300 6324 4302
rect 4982 3810 5038 3812
rect 5062 3810 5118 3812
rect 5142 3810 5198 3812
rect 5222 3810 5278 3812
rect 5302 3810 5358 3812
rect 4982 3758 4984 3810
rect 4984 3758 5036 3810
rect 5036 3758 5038 3810
rect 5062 3758 5100 3810
rect 5100 3758 5112 3810
rect 5112 3758 5118 3810
rect 5142 3758 5164 3810
rect 5164 3758 5176 3810
rect 5176 3758 5198 3810
rect 5222 3758 5228 3810
rect 5228 3758 5240 3810
rect 5240 3758 5278 3810
rect 5302 3758 5304 3810
rect 5304 3758 5356 3810
rect 5356 3758 5358 3810
rect 4982 3756 5038 3758
rect 5062 3756 5118 3758
rect 5142 3756 5198 3758
rect 5222 3756 5278 3758
rect 5302 3756 5358 3758
rect 7878 5442 7934 5444
rect 7958 5442 8014 5444
rect 8038 5442 8094 5444
rect 8118 5442 8174 5444
rect 8198 5442 8254 5444
rect 7878 5390 7880 5442
rect 7880 5390 7932 5442
rect 7932 5390 7934 5442
rect 7958 5390 7996 5442
rect 7996 5390 8008 5442
rect 8008 5390 8014 5442
rect 8038 5390 8060 5442
rect 8060 5390 8072 5442
rect 8072 5390 8094 5442
rect 8118 5390 8124 5442
rect 8124 5390 8136 5442
rect 8136 5390 8174 5442
rect 8198 5390 8200 5442
rect 8200 5390 8252 5442
rect 8252 5390 8254 5442
rect 7878 5388 7934 5390
rect 7958 5388 8014 5390
rect 8038 5388 8094 5390
rect 8118 5388 8174 5390
rect 8198 5388 8254 5390
rect 6913 4898 6969 4900
rect 6993 4898 7049 4900
rect 7073 4898 7129 4900
rect 7153 4898 7209 4900
rect 7233 4898 7289 4900
rect 6913 4846 6915 4898
rect 6915 4846 6967 4898
rect 6967 4846 6969 4898
rect 6993 4846 7031 4898
rect 7031 4846 7043 4898
rect 7043 4846 7049 4898
rect 7073 4846 7095 4898
rect 7095 4846 7107 4898
rect 7107 4846 7129 4898
rect 7153 4846 7159 4898
rect 7159 4846 7171 4898
rect 7171 4846 7209 4898
rect 7233 4846 7235 4898
rect 7235 4846 7287 4898
rect 7287 4846 7289 4898
rect 6913 4844 6969 4846
rect 6993 4844 7049 4846
rect 7073 4844 7129 4846
rect 7153 4844 7209 4846
rect 7233 4844 7289 4846
rect 6913 3810 6969 3812
rect 6993 3810 7049 3812
rect 7073 3810 7129 3812
rect 7153 3810 7209 3812
rect 7233 3810 7289 3812
rect 6913 3758 6915 3810
rect 6915 3758 6967 3810
rect 6967 3758 6969 3810
rect 6993 3758 7031 3810
rect 7031 3758 7043 3810
rect 7043 3758 7049 3810
rect 7073 3758 7095 3810
rect 7095 3758 7107 3810
rect 7107 3758 7129 3810
rect 7153 3758 7159 3810
rect 7159 3758 7171 3810
rect 7171 3758 7209 3810
rect 7233 3758 7235 3810
rect 7235 3758 7287 3810
rect 7287 3758 7289 3810
rect 6913 3756 6969 3758
rect 6993 3756 7049 3758
rect 7073 3756 7129 3758
rect 7153 3756 7209 3758
rect 7233 3756 7289 3758
rect 7878 4354 7934 4356
rect 7958 4354 8014 4356
rect 8038 4354 8094 4356
rect 8118 4354 8174 4356
rect 8198 4354 8254 4356
rect 7878 4302 7880 4354
rect 7880 4302 7932 4354
rect 7932 4302 7934 4354
rect 7958 4302 7996 4354
rect 7996 4302 8008 4354
rect 8008 4302 8014 4354
rect 8038 4302 8060 4354
rect 8060 4302 8072 4354
rect 8072 4302 8094 4354
rect 8118 4302 8124 4354
rect 8124 4302 8136 4354
rect 8136 4302 8174 4354
rect 8198 4302 8200 4354
rect 8200 4302 8252 4354
rect 8252 4302 8254 4354
rect 7878 4300 7934 4302
rect 7958 4300 8014 4302
rect 8038 4300 8094 4302
rect 8118 4300 8174 4302
rect 8198 4300 8254 4302
rect 4017 3266 4073 3268
rect 4097 3266 4153 3268
rect 4177 3266 4233 3268
rect 4257 3266 4313 3268
rect 4337 3266 4393 3268
rect 4017 3214 4019 3266
rect 4019 3214 4071 3266
rect 4071 3214 4073 3266
rect 4097 3214 4135 3266
rect 4135 3214 4147 3266
rect 4147 3214 4153 3266
rect 4177 3214 4199 3266
rect 4199 3214 4211 3266
rect 4211 3214 4233 3266
rect 4257 3214 4263 3266
rect 4263 3214 4275 3266
rect 4275 3214 4313 3266
rect 4337 3214 4339 3266
rect 4339 3214 4391 3266
rect 4391 3214 4393 3266
rect 4017 3212 4073 3214
rect 4097 3212 4153 3214
rect 4177 3212 4233 3214
rect 4257 3212 4313 3214
rect 4337 3212 4393 3214
rect 5948 3266 6004 3268
rect 6028 3266 6084 3268
rect 6108 3266 6164 3268
rect 6188 3266 6244 3268
rect 6268 3266 6324 3268
rect 5948 3214 5950 3266
rect 5950 3214 6002 3266
rect 6002 3214 6004 3266
rect 6028 3214 6066 3266
rect 6066 3214 6078 3266
rect 6078 3214 6084 3266
rect 6108 3214 6130 3266
rect 6130 3214 6142 3266
rect 6142 3214 6164 3266
rect 6188 3214 6194 3266
rect 6194 3214 6206 3266
rect 6206 3214 6244 3266
rect 6268 3214 6270 3266
rect 6270 3214 6322 3266
rect 6322 3214 6324 3266
rect 5948 3212 6004 3214
rect 6028 3212 6084 3214
rect 6108 3212 6164 3214
rect 6188 3212 6244 3214
rect 6268 3212 6324 3214
rect 7878 3266 7934 3268
rect 7958 3266 8014 3268
rect 8038 3266 8094 3268
rect 8118 3266 8174 3268
rect 8198 3266 8254 3268
rect 7878 3214 7880 3266
rect 7880 3214 7932 3266
rect 7932 3214 7934 3266
rect 7958 3214 7996 3266
rect 7996 3214 8008 3266
rect 8008 3214 8014 3266
rect 8038 3214 8060 3266
rect 8060 3214 8072 3266
rect 8072 3214 8094 3266
rect 8118 3214 8124 3266
rect 8124 3214 8136 3266
rect 8136 3214 8174 3266
rect 8198 3214 8200 3266
rect 8200 3214 8252 3266
rect 8252 3214 8254 3266
rect 7878 3212 7934 3214
rect 7958 3212 8014 3214
rect 8038 3212 8094 3214
rect 8118 3212 8174 3214
rect 8198 3212 8254 3214
<< metal3 >>
rect 0 9736 12184 9744
rect 0 9672 8 9736
rect 72 9672 88 9736
rect 152 9672 168 9736
rect 232 9672 248 9736
rect 312 9672 328 9736
rect 392 9672 408 9736
rect 472 9672 488 9736
rect 552 9672 568 9736
rect 632 9672 648 9736
rect 712 9672 728 9736
rect 792 9672 4978 9736
rect 5042 9672 5058 9736
rect 5122 9672 5138 9736
rect 5202 9672 5218 9736
rect 5282 9672 5298 9736
rect 5362 9672 6909 9736
rect 6973 9672 6989 9736
rect 7053 9672 7069 9736
rect 7133 9672 7149 9736
rect 7213 9672 7229 9736
rect 7293 9672 11392 9736
rect 11456 9672 11472 9736
rect 11536 9672 11552 9736
rect 11616 9672 11632 9736
rect 11696 9672 11712 9736
rect 11776 9672 11792 9736
rect 11856 9672 11872 9736
rect 11936 9672 11952 9736
rect 12016 9672 12032 9736
rect 12096 9672 12112 9736
rect 12176 9672 12184 9736
rect 0 9656 12184 9672
rect 0 9592 8 9656
rect 72 9592 88 9656
rect 152 9592 168 9656
rect 232 9592 248 9656
rect 312 9592 328 9656
rect 392 9592 408 9656
rect 472 9592 488 9656
rect 552 9592 568 9656
rect 632 9592 648 9656
rect 712 9592 728 9656
rect 792 9592 4978 9656
rect 5042 9592 5058 9656
rect 5122 9592 5138 9656
rect 5202 9592 5218 9656
rect 5282 9592 5298 9656
rect 5362 9592 6909 9656
rect 6973 9592 6989 9656
rect 7053 9592 7069 9656
rect 7133 9592 7149 9656
rect 7213 9592 7229 9656
rect 7293 9592 11392 9656
rect 11456 9592 11472 9656
rect 11536 9592 11552 9656
rect 11616 9592 11632 9656
rect 11696 9592 11712 9656
rect 11776 9592 11792 9656
rect 11856 9592 11872 9656
rect 11936 9592 11952 9656
rect 12016 9592 12032 9656
rect 12096 9592 12112 9656
rect 12176 9592 12184 9656
rect 0 9576 12184 9592
rect 0 9512 8 9576
rect 72 9512 88 9576
rect 152 9512 168 9576
rect 232 9512 248 9576
rect 312 9512 328 9576
rect 392 9512 408 9576
rect 472 9512 488 9576
rect 552 9512 568 9576
rect 632 9512 648 9576
rect 712 9512 728 9576
rect 792 9512 4978 9576
rect 5042 9512 5058 9576
rect 5122 9512 5138 9576
rect 5202 9512 5218 9576
rect 5282 9512 5298 9576
rect 5362 9512 6909 9576
rect 6973 9512 6989 9576
rect 7053 9512 7069 9576
rect 7133 9512 7149 9576
rect 7213 9512 7229 9576
rect 7293 9512 11392 9576
rect 11456 9512 11472 9576
rect 11536 9512 11552 9576
rect 11616 9512 11632 9576
rect 11696 9512 11712 9576
rect 11776 9512 11792 9576
rect 11856 9512 11872 9576
rect 11936 9512 11952 9576
rect 12016 9512 12032 9576
rect 12096 9512 12112 9576
rect 12176 9512 12184 9576
rect 0 9496 12184 9512
rect 0 9432 8 9496
rect 72 9432 88 9496
rect 152 9432 168 9496
rect 232 9432 248 9496
rect 312 9432 328 9496
rect 392 9432 408 9496
rect 472 9432 488 9496
rect 552 9432 568 9496
rect 632 9432 648 9496
rect 712 9432 728 9496
rect 792 9432 4978 9496
rect 5042 9432 5058 9496
rect 5122 9432 5138 9496
rect 5202 9432 5218 9496
rect 5282 9432 5298 9496
rect 5362 9432 6909 9496
rect 6973 9432 6989 9496
rect 7053 9432 7069 9496
rect 7133 9432 7149 9496
rect 7213 9432 7229 9496
rect 7293 9432 11392 9496
rect 11456 9432 11472 9496
rect 11536 9432 11552 9496
rect 11616 9432 11632 9496
rect 11696 9432 11712 9496
rect 11776 9432 11792 9496
rect 11856 9432 11872 9496
rect 11936 9432 11952 9496
rect 12016 9432 12032 9496
rect 12096 9432 12112 9496
rect 12176 9432 12184 9496
rect 0 9416 12184 9432
rect 0 9352 8 9416
rect 72 9352 88 9416
rect 152 9352 168 9416
rect 232 9352 248 9416
rect 312 9352 328 9416
rect 392 9352 408 9416
rect 472 9352 488 9416
rect 552 9352 568 9416
rect 632 9352 648 9416
rect 712 9352 728 9416
rect 792 9352 4978 9416
rect 5042 9352 5058 9416
rect 5122 9352 5138 9416
rect 5202 9352 5218 9416
rect 5282 9352 5298 9416
rect 5362 9352 6909 9416
rect 6973 9352 6989 9416
rect 7053 9352 7069 9416
rect 7133 9352 7149 9416
rect 7213 9352 7229 9416
rect 7293 9352 11392 9416
rect 11456 9352 11472 9416
rect 11536 9352 11552 9416
rect 11616 9352 11632 9416
rect 11696 9352 11712 9416
rect 11776 9352 11792 9416
rect 11856 9352 11872 9416
rect 11936 9352 11952 9416
rect 12016 9352 12032 9416
rect 12096 9352 12112 9416
rect 12176 9352 12184 9416
rect 0 9336 12184 9352
rect 0 9272 8 9336
rect 72 9272 88 9336
rect 152 9272 168 9336
rect 232 9272 248 9336
rect 312 9272 328 9336
rect 392 9272 408 9336
rect 472 9272 488 9336
rect 552 9272 568 9336
rect 632 9272 648 9336
rect 712 9272 728 9336
rect 792 9272 4978 9336
rect 5042 9272 5058 9336
rect 5122 9272 5138 9336
rect 5202 9272 5218 9336
rect 5282 9272 5298 9336
rect 5362 9272 6909 9336
rect 6973 9272 6989 9336
rect 7053 9272 7069 9336
rect 7133 9272 7149 9336
rect 7213 9272 7229 9336
rect 7293 9272 11392 9336
rect 11456 9272 11472 9336
rect 11536 9272 11552 9336
rect 11616 9272 11632 9336
rect 11696 9272 11712 9336
rect 11776 9272 11792 9336
rect 11856 9272 11872 9336
rect 11936 9272 11952 9336
rect 12016 9272 12032 9336
rect 12096 9272 12112 9336
rect 12176 9272 12184 9336
rect 0 9256 12184 9272
rect 0 9192 8 9256
rect 72 9192 88 9256
rect 152 9192 168 9256
rect 232 9192 248 9256
rect 312 9192 328 9256
rect 392 9192 408 9256
rect 472 9192 488 9256
rect 552 9192 568 9256
rect 632 9192 648 9256
rect 712 9192 728 9256
rect 792 9192 4978 9256
rect 5042 9192 5058 9256
rect 5122 9192 5138 9256
rect 5202 9192 5218 9256
rect 5282 9192 5298 9256
rect 5362 9192 6909 9256
rect 6973 9192 6989 9256
rect 7053 9192 7069 9256
rect 7133 9192 7149 9256
rect 7213 9192 7229 9256
rect 7293 9192 11392 9256
rect 11456 9192 11472 9256
rect 11536 9192 11552 9256
rect 11616 9192 11632 9256
rect 11696 9192 11712 9256
rect 11776 9192 11792 9256
rect 11856 9192 11872 9256
rect 11936 9192 11952 9256
rect 12016 9192 12032 9256
rect 12096 9192 12112 9256
rect 12176 9192 12184 9256
rect 0 9176 12184 9192
rect 0 9112 8 9176
rect 72 9112 88 9176
rect 152 9112 168 9176
rect 232 9112 248 9176
rect 312 9112 328 9176
rect 392 9112 408 9176
rect 472 9112 488 9176
rect 552 9112 568 9176
rect 632 9112 648 9176
rect 712 9112 728 9176
rect 792 9112 4978 9176
rect 5042 9112 5058 9176
rect 5122 9112 5138 9176
rect 5202 9112 5218 9176
rect 5282 9112 5298 9176
rect 5362 9112 6909 9176
rect 6973 9112 6989 9176
rect 7053 9112 7069 9176
rect 7133 9112 7149 9176
rect 7213 9112 7229 9176
rect 7293 9112 11392 9176
rect 11456 9112 11472 9176
rect 11536 9112 11552 9176
rect 11616 9112 11632 9176
rect 11696 9112 11712 9176
rect 11776 9112 11792 9176
rect 11856 9112 11872 9176
rect 11936 9112 11952 9176
rect 12016 9112 12032 9176
rect 12096 9112 12112 9176
rect 12176 9112 12184 9176
rect 0 9096 12184 9112
rect 0 9032 8 9096
rect 72 9032 88 9096
rect 152 9032 168 9096
rect 232 9032 248 9096
rect 312 9032 328 9096
rect 392 9032 408 9096
rect 472 9032 488 9096
rect 552 9032 568 9096
rect 632 9032 648 9096
rect 712 9032 728 9096
rect 792 9032 4978 9096
rect 5042 9032 5058 9096
rect 5122 9032 5138 9096
rect 5202 9032 5218 9096
rect 5282 9032 5298 9096
rect 5362 9032 6909 9096
rect 6973 9032 6989 9096
rect 7053 9032 7069 9096
rect 7133 9032 7149 9096
rect 7213 9032 7229 9096
rect 7293 9032 11392 9096
rect 11456 9032 11472 9096
rect 11536 9032 11552 9096
rect 11616 9032 11632 9096
rect 11696 9032 11712 9096
rect 11776 9032 11792 9096
rect 11856 9032 11872 9096
rect 11936 9032 11952 9096
rect 12016 9032 12032 9096
rect 12096 9032 12112 9096
rect 12176 9032 12184 9096
rect 0 9016 12184 9032
rect 0 8952 8 9016
rect 72 8952 88 9016
rect 152 8952 168 9016
rect 232 8952 248 9016
rect 312 8952 328 9016
rect 392 8952 408 9016
rect 472 8952 488 9016
rect 552 8952 568 9016
rect 632 8952 648 9016
rect 712 8952 728 9016
rect 792 8952 4978 9016
rect 5042 8952 5058 9016
rect 5122 8952 5138 9016
rect 5202 8952 5218 9016
rect 5282 8952 5298 9016
rect 5362 8952 6909 9016
rect 6973 8952 6989 9016
rect 7053 8952 7069 9016
rect 7133 8952 7149 9016
rect 7213 8952 7229 9016
rect 7293 8952 11392 9016
rect 11456 8952 11472 9016
rect 11536 8952 11552 9016
rect 11616 8952 11632 9016
rect 11696 8952 11712 9016
rect 11776 8952 11792 9016
rect 11856 8952 11872 9016
rect 11936 8952 11952 9016
rect 12016 8952 12032 9016
rect 12096 8952 12112 9016
rect 12176 8952 12184 9016
rect 0 8944 12184 8952
rect 1140 8596 11044 8604
rect 1140 8532 1148 8596
rect 1212 8532 1228 8596
rect 1292 8532 1308 8596
rect 1372 8532 1388 8596
rect 1452 8532 1468 8596
rect 1532 8532 1548 8596
rect 1612 8532 1628 8596
rect 1692 8532 1708 8596
rect 1772 8532 1788 8596
rect 1852 8532 1868 8596
rect 1932 8532 4013 8596
rect 4077 8532 4093 8596
rect 4157 8532 4173 8596
rect 4237 8532 4253 8596
rect 4317 8532 4333 8596
rect 4397 8532 5944 8596
rect 6008 8532 6024 8596
rect 6088 8532 6104 8596
rect 6168 8532 6184 8596
rect 6248 8532 6264 8596
rect 6328 8532 7874 8596
rect 7938 8532 7954 8596
rect 8018 8532 8034 8596
rect 8098 8532 8114 8596
rect 8178 8532 8194 8596
rect 8258 8532 10252 8596
rect 10316 8532 10332 8596
rect 10396 8532 10412 8596
rect 10476 8532 10492 8596
rect 10556 8532 10572 8596
rect 10636 8532 10652 8596
rect 10716 8532 10732 8596
rect 10796 8532 10812 8596
rect 10876 8532 10892 8596
rect 10956 8532 10972 8596
rect 11036 8532 11044 8596
rect 1140 8516 11044 8532
rect 1140 8452 1148 8516
rect 1212 8452 1228 8516
rect 1292 8452 1308 8516
rect 1372 8452 1388 8516
rect 1452 8452 1468 8516
rect 1532 8452 1548 8516
rect 1612 8452 1628 8516
rect 1692 8452 1708 8516
rect 1772 8452 1788 8516
rect 1852 8452 1868 8516
rect 1932 8452 4013 8516
rect 4077 8452 4093 8516
rect 4157 8452 4173 8516
rect 4237 8452 4253 8516
rect 4317 8452 4333 8516
rect 4397 8452 5944 8516
rect 6008 8452 6024 8516
rect 6088 8452 6104 8516
rect 6168 8452 6184 8516
rect 6248 8452 6264 8516
rect 6328 8452 7874 8516
rect 7938 8452 7954 8516
rect 8018 8452 8034 8516
rect 8098 8452 8114 8516
rect 8178 8452 8194 8516
rect 8258 8452 10252 8516
rect 10316 8452 10332 8516
rect 10396 8452 10412 8516
rect 10476 8452 10492 8516
rect 10556 8452 10572 8516
rect 10636 8452 10652 8516
rect 10716 8452 10732 8516
rect 10796 8452 10812 8516
rect 10876 8452 10892 8516
rect 10956 8452 10972 8516
rect 11036 8452 11044 8516
rect 1140 8436 11044 8452
rect 1140 8372 1148 8436
rect 1212 8372 1228 8436
rect 1292 8372 1308 8436
rect 1372 8372 1388 8436
rect 1452 8372 1468 8436
rect 1532 8372 1548 8436
rect 1612 8372 1628 8436
rect 1692 8372 1708 8436
rect 1772 8372 1788 8436
rect 1852 8372 1868 8436
rect 1932 8372 4013 8436
rect 4077 8372 4093 8436
rect 4157 8372 4173 8436
rect 4237 8372 4253 8436
rect 4317 8372 4333 8436
rect 4397 8372 5944 8436
rect 6008 8372 6024 8436
rect 6088 8372 6104 8436
rect 6168 8372 6184 8436
rect 6248 8372 6264 8436
rect 6328 8372 7874 8436
rect 7938 8372 7954 8436
rect 8018 8372 8034 8436
rect 8098 8372 8114 8436
rect 8178 8372 8194 8436
rect 8258 8372 10252 8436
rect 10316 8372 10332 8436
rect 10396 8372 10412 8436
rect 10476 8372 10492 8436
rect 10556 8372 10572 8436
rect 10636 8372 10652 8436
rect 10716 8372 10732 8436
rect 10796 8372 10812 8436
rect 10876 8372 10892 8436
rect 10956 8372 10972 8436
rect 11036 8372 11044 8436
rect 1140 8356 11044 8372
rect 1140 8292 1148 8356
rect 1212 8292 1228 8356
rect 1292 8292 1308 8356
rect 1372 8292 1388 8356
rect 1452 8292 1468 8356
rect 1532 8292 1548 8356
rect 1612 8292 1628 8356
rect 1692 8292 1708 8356
rect 1772 8292 1788 8356
rect 1852 8292 1868 8356
rect 1932 8292 4013 8356
rect 4077 8292 4093 8356
rect 4157 8292 4173 8356
rect 4237 8292 4253 8356
rect 4317 8292 4333 8356
rect 4397 8292 5944 8356
rect 6008 8292 6024 8356
rect 6088 8292 6104 8356
rect 6168 8292 6184 8356
rect 6248 8292 6264 8356
rect 6328 8292 7874 8356
rect 7938 8292 7954 8356
rect 8018 8292 8034 8356
rect 8098 8292 8114 8356
rect 8178 8292 8194 8356
rect 8258 8292 10252 8356
rect 10316 8292 10332 8356
rect 10396 8292 10412 8356
rect 10476 8292 10492 8356
rect 10556 8292 10572 8356
rect 10636 8292 10652 8356
rect 10716 8292 10732 8356
rect 10796 8292 10812 8356
rect 10876 8292 10892 8356
rect 10956 8292 10972 8356
rect 11036 8292 11044 8356
rect 1140 8276 11044 8292
rect 1140 8212 1148 8276
rect 1212 8212 1228 8276
rect 1292 8212 1308 8276
rect 1372 8212 1388 8276
rect 1452 8212 1468 8276
rect 1532 8212 1548 8276
rect 1612 8212 1628 8276
rect 1692 8212 1708 8276
rect 1772 8212 1788 8276
rect 1852 8212 1868 8276
rect 1932 8212 4013 8276
rect 4077 8212 4093 8276
rect 4157 8212 4173 8276
rect 4237 8212 4253 8276
rect 4317 8212 4333 8276
rect 4397 8212 5944 8276
rect 6008 8212 6024 8276
rect 6088 8212 6104 8276
rect 6168 8212 6184 8276
rect 6248 8212 6264 8276
rect 6328 8212 7874 8276
rect 7938 8212 7954 8276
rect 8018 8212 8034 8276
rect 8098 8212 8114 8276
rect 8178 8212 8194 8276
rect 8258 8212 10252 8276
rect 10316 8212 10332 8276
rect 10396 8212 10412 8276
rect 10476 8212 10492 8276
rect 10556 8212 10572 8276
rect 10636 8212 10652 8276
rect 10716 8212 10732 8276
rect 10796 8212 10812 8276
rect 10876 8212 10892 8276
rect 10956 8212 10972 8276
rect 11036 8212 11044 8276
rect 1140 8196 11044 8212
rect 1140 8132 1148 8196
rect 1212 8132 1228 8196
rect 1292 8132 1308 8196
rect 1372 8132 1388 8196
rect 1452 8132 1468 8196
rect 1532 8132 1548 8196
rect 1612 8132 1628 8196
rect 1692 8132 1708 8196
rect 1772 8132 1788 8196
rect 1852 8132 1868 8196
rect 1932 8132 4013 8196
rect 4077 8132 4093 8196
rect 4157 8132 4173 8196
rect 4237 8132 4253 8196
rect 4317 8132 4333 8196
rect 4397 8132 5944 8196
rect 6008 8132 6024 8196
rect 6088 8132 6104 8196
rect 6168 8132 6184 8196
rect 6248 8132 6264 8196
rect 6328 8132 7874 8196
rect 7938 8132 7954 8196
rect 8018 8132 8034 8196
rect 8098 8132 8114 8196
rect 8178 8132 8194 8196
rect 8258 8132 10252 8196
rect 10316 8132 10332 8196
rect 10396 8132 10412 8196
rect 10476 8132 10492 8196
rect 10556 8132 10572 8196
rect 10636 8132 10652 8196
rect 10716 8132 10732 8196
rect 10796 8132 10812 8196
rect 10876 8132 10892 8196
rect 10956 8132 10972 8196
rect 11036 8132 11044 8196
rect 1140 8116 11044 8132
rect 1140 8052 1148 8116
rect 1212 8052 1228 8116
rect 1292 8052 1308 8116
rect 1372 8052 1388 8116
rect 1452 8052 1468 8116
rect 1532 8052 1548 8116
rect 1612 8052 1628 8116
rect 1692 8052 1708 8116
rect 1772 8052 1788 8116
rect 1852 8052 1868 8116
rect 1932 8052 4013 8116
rect 4077 8052 4093 8116
rect 4157 8052 4173 8116
rect 4237 8052 4253 8116
rect 4317 8052 4333 8116
rect 4397 8052 5944 8116
rect 6008 8052 6024 8116
rect 6088 8052 6104 8116
rect 6168 8052 6184 8116
rect 6248 8052 6264 8116
rect 6328 8052 7874 8116
rect 7938 8052 7954 8116
rect 8018 8052 8034 8116
rect 8098 8052 8114 8116
rect 8178 8052 8194 8116
rect 8258 8052 10252 8116
rect 10316 8052 10332 8116
rect 10396 8052 10412 8116
rect 10476 8052 10492 8116
rect 10556 8052 10572 8116
rect 10636 8052 10652 8116
rect 10716 8052 10732 8116
rect 10796 8052 10812 8116
rect 10876 8052 10892 8116
rect 10956 8052 10972 8116
rect 11036 8052 11044 8116
rect 1140 8036 11044 8052
rect 1140 7972 1148 8036
rect 1212 7972 1228 8036
rect 1292 7972 1308 8036
rect 1372 7972 1388 8036
rect 1452 7972 1468 8036
rect 1532 7972 1548 8036
rect 1612 7972 1628 8036
rect 1692 7972 1708 8036
rect 1772 7972 1788 8036
rect 1852 7972 1868 8036
rect 1932 7972 4013 8036
rect 4077 7972 4093 8036
rect 4157 7972 4173 8036
rect 4237 7972 4253 8036
rect 4317 7972 4333 8036
rect 4397 7972 5944 8036
rect 6008 7972 6024 8036
rect 6088 7972 6104 8036
rect 6168 7972 6184 8036
rect 6248 7972 6264 8036
rect 6328 7972 7874 8036
rect 7938 7972 7954 8036
rect 8018 7972 8034 8036
rect 8098 7972 8114 8036
rect 8178 7972 8194 8036
rect 8258 7972 10252 8036
rect 10316 7972 10332 8036
rect 10396 7972 10412 8036
rect 10476 7972 10492 8036
rect 10556 7972 10572 8036
rect 10636 7972 10652 8036
rect 10716 7972 10732 8036
rect 10796 7972 10812 8036
rect 10876 7972 10892 8036
rect 10956 7972 10972 8036
rect 11036 7972 11044 8036
rect 1140 7956 11044 7972
rect 1140 7892 1148 7956
rect 1212 7892 1228 7956
rect 1292 7892 1308 7956
rect 1372 7892 1388 7956
rect 1452 7892 1468 7956
rect 1532 7892 1548 7956
rect 1612 7892 1628 7956
rect 1692 7892 1708 7956
rect 1772 7892 1788 7956
rect 1852 7892 1868 7956
rect 1932 7892 4013 7956
rect 4077 7892 4093 7956
rect 4157 7892 4173 7956
rect 4237 7892 4253 7956
rect 4317 7892 4333 7956
rect 4397 7892 5944 7956
rect 6008 7892 6024 7956
rect 6088 7892 6104 7956
rect 6168 7892 6184 7956
rect 6248 7892 6264 7956
rect 6328 7892 7874 7956
rect 7938 7892 7954 7956
rect 8018 7892 8034 7956
rect 8098 7892 8114 7956
rect 8178 7892 8194 7956
rect 8258 7892 10252 7956
rect 10316 7892 10332 7956
rect 10396 7892 10412 7956
rect 10476 7892 10492 7956
rect 10556 7892 10572 7956
rect 10636 7892 10652 7956
rect 10716 7892 10732 7956
rect 10796 7892 10812 7956
rect 10876 7892 10892 7956
rect 10956 7892 10972 7956
rect 11036 7892 11044 7956
rect 1140 7876 11044 7892
rect 1140 7812 1148 7876
rect 1212 7812 1228 7876
rect 1292 7812 1308 7876
rect 1372 7812 1388 7876
rect 1452 7812 1468 7876
rect 1532 7812 1548 7876
rect 1612 7812 1628 7876
rect 1692 7812 1708 7876
rect 1772 7812 1788 7876
rect 1852 7812 1868 7876
rect 1932 7812 4013 7876
rect 4077 7812 4093 7876
rect 4157 7812 4173 7876
rect 4237 7812 4253 7876
rect 4317 7812 4333 7876
rect 4397 7812 5944 7876
rect 6008 7812 6024 7876
rect 6088 7812 6104 7876
rect 6168 7812 6184 7876
rect 6248 7812 6264 7876
rect 6328 7812 7874 7876
rect 7938 7812 7954 7876
rect 8018 7812 8034 7876
rect 8098 7812 8114 7876
rect 8178 7812 8194 7876
rect 8258 7812 10252 7876
rect 10316 7812 10332 7876
rect 10396 7812 10412 7876
rect 10476 7812 10492 7876
rect 10556 7812 10572 7876
rect 10636 7812 10652 7876
rect 10716 7812 10732 7876
rect 10796 7812 10812 7876
rect 10876 7812 10892 7876
rect 10956 7812 10972 7876
rect 11036 7812 11044 7876
rect 1140 7804 11044 7812
rect 3995 6536 4415 6537
rect 3995 6472 4013 6536
rect 4077 6472 4093 6536
rect 4157 6472 4173 6536
rect 4237 6472 4253 6536
rect 4317 6472 4333 6536
rect 4397 6472 4415 6536
rect 3995 6471 4415 6472
rect 5926 6536 6346 6537
rect 5926 6472 5944 6536
rect 6008 6472 6024 6536
rect 6088 6472 6104 6536
rect 6168 6472 6184 6536
rect 6248 6472 6264 6536
rect 6328 6472 6346 6536
rect 5926 6471 6346 6472
rect 7856 6536 8276 6537
rect 7856 6472 7874 6536
rect 7938 6472 7954 6536
rect 8018 6472 8034 6536
rect 8098 6472 8114 6536
rect 8178 6472 8194 6536
rect 8258 6472 8276 6536
rect 7856 6471 8276 6472
rect 4960 5992 5380 5993
rect 4960 5928 4978 5992
rect 5042 5928 5058 5992
rect 5122 5928 5138 5992
rect 5202 5928 5218 5992
rect 5282 5928 5298 5992
rect 5362 5928 5380 5992
rect 4960 5927 5380 5928
rect 6891 5992 7311 5993
rect 6891 5928 6909 5992
rect 6973 5928 6989 5992
rect 7053 5928 7069 5992
rect 7133 5928 7149 5992
rect 7213 5928 7229 5992
rect 7293 5928 7311 5992
rect 6891 5927 7311 5928
rect 3995 5448 4415 5449
rect 3995 5384 4013 5448
rect 4077 5384 4093 5448
rect 4157 5384 4173 5448
rect 4237 5384 4253 5448
rect 4317 5384 4333 5448
rect 4397 5384 4415 5448
rect 3995 5383 4415 5384
rect 5926 5448 6346 5449
rect 5926 5384 5944 5448
rect 6008 5384 6024 5448
rect 6088 5384 6104 5448
rect 6168 5384 6184 5448
rect 6248 5384 6264 5448
rect 6328 5384 6346 5448
rect 5926 5383 6346 5384
rect 7856 5448 8276 5449
rect 7856 5384 7874 5448
rect 7938 5384 7954 5448
rect 8018 5384 8034 5448
rect 8098 5384 8114 5448
rect 8178 5384 8194 5448
rect 8258 5384 8276 5448
rect 7856 5383 8276 5384
rect 4960 4904 5380 4905
rect 4960 4840 4978 4904
rect 5042 4840 5058 4904
rect 5122 4840 5138 4904
rect 5202 4840 5218 4904
rect 5282 4840 5298 4904
rect 5362 4840 5380 4904
rect 4960 4839 5380 4840
rect 6891 4904 7311 4905
rect 6891 4840 6909 4904
rect 6973 4840 6989 4904
rect 7053 4840 7069 4904
rect 7133 4840 7149 4904
rect 7213 4840 7229 4904
rect 7293 4840 7311 4904
rect 6891 4839 7311 4840
rect 3995 4360 4415 4361
rect 3995 4296 4013 4360
rect 4077 4296 4093 4360
rect 4157 4296 4173 4360
rect 4237 4296 4253 4360
rect 4317 4296 4333 4360
rect 4397 4296 4415 4360
rect 3995 4295 4415 4296
rect 5926 4360 6346 4361
rect 5926 4296 5944 4360
rect 6008 4296 6024 4360
rect 6088 4296 6104 4360
rect 6168 4296 6184 4360
rect 6248 4296 6264 4360
rect 6328 4296 6346 4360
rect 5926 4295 6346 4296
rect 7856 4360 8276 4361
rect 7856 4296 7874 4360
rect 7938 4296 7954 4360
rect 8018 4296 8034 4360
rect 8098 4296 8114 4360
rect 8178 4296 8194 4360
rect 8258 4296 8276 4360
rect 7856 4295 8276 4296
rect 4960 3816 5380 3817
rect 4960 3752 4978 3816
rect 5042 3752 5058 3816
rect 5122 3752 5138 3816
rect 5202 3752 5218 3816
rect 5282 3752 5298 3816
rect 5362 3752 5380 3816
rect 4960 3751 5380 3752
rect 6891 3816 7311 3817
rect 6891 3752 6909 3816
rect 6973 3752 6989 3816
rect 7053 3752 7069 3816
rect 7133 3752 7149 3816
rect 7213 3752 7229 3816
rect 7293 3752 7311 3816
rect 6891 3751 7311 3752
rect 3995 3272 4415 3273
rect 3995 3208 4013 3272
rect 4077 3208 4093 3272
rect 4157 3208 4173 3272
rect 4237 3208 4253 3272
rect 4317 3208 4333 3272
rect 4397 3208 4415 3272
rect 3995 3207 4415 3208
rect 5926 3272 6346 3273
rect 5926 3208 5944 3272
rect 6008 3208 6024 3272
rect 6088 3208 6104 3272
rect 6168 3208 6184 3272
rect 6248 3208 6264 3272
rect 6328 3208 6346 3272
rect 5926 3207 6346 3208
rect 7856 3272 8276 3273
rect 7856 3208 7874 3272
rect 7938 3208 7954 3272
rect 8018 3208 8034 3272
rect 8098 3208 8114 3272
rect 8178 3208 8194 3272
rect 8258 3208 8276 3272
rect 7856 3207 8276 3208
rect 1140 1932 11044 1940
rect 1140 1868 1148 1932
rect 1212 1868 1228 1932
rect 1292 1868 1308 1932
rect 1372 1868 1388 1932
rect 1452 1868 1468 1932
rect 1532 1868 1548 1932
rect 1612 1868 1628 1932
rect 1692 1868 1708 1932
rect 1772 1868 1788 1932
rect 1852 1868 1868 1932
rect 1932 1868 4013 1932
rect 4077 1868 4093 1932
rect 4157 1868 4173 1932
rect 4237 1868 4253 1932
rect 4317 1868 4333 1932
rect 4397 1868 5944 1932
rect 6008 1868 6024 1932
rect 6088 1868 6104 1932
rect 6168 1868 6184 1932
rect 6248 1868 6264 1932
rect 6328 1868 7874 1932
rect 7938 1868 7954 1932
rect 8018 1868 8034 1932
rect 8098 1868 8114 1932
rect 8178 1868 8194 1932
rect 8258 1868 10252 1932
rect 10316 1868 10332 1932
rect 10396 1868 10412 1932
rect 10476 1868 10492 1932
rect 10556 1868 10572 1932
rect 10636 1868 10652 1932
rect 10716 1868 10732 1932
rect 10796 1868 10812 1932
rect 10876 1868 10892 1932
rect 10956 1868 10972 1932
rect 11036 1868 11044 1932
rect 1140 1852 11044 1868
rect 1140 1788 1148 1852
rect 1212 1788 1228 1852
rect 1292 1788 1308 1852
rect 1372 1788 1388 1852
rect 1452 1788 1468 1852
rect 1532 1788 1548 1852
rect 1612 1788 1628 1852
rect 1692 1788 1708 1852
rect 1772 1788 1788 1852
rect 1852 1788 1868 1852
rect 1932 1788 4013 1852
rect 4077 1788 4093 1852
rect 4157 1788 4173 1852
rect 4237 1788 4253 1852
rect 4317 1788 4333 1852
rect 4397 1788 5944 1852
rect 6008 1788 6024 1852
rect 6088 1788 6104 1852
rect 6168 1788 6184 1852
rect 6248 1788 6264 1852
rect 6328 1788 7874 1852
rect 7938 1788 7954 1852
rect 8018 1788 8034 1852
rect 8098 1788 8114 1852
rect 8178 1788 8194 1852
rect 8258 1788 10252 1852
rect 10316 1788 10332 1852
rect 10396 1788 10412 1852
rect 10476 1788 10492 1852
rect 10556 1788 10572 1852
rect 10636 1788 10652 1852
rect 10716 1788 10732 1852
rect 10796 1788 10812 1852
rect 10876 1788 10892 1852
rect 10956 1788 10972 1852
rect 11036 1788 11044 1852
rect 1140 1772 11044 1788
rect 1140 1708 1148 1772
rect 1212 1708 1228 1772
rect 1292 1708 1308 1772
rect 1372 1708 1388 1772
rect 1452 1708 1468 1772
rect 1532 1708 1548 1772
rect 1612 1708 1628 1772
rect 1692 1708 1708 1772
rect 1772 1708 1788 1772
rect 1852 1708 1868 1772
rect 1932 1708 4013 1772
rect 4077 1708 4093 1772
rect 4157 1708 4173 1772
rect 4237 1708 4253 1772
rect 4317 1708 4333 1772
rect 4397 1708 5944 1772
rect 6008 1708 6024 1772
rect 6088 1708 6104 1772
rect 6168 1708 6184 1772
rect 6248 1708 6264 1772
rect 6328 1708 7874 1772
rect 7938 1708 7954 1772
rect 8018 1708 8034 1772
rect 8098 1708 8114 1772
rect 8178 1708 8194 1772
rect 8258 1708 10252 1772
rect 10316 1708 10332 1772
rect 10396 1708 10412 1772
rect 10476 1708 10492 1772
rect 10556 1708 10572 1772
rect 10636 1708 10652 1772
rect 10716 1708 10732 1772
rect 10796 1708 10812 1772
rect 10876 1708 10892 1772
rect 10956 1708 10972 1772
rect 11036 1708 11044 1772
rect 1140 1692 11044 1708
rect 1140 1628 1148 1692
rect 1212 1628 1228 1692
rect 1292 1628 1308 1692
rect 1372 1628 1388 1692
rect 1452 1628 1468 1692
rect 1532 1628 1548 1692
rect 1612 1628 1628 1692
rect 1692 1628 1708 1692
rect 1772 1628 1788 1692
rect 1852 1628 1868 1692
rect 1932 1628 4013 1692
rect 4077 1628 4093 1692
rect 4157 1628 4173 1692
rect 4237 1628 4253 1692
rect 4317 1628 4333 1692
rect 4397 1628 5944 1692
rect 6008 1628 6024 1692
rect 6088 1628 6104 1692
rect 6168 1628 6184 1692
rect 6248 1628 6264 1692
rect 6328 1628 7874 1692
rect 7938 1628 7954 1692
rect 8018 1628 8034 1692
rect 8098 1628 8114 1692
rect 8178 1628 8194 1692
rect 8258 1628 10252 1692
rect 10316 1628 10332 1692
rect 10396 1628 10412 1692
rect 10476 1628 10492 1692
rect 10556 1628 10572 1692
rect 10636 1628 10652 1692
rect 10716 1628 10732 1692
rect 10796 1628 10812 1692
rect 10876 1628 10892 1692
rect 10956 1628 10972 1692
rect 11036 1628 11044 1692
rect 1140 1612 11044 1628
rect 1140 1548 1148 1612
rect 1212 1548 1228 1612
rect 1292 1548 1308 1612
rect 1372 1548 1388 1612
rect 1452 1548 1468 1612
rect 1532 1548 1548 1612
rect 1612 1548 1628 1612
rect 1692 1548 1708 1612
rect 1772 1548 1788 1612
rect 1852 1548 1868 1612
rect 1932 1548 4013 1612
rect 4077 1548 4093 1612
rect 4157 1548 4173 1612
rect 4237 1548 4253 1612
rect 4317 1548 4333 1612
rect 4397 1548 5944 1612
rect 6008 1548 6024 1612
rect 6088 1548 6104 1612
rect 6168 1548 6184 1612
rect 6248 1548 6264 1612
rect 6328 1548 7874 1612
rect 7938 1548 7954 1612
rect 8018 1548 8034 1612
rect 8098 1548 8114 1612
rect 8178 1548 8194 1612
rect 8258 1548 10252 1612
rect 10316 1548 10332 1612
rect 10396 1548 10412 1612
rect 10476 1548 10492 1612
rect 10556 1548 10572 1612
rect 10636 1548 10652 1612
rect 10716 1548 10732 1612
rect 10796 1548 10812 1612
rect 10876 1548 10892 1612
rect 10956 1548 10972 1612
rect 11036 1548 11044 1612
rect 1140 1532 11044 1548
rect 1140 1468 1148 1532
rect 1212 1468 1228 1532
rect 1292 1468 1308 1532
rect 1372 1468 1388 1532
rect 1452 1468 1468 1532
rect 1532 1468 1548 1532
rect 1612 1468 1628 1532
rect 1692 1468 1708 1532
rect 1772 1468 1788 1532
rect 1852 1468 1868 1532
rect 1932 1468 4013 1532
rect 4077 1468 4093 1532
rect 4157 1468 4173 1532
rect 4237 1468 4253 1532
rect 4317 1468 4333 1532
rect 4397 1468 5944 1532
rect 6008 1468 6024 1532
rect 6088 1468 6104 1532
rect 6168 1468 6184 1532
rect 6248 1468 6264 1532
rect 6328 1468 7874 1532
rect 7938 1468 7954 1532
rect 8018 1468 8034 1532
rect 8098 1468 8114 1532
rect 8178 1468 8194 1532
rect 8258 1468 10252 1532
rect 10316 1468 10332 1532
rect 10396 1468 10412 1532
rect 10476 1468 10492 1532
rect 10556 1468 10572 1532
rect 10636 1468 10652 1532
rect 10716 1468 10732 1532
rect 10796 1468 10812 1532
rect 10876 1468 10892 1532
rect 10956 1468 10972 1532
rect 11036 1468 11044 1532
rect 1140 1452 11044 1468
rect 1140 1388 1148 1452
rect 1212 1388 1228 1452
rect 1292 1388 1308 1452
rect 1372 1388 1388 1452
rect 1452 1388 1468 1452
rect 1532 1388 1548 1452
rect 1612 1388 1628 1452
rect 1692 1388 1708 1452
rect 1772 1388 1788 1452
rect 1852 1388 1868 1452
rect 1932 1388 4013 1452
rect 4077 1388 4093 1452
rect 4157 1388 4173 1452
rect 4237 1388 4253 1452
rect 4317 1388 4333 1452
rect 4397 1388 5944 1452
rect 6008 1388 6024 1452
rect 6088 1388 6104 1452
rect 6168 1388 6184 1452
rect 6248 1388 6264 1452
rect 6328 1388 7874 1452
rect 7938 1388 7954 1452
rect 8018 1388 8034 1452
rect 8098 1388 8114 1452
rect 8178 1388 8194 1452
rect 8258 1388 10252 1452
rect 10316 1388 10332 1452
rect 10396 1388 10412 1452
rect 10476 1388 10492 1452
rect 10556 1388 10572 1452
rect 10636 1388 10652 1452
rect 10716 1388 10732 1452
rect 10796 1388 10812 1452
rect 10876 1388 10892 1452
rect 10956 1388 10972 1452
rect 11036 1388 11044 1452
rect 1140 1372 11044 1388
rect 1140 1308 1148 1372
rect 1212 1308 1228 1372
rect 1292 1308 1308 1372
rect 1372 1308 1388 1372
rect 1452 1308 1468 1372
rect 1532 1308 1548 1372
rect 1612 1308 1628 1372
rect 1692 1308 1708 1372
rect 1772 1308 1788 1372
rect 1852 1308 1868 1372
rect 1932 1308 4013 1372
rect 4077 1308 4093 1372
rect 4157 1308 4173 1372
rect 4237 1308 4253 1372
rect 4317 1308 4333 1372
rect 4397 1308 5944 1372
rect 6008 1308 6024 1372
rect 6088 1308 6104 1372
rect 6168 1308 6184 1372
rect 6248 1308 6264 1372
rect 6328 1308 7874 1372
rect 7938 1308 7954 1372
rect 8018 1308 8034 1372
rect 8098 1308 8114 1372
rect 8178 1308 8194 1372
rect 8258 1308 10252 1372
rect 10316 1308 10332 1372
rect 10396 1308 10412 1372
rect 10476 1308 10492 1372
rect 10556 1308 10572 1372
rect 10636 1308 10652 1372
rect 10716 1308 10732 1372
rect 10796 1308 10812 1372
rect 10876 1308 10892 1372
rect 10956 1308 10972 1372
rect 11036 1308 11044 1372
rect 1140 1292 11044 1308
rect 1140 1228 1148 1292
rect 1212 1228 1228 1292
rect 1292 1228 1308 1292
rect 1372 1228 1388 1292
rect 1452 1228 1468 1292
rect 1532 1228 1548 1292
rect 1612 1228 1628 1292
rect 1692 1228 1708 1292
rect 1772 1228 1788 1292
rect 1852 1228 1868 1292
rect 1932 1228 4013 1292
rect 4077 1228 4093 1292
rect 4157 1228 4173 1292
rect 4237 1228 4253 1292
rect 4317 1228 4333 1292
rect 4397 1228 5944 1292
rect 6008 1228 6024 1292
rect 6088 1228 6104 1292
rect 6168 1228 6184 1292
rect 6248 1228 6264 1292
rect 6328 1228 7874 1292
rect 7938 1228 7954 1292
rect 8018 1228 8034 1292
rect 8098 1228 8114 1292
rect 8178 1228 8194 1292
rect 8258 1228 10252 1292
rect 10316 1228 10332 1292
rect 10396 1228 10412 1292
rect 10476 1228 10492 1292
rect 10556 1228 10572 1292
rect 10636 1228 10652 1292
rect 10716 1228 10732 1292
rect 10796 1228 10812 1292
rect 10876 1228 10892 1292
rect 10956 1228 10972 1292
rect 11036 1228 11044 1292
rect 1140 1212 11044 1228
rect 1140 1148 1148 1212
rect 1212 1148 1228 1212
rect 1292 1148 1308 1212
rect 1372 1148 1388 1212
rect 1452 1148 1468 1212
rect 1532 1148 1548 1212
rect 1612 1148 1628 1212
rect 1692 1148 1708 1212
rect 1772 1148 1788 1212
rect 1852 1148 1868 1212
rect 1932 1148 4013 1212
rect 4077 1148 4093 1212
rect 4157 1148 4173 1212
rect 4237 1148 4253 1212
rect 4317 1148 4333 1212
rect 4397 1148 5944 1212
rect 6008 1148 6024 1212
rect 6088 1148 6104 1212
rect 6168 1148 6184 1212
rect 6248 1148 6264 1212
rect 6328 1148 7874 1212
rect 7938 1148 7954 1212
rect 8018 1148 8034 1212
rect 8098 1148 8114 1212
rect 8178 1148 8194 1212
rect 8258 1148 10252 1212
rect 10316 1148 10332 1212
rect 10396 1148 10412 1212
rect 10476 1148 10492 1212
rect 10556 1148 10572 1212
rect 10636 1148 10652 1212
rect 10716 1148 10732 1212
rect 10796 1148 10812 1212
rect 10876 1148 10892 1212
rect 10956 1148 10972 1212
rect 11036 1148 11044 1212
rect 1140 1140 11044 1148
rect 0 792 12184 800
rect 0 728 8 792
rect 72 728 88 792
rect 152 728 168 792
rect 232 728 248 792
rect 312 728 328 792
rect 392 728 408 792
rect 472 728 488 792
rect 552 728 568 792
rect 632 728 648 792
rect 712 728 728 792
rect 792 728 4978 792
rect 5042 728 5058 792
rect 5122 728 5138 792
rect 5202 728 5218 792
rect 5282 728 5298 792
rect 5362 728 6909 792
rect 6973 728 6989 792
rect 7053 728 7069 792
rect 7133 728 7149 792
rect 7213 728 7229 792
rect 7293 728 11392 792
rect 11456 728 11472 792
rect 11536 728 11552 792
rect 11616 728 11632 792
rect 11696 728 11712 792
rect 11776 728 11792 792
rect 11856 728 11872 792
rect 11936 728 11952 792
rect 12016 728 12032 792
rect 12096 728 12112 792
rect 12176 728 12184 792
rect 0 712 12184 728
rect 0 648 8 712
rect 72 648 88 712
rect 152 648 168 712
rect 232 648 248 712
rect 312 648 328 712
rect 392 648 408 712
rect 472 648 488 712
rect 552 648 568 712
rect 632 648 648 712
rect 712 648 728 712
rect 792 648 4978 712
rect 5042 648 5058 712
rect 5122 648 5138 712
rect 5202 648 5218 712
rect 5282 648 5298 712
rect 5362 648 6909 712
rect 6973 648 6989 712
rect 7053 648 7069 712
rect 7133 648 7149 712
rect 7213 648 7229 712
rect 7293 648 11392 712
rect 11456 648 11472 712
rect 11536 648 11552 712
rect 11616 648 11632 712
rect 11696 648 11712 712
rect 11776 648 11792 712
rect 11856 648 11872 712
rect 11936 648 11952 712
rect 12016 648 12032 712
rect 12096 648 12112 712
rect 12176 648 12184 712
rect 0 632 12184 648
rect 0 568 8 632
rect 72 568 88 632
rect 152 568 168 632
rect 232 568 248 632
rect 312 568 328 632
rect 392 568 408 632
rect 472 568 488 632
rect 552 568 568 632
rect 632 568 648 632
rect 712 568 728 632
rect 792 568 4978 632
rect 5042 568 5058 632
rect 5122 568 5138 632
rect 5202 568 5218 632
rect 5282 568 5298 632
rect 5362 568 6909 632
rect 6973 568 6989 632
rect 7053 568 7069 632
rect 7133 568 7149 632
rect 7213 568 7229 632
rect 7293 568 11392 632
rect 11456 568 11472 632
rect 11536 568 11552 632
rect 11616 568 11632 632
rect 11696 568 11712 632
rect 11776 568 11792 632
rect 11856 568 11872 632
rect 11936 568 11952 632
rect 12016 568 12032 632
rect 12096 568 12112 632
rect 12176 568 12184 632
rect 0 552 12184 568
rect 0 488 8 552
rect 72 488 88 552
rect 152 488 168 552
rect 232 488 248 552
rect 312 488 328 552
rect 392 488 408 552
rect 472 488 488 552
rect 552 488 568 552
rect 632 488 648 552
rect 712 488 728 552
rect 792 488 4978 552
rect 5042 488 5058 552
rect 5122 488 5138 552
rect 5202 488 5218 552
rect 5282 488 5298 552
rect 5362 488 6909 552
rect 6973 488 6989 552
rect 7053 488 7069 552
rect 7133 488 7149 552
rect 7213 488 7229 552
rect 7293 488 11392 552
rect 11456 488 11472 552
rect 11536 488 11552 552
rect 11616 488 11632 552
rect 11696 488 11712 552
rect 11776 488 11792 552
rect 11856 488 11872 552
rect 11936 488 11952 552
rect 12016 488 12032 552
rect 12096 488 12112 552
rect 12176 488 12184 552
rect 0 472 12184 488
rect 0 408 8 472
rect 72 408 88 472
rect 152 408 168 472
rect 232 408 248 472
rect 312 408 328 472
rect 392 408 408 472
rect 472 408 488 472
rect 552 408 568 472
rect 632 408 648 472
rect 712 408 728 472
rect 792 408 4978 472
rect 5042 408 5058 472
rect 5122 408 5138 472
rect 5202 408 5218 472
rect 5282 408 5298 472
rect 5362 408 6909 472
rect 6973 408 6989 472
rect 7053 408 7069 472
rect 7133 408 7149 472
rect 7213 408 7229 472
rect 7293 408 11392 472
rect 11456 408 11472 472
rect 11536 408 11552 472
rect 11616 408 11632 472
rect 11696 408 11712 472
rect 11776 408 11792 472
rect 11856 408 11872 472
rect 11936 408 11952 472
rect 12016 408 12032 472
rect 12096 408 12112 472
rect 12176 408 12184 472
rect 0 392 12184 408
rect 0 328 8 392
rect 72 328 88 392
rect 152 328 168 392
rect 232 328 248 392
rect 312 328 328 392
rect 392 328 408 392
rect 472 328 488 392
rect 552 328 568 392
rect 632 328 648 392
rect 712 328 728 392
rect 792 328 4978 392
rect 5042 328 5058 392
rect 5122 328 5138 392
rect 5202 328 5218 392
rect 5282 328 5298 392
rect 5362 328 6909 392
rect 6973 328 6989 392
rect 7053 328 7069 392
rect 7133 328 7149 392
rect 7213 328 7229 392
rect 7293 328 11392 392
rect 11456 328 11472 392
rect 11536 328 11552 392
rect 11616 328 11632 392
rect 11696 328 11712 392
rect 11776 328 11792 392
rect 11856 328 11872 392
rect 11936 328 11952 392
rect 12016 328 12032 392
rect 12096 328 12112 392
rect 12176 328 12184 392
rect 0 312 12184 328
rect 0 248 8 312
rect 72 248 88 312
rect 152 248 168 312
rect 232 248 248 312
rect 312 248 328 312
rect 392 248 408 312
rect 472 248 488 312
rect 552 248 568 312
rect 632 248 648 312
rect 712 248 728 312
rect 792 248 4978 312
rect 5042 248 5058 312
rect 5122 248 5138 312
rect 5202 248 5218 312
rect 5282 248 5298 312
rect 5362 248 6909 312
rect 6973 248 6989 312
rect 7053 248 7069 312
rect 7133 248 7149 312
rect 7213 248 7229 312
rect 7293 248 11392 312
rect 11456 248 11472 312
rect 11536 248 11552 312
rect 11616 248 11632 312
rect 11696 248 11712 312
rect 11776 248 11792 312
rect 11856 248 11872 312
rect 11936 248 11952 312
rect 12016 248 12032 312
rect 12096 248 12112 312
rect 12176 248 12184 312
rect 0 232 12184 248
rect 0 168 8 232
rect 72 168 88 232
rect 152 168 168 232
rect 232 168 248 232
rect 312 168 328 232
rect 392 168 408 232
rect 472 168 488 232
rect 552 168 568 232
rect 632 168 648 232
rect 712 168 728 232
rect 792 168 4978 232
rect 5042 168 5058 232
rect 5122 168 5138 232
rect 5202 168 5218 232
rect 5282 168 5298 232
rect 5362 168 6909 232
rect 6973 168 6989 232
rect 7053 168 7069 232
rect 7133 168 7149 232
rect 7213 168 7229 232
rect 7293 168 11392 232
rect 11456 168 11472 232
rect 11536 168 11552 232
rect 11616 168 11632 232
rect 11696 168 11712 232
rect 11776 168 11792 232
rect 11856 168 11872 232
rect 11936 168 11952 232
rect 12016 168 12032 232
rect 12096 168 12112 232
rect 12176 168 12184 232
rect 0 152 12184 168
rect 0 88 8 152
rect 72 88 88 152
rect 152 88 168 152
rect 232 88 248 152
rect 312 88 328 152
rect 392 88 408 152
rect 472 88 488 152
rect 552 88 568 152
rect 632 88 648 152
rect 712 88 728 152
rect 792 88 4978 152
rect 5042 88 5058 152
rect 5122 88 5138 152
rect 5202 88 5218 152
rect 5282 88 5298 152
rect 5362 88 6909 152
rect 6973 88 6989 152
rect 7053 88 7069 152
rect 7133 88 7149 152
rect 7213 88 7229 152
rect 7293 88 11392 152
rect 11456 88 11472 152
rect 11536 88 11552 152
rect 11616 88 11632 152
rect 11696 88 11712 152
rect 11776 88 11792 152
rect 11856 88 11872 152
rect 11936 88 11952 152
rect 12016 88 12032 152
rect 12096 88 12112 152
rect 12176 88 12184 152
rect 0 72 12184 88
rect 0 8 8 72
rect 72 8 88 72
rect 152 8 168 72
rect 232 8 248 72
rect 312 8 328 72
rect 392 8 408 72
rect 472 8 488 72
rect 552 8 568 72
rect 632 8 648 72
rect 712 8 728 72
rect 792 8 4978 72
rect 5042 8 5058 72
rect 5122 8 5138 72
rect 5202 8 5218 72
rect 5282 8 5298 72
rect 5362 8 6909 72
rect 6973 8 6989 72
rect 7053 8 7069 72
rect 7133 8 7149 72
rect 7213 8 7229 72
rect 7293 8 11392 72
rect 11456 8 11472 72
rect 11536 8 11552 72
rect 11616 8 11632 72
rect 11696 8 11712 72
rect 11776 8 11792 72
rect 11856 8 11872 72
rect 11936 8 11952 72
rect 12016 8 12032 72
rect 12096 8 12112 72
rect 12176 8 12184 72
rect 0 0 12184 8
<< via3 >>
rect 8 9672 72 9736
rect 88 9672 152 9736
rect 168 9672 232 9736
rect 248 9672 312 9736
rect 328 9672 392 9736
rect 408 9672 472 9736
rect 488 9672 552 9736
rect 568 9672 632 9736
rect 648 9672 712 9736
rect 728 9672 792 9736
rect 4978 9672 5042 9736
rect 5058 9672 5122 9736
rect 5138 9672 5202 9736
rect 5218 9672 5282 9736
rect 5298 9672 5362 9736
rect 6909 9672 6973 9736
rect 6989 9672 7053 9736
rect 7069 9672 7133 9736
rect 7149 9672 7213 9736
rect 7229 9672 7293 9736
rect 11392 9672 11456 9736
rect 11472 9672 11536 9736
rect 11552 9672 11616 9736
rect 11632 9672 11696 9736
rect 11712 9672 11776 9736
rect 11792 9672 11856 9736
rect 11872 9672 11936 9736
rect 11952 9672 12016 9736
rect 12032 9672 12096 9736
rect 12112 9672 12176 9736
rect 8 9592 72 9656
rect 88 9592 152 9656
rect 168 9592 232 9656
rect 248 9592 312 9656
rect 328 9592 392 9656
rect 408 9592 472 9656
rect 488 9592 552 9656
rect 568 9592 632 9656
rect 648 9592 712 9656
rect 728 9592 792 9656
rect 4978 9592 5042 9656
rect 5058 9592 5122 9656
rect 5138 9592 5202 9656
rect 5218 9592 5282 9656
rect 5298 9592 5362 9656
rect 6909 9592 6973 9656
rect 6989 9592 7053 9656
rect 7069 9592 7133 9656
rect 7149 9592 7213 9656
rect 7229 9592 7293 9656
rect 11392 9592 11456 9656
rect 11472 9592 11536 9656
rect 11552 9592 11616 9656
rect 11632 9592 11696 9656
rect 11712 9592 11776 9656
rect 11792 9592 11856 9656
rect 11872 9592 11936 9656
rect 11952 9592 12016 9656
rect 12032 9592 12096 9656
rect 12112 9592 12176 9656
rect 8 9512 72 9576
rect 88 9512 152 9576
rect 168 9512 232 9576
rect 248 9512 312 9576
rect 328 9512 392 9576
rect 408 9512 472 9576
rect 488 9512 552 9576
rect 568 9512 632 9576
rect 648 9512 712 9576
rect 728 9512 792 9576
rect 4978 9512 5042 9576
rect 5058 9512 5122 9576
rect 5138 9512 5202 9576
rect 5218 9512 5282 9576
rect 5298 9512 5362 9576
rect 6909 9512 6973 9576
rect 6989 9512 7053 9576
rect 7069 9512 7133 9576
rect 7149 9512 7213 9576
rect 7229 9512 7293 9576
rect 11392 9512 11456 9576
rect 11472 9512 11536 9576
rect 11552 9512 11616 9576
rect 11632 9512 11696 9576
rect 11712 9512 11776 9576
rect 11792 9512 11856 9576
rect 11872 9512 11936 9576
rect 11952 9512 12016 9576
rect 12032 9512 12096 9576
rect 12112 9512 12176 9576
rect 8 9432 72 9496
rect 88 9432 152 9496
rect 168 9432 232 9496
rect 248 9432 312 9496
rect 328 9432 392 9496
rect 408 9432 472 9496
rect 488 9432 552 9496
rect 568 9432 632 9496
rect 648 9432 712 9496
rect 728 9432 792 9496
rect 4978 9432 5042 9496
rect 5058 9432 5122 9496
rect 5138 9432 5202 9496
rect 5218 9432 5282 9496
rect 5298 9432 5362 9496
rect 6909 9432 6973 9496
rect 6989 9432 7053 9496
rect 7069 9432 7133 9496
rect 7149 9432 7213 9496
rect 7229 9432 7293 9496
rect 11392 9432 11456 9496
rect 11472 9432 11536 9496
rect 11552 9432 11616 9496
rect 11632 9432 11696 9496
rect 11712 9432 11776 9496
rect 11792 9432 11856 9496
rect 11872 9432 11936 9496
rect 11952 9432 12016 9496
rect 12032 9432 12096 9496
rect 12112 9432 12176 9496
rect 8 9352 72 9416
rect 88 9352 152 9416
rect 168 9352 232 9416
rect 248 9352 312 9416
rect 328 9352 392 9416
rect 408 9352 472 9416
rect 488 9352 552 9416
rect 568 9352 632 9416
rect 648 9352 712 9416
rect 728 9352 792 9416
rect 4978 9352 5042 9416
rect 5058 9352 5122 9416
rect 5138 9352 5202 9416
rect 5218 9352 5282 9416
rect 5298 9352 5362 9416
rect 6909 9352 6973 9416
rect 6989 9352 7053 9416
rect 7069 9352 7133 9416
rect 7149 9352 7213 9416
rect 7229 9352 7293 9416
rect 11392 9352 11456 9416
rect 11472 9352 11536 9416
rect 11552 9352 11616 9416
rect 11632 9352 11696 9416
rect 11712 9352 11776 9416
rect 11792 9352 11856 9416
rect 11872 9352 11936 9416
rect 11952 9352 12016 9416
rect 12032 9352 12096 9416
rect 12112 9352 12176 9416
rect 8 9272 72 9336
rect 88 9272 152 9336
rect 168 9272 232 9336
rect 248 9272 312 9336
rect 328 9272 392 9336
rect 408 9272 472 9336
rect 488 9272 552 9336
rect 568 9272 632 9336
rect 648 9272 712 9336
rect 728 9272 792 9336
rect 4978 9272 5042 9336
rect 5058 9272 5122 9336
rect 5138 9272 5202 9336
rect 5218 9272 5282 9336
rect 5298 9272 5362 9336
rect 6909 9272 6973 9336
rect 6989 9272 7053 9336
rect 7069 9272 7133 9336
rect 7149 9272 7213 9336
rect 7229 9272 7293 9336
rect 11392 9272 11456 9336
rect 11472 9272 11536 9336
rect 11552 9272 11616 9336
rect 11632 9272 11696 9336
rect 11712 9272 11776 9336
rect 11792 9272 11856 9336
rect 11872 9272 11936 9336
rect 11952 9272 12016 9336
rect 12032 9272 12096 9336
rect 12112 9272 12176 9336
rect 8 9192 72 9256
rect 88 9192 152 9256
rect 168 9192 232 9256
rect 248 9192 312 9256
rect 328 9192 392 9256
rect 408 9192 472 9256
rect 488 9192 552 9256
rect 568 9192 632 9256
rect 648 9192 712 9256
rect 728 9192 792 9256
rect 4978 9192 5042 9256
rect 5058 9192 5122 9256
rect 5138 9192 5202 9256
rect 5218 9192 5282 9256
rect 5298 9192 5362 9256
rect 6909 9192 6973 9256
rect 6989 9192 7053 9256
rect 7069 9192 7133 9256
rect 7149 9192 7213 9256
rect 7229 9192 7293 9256
rect 11392 9192 11456 9256
rect 11472 9192 11536 9256
rect 11552 9192 11616 9256
rect 11632 9192 11696 9256
rect 11712 9192 11776 9256
rect 11792 9192 11856 9256
rect 11872 9192 11936 9256
rect 11952 9192 12016 9256
rect 12032 9192 12096 9256
rect 12112 9192 12176 9256
rect 8 9112 72 9176
rect 88 9112 152 9176
rect 168 9112 232 9176
rect 248 9112 312 9176
rect 328 9112 392 9176
rect 408 9112 472 9176
rect 488 9112 552 9176
rect 568 9112 632 9176
rect 648 9112 712 9176
rect 728 9112 792 9176
rect 4978 9112 5042 9176
rect 5058 9112 5122 9176
rect 5138 9112 5202 9176
rect 5218 9112 5282 9176
rect 5298 9112 5362 9176
rect 6909 9112 6973 9176
rect 6989 9112 7053 9176
rect 7069 9112 7133 9176
rect 7149 9112 7213 9176
rect 7229 9112 7293 9176
rect 11392 9112 11456 9176
rect 11472 9112 11536 9176
rect 11552 9112 11616 9176
rect 11632 9112 11696 9176
rect 11712 9112 11776 9176
rect 11792 9112 11856 9176
rect 11872 9112 11936 9176
rect 11952 9112 12016 9176
rect 12032 9112 12096 9176
rect 12112 9112 12176 9176
rect 8 9032 72 9096
rect 88 9032 152 9096
rect 168 9032 232 9096
rect 248 9032 312 9096
rect 328 9032 392 9096
rect 408 9032 472 9096
rect 488 9032 552 9096
rect 568 9032 632 9096
rect 648 9032 712 9096
rect 728 9032 792 9096
rect 4978 9032 5042 9096
rect 5058 9032 5122 9096
rect 5138 9032 5202 9096
rect 5218 9032 5282 9096
rect 5298 9032 5362 9096
rect 6909 9032 6973 9096
rect 6989 9032 7053 9096
rect 7069 9032 7133 9096
rect 7149 9032 7213 9096
rect 7229 9032 7293 9096
rect 11392 9032 11456 9096
rect 11472 9032 11536 9096
rect 11552 9032 11616 9096
rect 11632 9032 11696 9096
rect 11712 9032 11776 9096
rect 11792 9032 11856 9096
rect 11872 9032 11936 9096
rect 11952 9032 12016 9096
rect 12032 9032 12096 9096
rect 12112 9032 12176 9096
rect 8 8952 72 9016
rect 88 8952 152 9016
rect 168 8952 232 9016
rect 248 8952 312 9016
rect 328 8952 392 9016
rect 408 8952 472 9016
rect 488 8952 552 9016
rect 568 8952 632 9016
rect 648 8952 712 9016
rect 728 8952 792 9016
rect 4978 8952 5042 9016
rect 5058 8952 5122 9016
rect 5138 8952 5202 9016
rect 5218 8952 5282 9016
rect 5298 8952 5362 9016
rect 6909 8952 6973 9016
rect 6989 8952 7053 9016
rect 7069 8952 7133 9016
rect 7149 8952 7213 9016
rect 7229 8952 7293 9016
rect 11392 8952 11456 9016
rect 11472 8952 11536 9016
rect 11552 8952 11616 9016
rect 11632 8952 11696 9016
rect 11712 8952 11776 9016
rect 11792 8952 11856 9016
rect 11872 8952 11936 9016
rect 11952 8952 12016 9016
rect 12032 8952 12096 9016
rect 12112 8952 12176 9016
rect 1148 8532 1212 8596
rect 1228 8532 1292 8596
rect 1308 8532 1372 8596
rect 1388 8532 1452 8596
rect 1468 8532 1532 8596
rect 1548 8532 1612 8596
rect 1628 8532 1692 8596
rect 1708 8532 1772 8596
rect 1788 8532 1852 8596
rect 1868 8532 1932 8596
rect 4013 8532 4077 8596
rect 4093 8532 4157 8596
rect 4173 8532 4237 8596
rect 4253 8532 4317 8596
rect 4333 8532 4397 8596
rect 5944 8532 6008 8596
rect 6024 8532 6088 8596
rect 6104 8532 6168 8596
rect 6184 8532 6248 8596
rect 6264 8532 6328 8596
rect 7874 8532 7938 8596
rect 7954 8532 8018 8596
rect 8034 8532 8098 8596
rect 8114 8532 8178 8596
rect 8194 8532 8258 8596
rect 10252 8532 10316 8596
rect 10332 8532 10396 8596
rect 10412 8532 10476 8596
rect 10492 8532 10556 8596
rect 10572 8532 10636 8596
rect 10652 8532 10716 8596
rect 10732 8532 10796 8596
rect 10812 8532 10876 8596
rect 10892 8532 10956 8596
rect 10972 8532 11036 8596
rect 1148 8452 1212 8516
rect 1228 8452 1292 8516
rect 1308 8452 1372 8516
rect 1388 8452 1452 8516
rect 1468 8452 1532 8516
rect 1548 8452 1612 8516
rect 1628 8452 1692 8516
rect 1708 8452 1772 8516
rect 1788 8452 1852 8516
rect 1868 8452 1932 8516
rect 4013 8452 4077 8516
rect 4093 8452 4157 8516
rect 4173 8452 4237 8516
rect 4253 8452 4317 8516
rect 4333 8452 4397 8516
rect 5944 8452 6008 8516
rect 6024 8452 6088 8516
rect 6104 8452 6168 8516
rect 6184 8452 6248 8516
rect 6264 8452 6328 8516
rect 7874 8452 7938 8516
rect 7954 8452 8018 8516
rect 8034 8452 8098 8516
rect 8114 8452 8178 8516
rect 8194 8452 8258 8516
rect 10252 8452 10316 8516
rect 10332 8452 10396 8516
rect 10412 8452 10476 8516
rect 10492 8452 10556 8516
rect 10572 8452 10636 8516
rect 10652 8452 10716 8516
rect 10732 8452 10796 8516
rect 10812 8452 10876 8516
rect 10892 8452 10956 8516
rect 10972 8452 11036 8516
rect 1148 8372 1212 8436
rect 1228 8372 1292 8436
rect 1308 8372 1372 8436
rect 1388 8372 1452 8436
rect 1468 8372 1532 8436
rect 1548 8372 1612 8436
rect 1628 8372 1692 8436
rect 1708 8372 1772 8436
rect 1788 8372 1852 8436
rect 1868 8372 1932 8436
rect 4013 8372 4077 8436
rect 4093 8372 4157 8436
rect 4173 8372 4237 8436
rect 4253 8372 4317 8436
rect 4333 8372 4397 8436
rect 5944 8372 6008 8436
rect 6024 8372 6088 8436
rect 6104 8372 6168 8436
rect 6184 8372 6248 8436
rect 6264 8372 6328 8436
rect 7874 8372 7938 8436
rect 7954 8372 8018 8436
rect 8034 8372 8098 8436
rect 8114 8372 8178 8436
rect 8194 8372 8258 8436
rect 10252 8372 10316 8436
rect 10332 8372 10396 8436
rect 10412 8372 10476 8436
rect 10492 8372 10556 8436
rect 10572 8372 10636 8436
rect 10652 8372 10716 8436
rect 10732 8372 10796 8436
rect 10812 8372 10876 8436
rect 10892 8372 10956 8436
rect 10972 8372 11036 8436
rect 1148 8292 1212 8356
rect 1228 8292 1292 8356
rect 1308 8292 1372 8356
rect 1388 8292 1452 8356
rect 1468 8292 1532 8356
rect 1548 8292 1612 8356
rect 1628 8292 1692 8356
rect 1708 8292 1772 8356
rect 1788 8292 1852 8356
rect 1868 8292 1932 8356
rect 4013 8292 4077 8356
rect 4093 8292 4157 8356
rect 4173 8292 4237 8356
rect 4253 8292 4317 8356
rect 4333 8292 4397 8356
rect 5944 8292 6008 8356
rect 6024 8292 6088 8356
rect 6104 8292 6168 8356
rect 6184 8292 6248 8356
rect 6264 8292 6328 8356
rect 7874 8292 7938 8356
rect 7954 8292 8018 8356
rect 8034 8292 8098 8356
rect 8114 8292 8178 8356
rect 8194 8292 8258 8356
rect 10252 8292 10316 8356
rect 10332 8292 10396 8356
rect 10412 8292 10476 8356
rect 10492 8292 10556 8356
rect 10572 8292 10636 8356
rect 10652 8292 10716 8356
rect 10732 8292 10796 8356
rect 10812 8292 10876 8356
rect 10892 8292 10956 8356
rect 10972 8292 11036 8356
rect 1148 8212 1212 8276
rect 1228 8212 1292 8276
rect 1308 8212 1372 8276
rect 1388 8212 1452 8276
rect 1468 8212 1532 8276
rect 1548 8212 1612 8276
rect 1628 8212 1692 8276
rect 1708 8212 1772 8276
rect 1788 8212 1852 8276
rect 1868 8212 1932 8276
rect 4013 8212 4077 8276
rect 4093 8212 4157 8276
rect 4173 8212 4237 8276
rect 4253 8212 4317 8276
rect 4333 8212 4397 8276
rect 5944 8212 6008 8276
rect 6024 8212 6088 8276
rect 6104 8212 6168 8276
rect 6184 8212 6248 8276
rect 6264 8212 6328 8276
rect 7874 8212 7938 8276
rect 7954 8212 8018 8276
rect 8034 8212 8098 8276
rect 8114 8212 8178 8276
rect 8194 8212 8258 8276
rect 10252 8212 10316 8276
rect 10332 8212 10396 8276
rect 10412 8212 10476 8276
rect 10492 8212 10556 8276
rect 10572 8212 10636 8276
rect 10652 8212 10716 8276
rect 10732 8212 10796 8276
rect 10812 8212 10876 8276
rect 10892 8212 10956 8276
rect 10972 8212 11036 8276
rect 1148 8132 1212 8196
rect 1228 8132 1292 8196
rect 1308 8132 1372 8196
rect 1388 8132 1452 8196
rect 1468 8132 1532 8196
rect 1548 8132 1612 8196
rect 1628 8132 1692 8196
rect 1708 8132 1772 8196
rect 1788 8132 1852 8196
rect 1868 8132 1932 8196
rect 4013 8132 4077 8196
rect 4093 8132 4157 8196
rect 4173 8132 4237 8196
rect 4253 8132 4317 8196
rect 4333 8132 4397 8196
rect 5944 8132 6008 8196
rect 6024 8132 6088 8196
rect 6104 8132 6168 8196
rect 6184 8132 6248 8196
rect 6264 8132 6328 8196
rect 7874 8132 7938 8196
rect 7954 8132 8018 8196
rect 8034 8132 8098 8196
rect 8114 8132 8178 8196
rect 8194 8132 8258 8196
rect 10252 8132 10316 8196
rect 10332 8132 10396 8196
rect 10412 8132 10476 8196
rect 10492 8132 10556 8196
rect 10572 8132 10636 8196
rect 10652 8132 10716 8196
rect 10732 8132 10796 8196
rect 10812 8132 10876 8196
rect 10892 8132 10956 8196
rect 10972 8132 11036 8196
rect 1148 8052 1212 8116
rect 1228 8052 1292 8116
rect 1308 8052 1372 8116
rect 1388 8052 1452 8116
rect 1468 8052 1532 8116
rect 1548 8052 1612 8116
rect 1628 8052 1692 8116
rect 1708 8052 1772 8116
rect 1788 8052 1852 8116
rect 1868 8052 1932 8116
rect 4013 8052 4077 8116
rect 4093 8052 4157 8116
rect 4173 8052 4237 8116
rect 4253 8052 4317 8116
rect 4333 8052 4397 8116
rect 5944 8052 6008 8116
rect 6024 8052 6088 8116
rect 6104 8052 6168 8116
rect 6184 8052 6248 8116
rect 6264 8052 6328 8116
rect 7874 8052 7938 8116
rect 7954 8052 8018 8116
rect 8034 8052 8098 8116
rect 8114 8052 8178 8116
rect 8194 8052 8258 8116
rect 10252 8052 10316 8116
rect 10332 8052 10396 8116
rect 10412 8052 10476 8116
rect 10492 8052 10556 8116
rect 10572 8052 10636 8116
rect 10652 8052 10716 8116
rect 10732 8052 10796 8116
rect 10812 8052 10876 8116
rect 10892 8052 10956 8116
rect 10972 8052 11036 8116
rect 1148 7972 1212 8036
rect 1228 7972 1292 8036
rect 1308 7972 1372 8036
rect 1388 7972 1452 8036
rect 1468 7972 1532 8036
rect 1548 7972 1612 8036
rect 1628 7972 1692 8036
rect 1708 7972 1772 8036
rect 1788 7972 1852 8036
rect 1868 7972 1932 8036
rect 4013 7972 4077 8036
rect 4093 7972 4157 8036
rect 4173 7972 4237 8036
rect 4253 7972 4317 8036
rect 4333 7972 4397 8036
rect 5944 7972 6008 8036
rect 6024 7972 6088 8036
rect 6104 7972 6168 8036
rect 6184 7972 6248 8036
rect 6264 7972 6328 8036
rect 7874 7972 7938 8036
rect 7954 7972 8018 8036
rect 8034 7972 8098 8036
rect 8114 7972 8178 8036
rect 8194 7972 8258 8036
rect 10252 7972 10316 8036
rect 10332 7972 10396 8036
rect 10412 7972 10476 8036
rect 10492 7972 10556 8036
rect 10572 7972 10636 8036
rect 10652 7972 10716 8036
rect 10732 7972 10796 8036
rect 10812 7972 10876 8036
rect 10892 7972 10956 8036
rect 10972 7972 11036 8036
rect 1148 7892 1212 7956
rect 1228 7892 1292 7956
rect 1308 7892 1372 7956
rect 1388 7892 1452 7956
rect 1468 7892 1532 7956
rect 1548 7892 1612 7956
rect 1628 7892 1692 7956
rect 1708 7892 1772 7956
rect 1788 7892 1852 7956
rect 1868 7892 1932 7956
rect 4013 7892 4077 7956
rect 4093 7892 4157 7956
rect 4173 7892 4237 7956
rect 4253 7892 4317 7956
rect 4333 7892 4397 7956
rect 5944 7892 6008 7956
rect 6024 7892 6088 7956
rect 6104 7892 6168 7956
rect 6184 7892 6248 7956
rect 6264 7892 6328 7956
rect 7874 7892 7938 7956
rect 7954 7892 8018 7956
rect 8034 7892 8098 7956
rect 8114 7892 8178 7956
rect 8194 7892 8258 7956
rect 10252 7892 10316 7956
rect 10332 7892 10396 7956
rect 10412 7892 10476 7956
rect 10492 7892 10556 7956
rect 10572 7892 10636 7956
rect 10652 7892 10716 7956
rect 10732 7892 10796 7956
rect 10812 7892 10876 7956
rect 10892 7892 10956 7956
rect 10972 7892 11036 7956
rect 1148 7812 1212 7876
rect 1228 7812 1292 7876
rect 1308 7812 1372 7876
rect 1388 7812 1452 7876
rect 1468 7812 1532 7876
rect 1548 7812 1612 7876
rect 1628 7812 1692 7876
rect 1708 7812 1772 7876
rect 1788 7812 1852 7876
rect 1868 7812 1932 7876
rect 4013 7812 4077 7876
rect 4093 7812 4157 7876
rect 4173 7812 4237 7876
rect 4253 7812 4317 7876
rect 4333 7812 4397 7876
rect 5944 7812 6008 7876
rect 6024 7812 6088 7876
rect 6104 7812 6168 7876
rect 6184 7812 6248 7876
rect 6264 7812 6328 7876
rect 7874 7812 7938 7876
rect 7954 7812 8018 7876
rect 8034 7812 8098 7876
rect 8114 7812 8178 7876
rect 8194 7812 8258 7876
rect 10252 7812 10316 7876
rect 10332 7812 10396 7876
rect 10412 7812 10476 7876
rect 10492 7812 10556 7876
rect 10572 7812 10636 7876
rect 10652 7812 10716 7876
rect 10732 7812 10796 7876
rect 10812 7812 10876 7876
rect 10892 7812 10956 7876
rect 10972 7812 11036 7876
rect 4013 6532 4077 6536
rect 4013 6476 4017 6532
rect 4017 6476 4073 6532
rect 4073 6476 4077 6532
rect 4013 6472 4077 6476
rect 4093 6532 4157 6536
rect 4093 6476 4097 6532
rect 4097 6476 4153 6532
rect 4153 6476 4157 6532
rect 4093 6472 4157 6476
rect 4173 6532 4237 6536
rect 4173 6476 4177 6532
rect 4177 6476 4233 6532
rect 4233 6476 4237 6532
rect 4173 6472 4237 6476
rect 4253 6532 4317 6536
rect 4253 6476 4257 6532
rect 4257 6476 4313 6532
rect 4313 6476 4317 6532
rect 4253 6472 4317 6476
rect 4333 6532 4397 6536
rect 4333 6476 4337 6532
rect 4337 6476 4393 6532
rect 4393 6476 4397 6532
rect 4333 6472 4397 6476
rect 5944 6532 6008 6536
rect 5944 6476 5948 6532
rect 5948 6476 6004 6532
rect 6004 6476 6008 6532
rect 5944 6472 6008 6476
rect 6024 6532 6088 6536
rect 6024 6476 6028 6532
rect 6028 6476 6084 6532
rect 6084 6476 6088 6532
rect 6024 6472 6088 6476
rect 6104 6532 6168 6536
rect 6104 6476 6108 6532
rect 6108 6476 6164 6532
rect 6164 6476 6168 6532
rect 6104 6472 6168 6476
rect 6184 6532 6248 6536
rect 6184 6476 6188 6532
rect 6188 6476 6244 6532
rect 6244 6476 6248 6532
rect 6184 6472 6248 6476
rect 6264 6532 6328 6536
rect 6264 6476 6268 6532
rect 6268 6476 6324 6532
rect 6324 6476 6328 6532
rect 6264 6472 6328 6476
rect 7874 6532 7938 6536
rect 7874 6476 7878 6532
rect 7878 6476 7934 6532
rect 7934 6476 7938 6532
rect 7874 6472 7938 6476
rect 7954 6532 8018 6536
rect 7954 6476 7958 6532
rect 7958 6476 8014 6532
rect 8014 6476 8018 6532
rect 7954 6472 8018 6476
rect 8034 6532 8098 6536
rect 8034 6476 8038 6532
rect 8038 6476 8094 6532
rect 8094 6476 8098 6532
rect 8034 6472 8098 6476
rect 8114 6532 8178 6536
rect 8114 6476 8118 6532
rect 8118 6476 8174 6532
rect 8174 6476 8178 6532
rect 8114 6472 8178 6476
rect 8194 6532 8258 6536
rect 8194 6476 8198 6532
rect 8198 6476 8254 6532
rect 8254 6476 8258 6532
rect 8194 6472 8258 6476
rect 4978 5988 5042 5992
rect 4978 5932 4982 5988
rect 4982 5932 5038 5988
rect 5038 5932 5042 5988
rect 4978 5928 5042 5932
rect 5058 5988 5122 5992
rect 5058 5932 5062 5988
rect 5062 5932 5118 5988
rect 5118 5932 5122 5988
rect 5058 5928 5122 5932
rect 5138 5988 5202 5992
rect 5138 5932 5142 5988
rect 5142 5932 5198 5988
rect 5198 5932 5202 5988
rect 5138 5928 5202 5932
rect 5218 5988 5282 5992
rect 5218 5932 5222 5988
rect 5222 5932 5278 5988
rect 5278 5932 5282 5988
rect 5218 5928 5282 5932
rect 5298 5988 5362 5992
rect 5298 5932 5302 5988
rect 5302 5932 5358 5988
rect 5358 5932 5362 5988
rect 5298 5928 5362 5932
rect 6909 5988 6973 5992
rect 6909 5932 6913 5988
rect 6913 5932 6969 5988
rect 6969 5932 6973 5988
rect 6909 5928 6973 5932
rect 6989 5988 7053 5992
rect 6989 5932 6993 5988
rect 6993 5932 7049 5988
rect 7049 5932 7053 5988
rect 6989 5928 7053 5932
rect 7069 5988 7133 5992
rect 7069 5932 7073 5988
rect 7073 5932 7129 5988
rect 7129 5932 7133 5988
rect 7069 5928 7133 5932
rect 7149 5988 7213 5992
rect 7149 5932 7153 5988
rect 7153 5932 7209 5988
rect 7209 5932 7213 5988
rect 7149 5928 7213 5932
rect 7229 5988 7293 5992
rect 7229 5932 7233 5988
rect 7233 5932 7289 5988
rect 7289 5932 7293 5988
rect 7229 5928 7293 5932
rect 4013 5444 4077 5448
rect 4013 5388 4017 5444
rect 4017 5388 4073 5444
rect 4073 5388 4077 5444
rect 4013 5384 4077 5388
rect 4093 5444 4157 5448
rect 4093 5388 4097 5444
rect 4097 5388 4153 5444
rect 4153 5388 4157 5444
rect 4093 5384 4157 5388
rect 4173 5444 4237 5448
rect 4173 5388 4177 5444
rect 4177 5388 4233 5444
rect 4233 5388 4237 5444
rect 4173 5384 4237 5388
rect 4253 5444 4317 5448
rect 4253 5388 4257 5444
rect 4257 5388 4313 5444
rect 4313 5388 4317 5444
rect 4253 5384 4317 5388
rect 4333 5444 4397 5448
rect 4333 5388 4337 5444
rect 4337 5388 4393 5444
rect 4393 5388 4397 5444
rect 4333 5384 4397 5388
rect 5944 5444 6008 5448
rect 5944 5388 5948 5444
rect 5948 5388 6004 5444
rect 6004 5388 6008 5444
rect 5944 5384 6008 5388
rect 6024 5444 6088 5448
rect 6024 5388 6028 5444
rect 6028 5388 6084 5444
rect 6084 5388 6088 5444
rect 6024 5384 6088 5388
rect 6104 5444 6168 5448
rect 6104 5388 6108 5444
rect 6108 5388 6164 5444
rect 6164 5388 6168 5444
rect 6104 5384 6168 5388
rect 6184 5444 6248 5448
rect 6184 5388 6188 5444
rect 6188 5388 6244 5444
rect 6244 5388 6248 5444
rect 6184 5384 6248 5388
rect 6264 5444 6328 5448
rect 6264 5388 6268 5444
rect 6268 5388 6324 5444
rect 6324 5388 6328 5444
rect 6264 5384 6328 5388
rect 7874 5444 7938 5448
rect 7874 5388 7878 5444
rect 7878 5388 7934 5444
rect 7934 5388 7938 5444
rect 7874 5384 7938 5388
rect 7954 5444 8018 5448
rect 7954 5388 7958 5444
rect 7958 5388 8014 5444
rect 8014 5388 8018 5444
rect 7954 5384 8018 5388
rect 8034 5444 8098 5448
rect 8034 5388 8038 5444
rect 8038 5388 8094 5444
rect 8094 5388 8098 5444
rect 8034 5384 8098 5388
rect 8114 5444 8178 5448
rect 8114 5388 8118 5444
rect 8118 5388 8174 5444
rect 8174 5388 8178 5444
rect 8114 5384 8178 5388
rect 8194 5444 8258 5448
rect 8194 5388 8198 5444
rect 8198 5388 8254 5444
rect 8254 5388 8258 5444
rect 8194 5384 8258 5388
rect 4978 4900 5042 4904
rect 4978 4844 4982 4900
rect 4982 4844 5038 4900
rect 5038 4844 5042 4900
rect 4978 4840 5042 4844
rect 5058 4900 5122 4904
rect 5058 4844 5062 4900
rect 5062 4844 5118 4900
rect 5118 4844 5122 4900
rect 5058 4840 5122 4844
rect 5138 4900 5202 4904
rect 5138 4844 5142 4900
rect 5142 4844 5198 4900
rect 5198 4844 5202 4900
rect 5138 4840 5202 4844
rect 5218 4900 5282 4904
rect 5218 4844 5222 4900
rect 5222 4844 5278 4900
rect 5278 4844 5282 4900
rect 5218 4840 5282 4844
rect 5298 4900 5362 4904
rect 5298 4844 5302 4900
rect 5302 4844 5358 4900
rect 5358 4844 5362 4900
rect 5298 4840 5362 4844
rect 6909 4900 6973 4904
rect 6909 4844 6913 4900
rect 6913 4844 6969 4900
rect 6969 4844 6973 4900
rect 6909 4840 6973 4844
rect 6989 4900 7053 4904
rect 6989 4844 6993 4900
rect 6993 4844 7049 4900
rect 7049 4844 7053 4900
rect 6989 4840 7053 4844
rect 7069 4900 7133 4904
rect 7069 4844 7073 4900
rect 7073 4844 7129 4900
rect 7129 4844 7133 4900
rect 7069 4840 7133 4844
rect 7149 4900 7213 4904
rect 7149 4844 7153 4900
rect 7153 4844 7209 4900
rect 7209 4844 7213 4900
rect 7149 4840 7213 4844
rect 7229 4900 7293 4904
rect 7229 4844 7233 4900
rect 7233 4844 7289 4900
rect 7289 4844 7293 4900
rect 7229 4840 7293 4844
rect 4013 4356 4077 4360
rect 4013 4300 4017 4356
rect 4017 4300 4073 4356
rect 4073 4300 4077 4356
rect 4013 4296 4077 4300
rect 4093 4356 4157 4360
rect 4093 4300 4097 4356
rect 4097 4300 4153 4356
rect 4153 4300 4157 4356
rect 4093 4296 4157 4300
rect 4173 4356 4237 4360
rect 4173 4300 4177 4356
rect 4177 4300 4233 4356
rect 4233 4300 4237 4356
rect 4173 4296 4237 4300
rect 4253 4356 4317 4360
rect 4253 4300 4257 4356
rect 4257 4300 4313 4356
rect 4313 4300 4317 4356
rect 4253 4296 4317 4300
rect 4333 4356 4397 4360
rect 4333 4300 4337 4356
rect 4337 4300 4393 4356
rect 4393 4300 4397 4356
rect 4333 4296 4397 4300
rect 5944 4356 6008 4360
rect 5944 4300 5948 4356
rect 5948 4300 6004 4356
rect 6004 4300 6008 4356
rect 5944 4296 6008 4300
rect 6024 4356 6088 4360
rect 6024 4300 6028 4356
rect 6028 4300 6084 4356
rect 6084 4300 6088 4356
rect 6024 4296 6088 4300
rect 6104 4356 6168 4360
rect 6104 4300 6108 4356
rect 6108 4300 6164 4356
rect 6164 4300 6168 4356
rect 6104 4296 6168 4300
rect 6184 4356 6248 4360
rect 6184 4300 6188 4356
rect 6188 4300 6244 4356
rect 6244 4300 6248 4356
rect 6184 4296 6248 4300
rect 6264 4356 6328 4360
rect 6264 4300 6268 4356
rect 6268 4300 6324 4356
rect 6324 4300 6328 4356
rect 6264 4296 6328 4300
rect 7874 4356 7938 4360
rect 7874 4300 7878 4356
rect 7878 4300 7934 4356
rect 7934 4300 7938 4356
rect 7874 4296 7938 4300
rect 7954 4356 8018 4360
rect 7954 4300 7958 4356
rect 7958 4300 8014 4356
rect 8014 4300 8018 4356
rect 7954 4296 8018 4300
rect 8034 4356 8098 4360
rect 8034 4300 8038 4356
rect 8038 4300 8094 4356
rect 8094 4300 8098 4356
rect 8034 4296 8098 4300
rect 8114 4356 8178 4360
rect 8114 4300 8118 4356
rect 8118 4300 8174 4356
rect 8174 4300 8178 4356
rect 8114 4296 8178 4300
rect 8194 4356 8258 4360
rect 8194 4300 8198 4356
rect 8198 4300 8254 4356
rect 8254 4300 8258 4356
rect 8194 4296 8258 4300
rect 4978 3812 5042 3816
rect 4978 3756 4982 3812
rect 4982 3756 5038 3812
rect 5038 3756 5042 3812
rect 4978 3752 5042 3756
rect 5058 3812 5122 3816
rect 5058 3756 5062 3812
rect 5062 3756 5118 3812
rect 5118 3756 5122 3812
rect 5058 3752 5122 3756
rect 5138 3812 5202 3816
rect 5138 3756 5142 3812
rect 5142 3756 5198 3812
rect 5198 3756 5202 3812
rect 5138 3752 5202 3756
rect 5218 3812 5282 3816
rect 5218 3756 5222 3812
rect 5222 3756 5278 3812
rect 5278 3756 5282 3812
rect 5218 3752 5282 3756
rect 5298 3812 5362 3816
rect 5298 3756 5302 3812
rect 5302 3756 5358 3812
rect 5358 3756 5362 3812
rect 5298 3752 5362 3756
rect 6909 3812 6973 3816
rect 6909 3756 6913 3812
rect 6913 3756 6969 3812
rect 6969 3756 6973 3812
rect 6909 3752 6973 3756
rect 6989 3812 7053 3816
rect 6989 3756 6993 3812
rect 6993 3756 7049 3812
rect 7049 3756 7053 3812
rect 6989 3752 7053 3756
rect 7069 3812 7133 3816
rect 7069 3756 7073 3812
rect 7073 3756 7129 3812
rect 7129 3756 7133 3812
rect 7069 3752 7133 3756
rect 7149 3812 7213 3816
rect 7149 3756 7153 3812
rect 7153 3756 7209 3812
rect 7209 3756 7213 3812
rect 7149 3752 7213 3756
rect 7229 3812 7293 3816
rect 7229 3756 7233 3812
rect 7233 3756 7289 3812
rect 7289 3756 7293 3812
rect 7229 3752 7293 3756
rect 4013 3268 4077 3272
rect 4013 3212 4017 3268
rect 4017 3212 4073 3268
rect 4073 3212 4077 3268
rect 4013 3208 4077 3212
rect 4093 3268 4157 3272
rect 4093 3212 4097 3268
rect 4097 3212 4153 3268
rect 4153 3212 4157 3268
rect 4093 3208 4157 3212
rect 4173 3268 4237 3272
rect 4173 3212 4177 3268
rect 4177 3212 4233 3268
rect 4233 3212 4237 3268
rect 4173 3208 4237 3212
rect 4253 3268 4317 3272
rect 4253 3212 4257 3268
rect 4257 3212 4313 3268
rect 4313 3212 4317 3268
rect 4253 3208 4317 3212
rect 4333 3268 4397 3272
rect 4333 3212 4337 3268
rect 4337 3212 4393 3268
rect 4393 3212 4397 3268
rect 4333 3208 4397 3212
rect 5944 3268 6008 3272
rect 5944 3212 5948 3268
rect 5948 3212 6004 3268
rect 6004 3212 6008 3268
rect 5944 3208 6008 3212
rect 6024 3268 6088 3272
rect 6024 3212 6028 3268
rect 6028 3212 6084 3268
rect 6084 3212 6088 3268
rect 6024 3208 6088 3212
rect 6104 3268 6168 3272
rect 6104 3212 6108 3268
rect 6108 3212 6164 3268
rect 6164 3212 6168 3268
rect 6104 3208 6168 3212
rect 6184 3268 6248 3272
rect 6184 3212 6188 3268
rect 6188 3212 6244 3268
rect 6244 3212 6248 3268
rect 6184 3208 6248 3212
rect 6264 3268 6328 3272
rect 6264 3212 6268 3268
rect 6268 3212 6324 3268
rect 6324 3212 6328 3268
rect 6264 3208 6328 3212
rect 7874 3268 7938 3272
rect 7874 3212 7878 3268
rect 7878 3212 7934 3268
rect 7934 3212 7938 3268
rect 7874 3208 7938 3212
rect 7954 3268 8018 3272
rect 7954 3212 7958 3268
rect 7958 3212 8014 3268
rect 8014 3212 8018 3268
rect 7954 3208 8018 3212
rect 8034 3268 8098 3272
rect 8034 3212 8038 3268
rect 8038 3212 8094 3268
rect 8094 3212 8098 3268
rect 8034 3208 8098 3212
rect 8114 3268 8178 3272
rect 8114 3212 8118 3268
rect 8118 3212 8174 3268
rect 8174 3212 8178 3268
rect 8114 3208 8178 3212
rect 8194 3268 8258 3272
rect 8194 3212 8198 3268
rect 8198 3212 8254 3268
rect 8254 3212 8258 3268
rect 8194 3208 8258 3212
rect 1148 1868 1212 1932
rect 1228 1868 1292 1932
rect 1308 1868 1372 1932
rect 1388 1868 1452 1932
rect 1468 1868 1532 1932
rect 1548 1868 1612 1932
rect 1628 1868 1692 1932
rect 1708 1868 1772 1932
rect 1788 1868 1852 1932
rect 1868 1868 1932 1932
rect 4013 1868 4077 1932
rect 4093 1868 4157 1932
rect 4173 1868 4237 1932
rect 4253 1868 4317 1932
rect 4333 1868 4397 1932
rect 5944 1868 6008 1932
rect 6024 1868 6088 1932
rect 6104 1868 6168 1932
rect 6184 1868 6248 1932
rect 6264 1868 6328 1932
rect 7874 1868 7938 1932
rect 7954 1868 8018 1932
rect 8034 1868 8098 1932
rect 8114 1868 8178 1932
rect 8194 1868 8258 1932
rect 10252 1868 10316 1932
rect 10332 1868 10396 1932
rect 10412 1868 10476 1932
rect 10492 1868 10556 1932
rect 10572 1868 10636 1932
rect 10652 1868 10716 1932
rect 10732 1868 10796 1932
rect 10812 1868 10876 1932
rect 10892 1868 10956 1932
rect 10972 1868 11036 1932
rect 1148 1788 1212 1852
rect 1228 1788 1292 1852
rect 1308 1788 1372 1852
rect 1388 1788 1452 1852
rect 1468 1788 1532 1852
rect 1548 1788 1612 1852
rect 1628 1788 1692 1852
rect 1708 1788 1772 1852
rect 1788 1788 1852 1852
rect 1868 1788 1932 1852
rect 4013 1788 4077 1852
rect 4093 1788 4157 1852
rect 4173 1788 4237 1852
rect 4253 1788 4317 1852
rect 4333 1788 4397 1852
rect 5944 1788 6008 1852
rect 6024 1788 6088 1852
rect 6104 1788 6168 1852
rect 6184 1788 6248 1852
rect 6264 1788 6328 1852
rect 7874 1788 7938 1852
rect 7954 1788 8018 1852
rect 8034 1788 8098 1852
rect 8114 1788 8178 1852
rect 8194 1788 8258 1852
rect 10252 1788 10316 1852
rect 10332 1788 10396 1852
rect 10412 1788 10476 1852
rect 10492 1788 10556 1852
rect 10572 1788 10636 1852
rect 10652 1788 10716 1852
rect 10732 1788 10796 1852
rect 10812 1788 10876 1852
rect 10892 1788 10956 1852
rect 10972 1788 11036 1852
rect 1148 1708 1212 1772
rect 1228 1708 1292 1772
rect 1308 1708 1372 1772
rect 1388 1708 1452 1772
rect 1468 1708 1532 1772
rect 1548 1708 1612 1772
rect 1628 1708 1692 1772
rect 1708 1708 1772 1772
rect 1788 1708 1852 1772
rect 1868 1708 1932 1772
rect 4013 1708 4077 1772
rect 4093 1708 4157 1772
rect 4173 1708 4237 1772
rect 4253 1708 4317 1772
rect 4333 1708 4397 1772
rect 5944 1708 6008 1772
rect 6024 1708 6088 1772
rect 6104 1708 6168 1772
rect 6184 1708 6248 1772
rect 6264 1708 6328 1772
rect 7874 1708 7938 1772
rect 7954 1708 8018 1772
rect 8034 1708 8098 1772
rect 8114 1708 8178 1772
rect 8194 1708 8258 1772
rect 10252 1708 10316 1772
rect 10332 1708 10396 1772
rect 10412 1708 10476 1772
rect 10492 1708 10556 1772
rect 10572 1708 10636 1772
rect 10652 1708 10716 1772
rect 10732 1708 10796 1772
rect 10812 1708 10876 1772
rect 10892 1708 10956 1772
rect 10972 1708 11036 1772
rect 1148 1628 1212 1692
rect 1228 1628 1292 1692
rect 1308 1628 1372 1692
rect 1388 1628 1452 1692
rect 1468 1628 1532 1692
rect 1548 1628 1612 1692
rect 1628 1628 1692 1692
rect 1708 1628 1772 1692
rect 1788 1628 1852 1692
rect 1868 1628 1932 1692
rect 4013 1628 4077 1692
rect 4093 1628 4157 1692
rect 4173 1628 4237 1692
rect 4253 1628 4317 1692
rect 4333 1628 4397 1692
rect 5944 1628 6008 1692
rect 6024 1628 6088 1692
rect 6104 1628 6168 1692
rect 6184 1628 6248 1692
rect 6264 1628 6328 1692
rect 7874 1628 7938 1692
rect 7954 1628 8018 1692
rect 8034 1628 8098 1692
rect 8114 1628 8178 1692
rect 8194 1628 8258 1692
rect 10252 1628 10316 1692
rect 10332 1628 10396 1692
rect 10412 1628 10476 1692
rect 10492 1628 10556 1692
rect 10572 1628 10636 1692
rect 10652 1628 10716 1692
rect 10732 1628 10796 1692
rect 10812 1628 10876 1692
rect 10892 1628 10956 1692
rect 10972 1628 11036 1692
rect 1148 1548 1212 1612
rect 1228 1548 1292 1612
rect 1308 1548 1372 1612
rect 1388 1548 1452 1612
rect 1468 1548 1532 1612
rect 1548 1548 1612 1612
rect 1628 1548 1692 1612
rect 1708 1548 1772 1612
rect 1788 1548 1852 1612
rect 1868 1548 1932 1612
rect 4013 1548 4077 1612
rect 4093 1548 4157 1612
rect 4173 1548 4237 1612
rect 4253 1548 4317 1612
rect 4333 1548 4397 1612
rect 5944 1548 6008 1612
rect 6024 1548 6088 1612
rect 6104 1548 6168 1612
rect 6184 1548 6248 1612
rect 6264 1548 6328 1612
rect 7874 1548 7938 1612
rect 7954 1548 8018 1612
rect 8034 1548 8098 1612
rect 8114 1548 8178 1612
rect 8194 1548 8258 1612
rect 10252 1548 10316 1612
rect 10332 1548 10396 1612
rect 10412 1548 10476 1612
rect 10492 1548 10556 1612
rect 10572 1548 10636 1612
rect 10652 1548 10716 1612
rect 10732 1548 10796 1612
rect 10812 1548 10876 1612
rect 10892 1548 10956 1612
rect 10972 1548 11036 1612
rect 1148 1468 1212 1532
rect 1228 1468 1292 1532
rect 1308 1468 1372 1532
rect 1388 1468 1452 1532
rect 1468 1468 1532 1532
rect 1548 1468 1612 1532
rect 1628 1468 1692 1532
rect 1708 1468 1772 1532
rect 1788 1468 1852 1532
rect 1868 1468 1932 1532
rect 4013 1468 4077 1532
rect 4093 1468 4157 1532
rect 4173 1468 4237 1532
rect 4253 1468 4317 1532
rect 4333 1468 4397 1532
rect 5944 1468 6008 1532
rect 6024 1468 6088 1532
rect 6104 1468 6168 1532
rect 6184 1468 6248 1532
rect 6264 1468 6328 1532
rect 7874 1468 7938 1532
rect 7954 1468 8018 1532
rect 8034 1468 8098 1532
rect 8114 1468 8178 1532
rect 8194 1468 8258 1532
rect 10252 1468 10316 1532
rect 10332 1468 10396 1532
rect 10412 1468 10476 1532
rect 10492 1468 10556 1532
rect 10572 1468 10636 1532
rect 10652 1468 10716 1532
rect 10732 1468 10796 1532
rect 10812 1468 10876 1532
rect 10892 1468 10956 1532
rect 10972 1468 11036 1532
rect 1148 1388 1212 1452
rect 1228 1388 1292 1452
rect 1308 1388 1372 1452
rect 1388 1388 1452 1452
rect 1468 1388 1532 1452
rect 1548 1388 1612 1452
rect 1628 1388 1692 1452
rect 1708 1388 1772 1452
rect 1788 1388 1852 1452
rect 1868 1388 1932 1452
rect 4013 1388 4077 1452
rect 4093 1388 4157 1452
rect 4173 1388 4237 1452
rect 4253 1388 4317 1452
rect 4333 1388 4397 1452
rect 5944 1388 6008 1452
rect 6024 1388 6088 1452
rect 6104 1388 6168 1452
rect 6184 1388 6248 1452
rect 6264 1388 6328 1452
rect 7874 1388 7938 1452
rect 7954 1388 8018 1452
rect 8034 1388 8098 1452
rect 8114 1388 8178 1452
rect 8194 1388 8258 1452
rect 10252 1388 10316 1452
rect 10332 1388 10396 1452
rect 10412 1388 10476 1452
rect 10492 1388 10556 1452
rect 10572 1388 10636 1452
rect 10652 1388 10716 1452
rect 10732 1388 10796 1452
rect 10812 1388 10876 1452
rect 10892 1388 10956 1452
rect 10972 1388 11036 1452
rect 1148 1308 1212 1372
rect 1228 1308 1292 1372
rect 1308 1308 1372 1372
rect 1388 1308 1452 1372
rect 1468 1308 1532 1372
rect 1548 1308 1612 1372
rect 1628 1308 1692 1372
rect 1708 1308 1772 1372
rect 1788 1308 1852 1372
rect 1868 1308 1932 1372
rect 4013 1308 4077 1372
rect 4093 1308 4157 1372
rect 4173 1308 4237 1372
rect 4253 1308 4317 1372
rect 4333 1308 4397 1372
rect 5944 1308 6008 1372
rect 6024 1308 6088 1372
rect 6104 1308 6168 1372
rect 6184 1308 6248 1372
rect 6264 1308 6328 1372
rect 7874 1308 7938 1372
rect 7954 1308 8018 1372
rect 8034 1308 8098 1372
rect 8114 1308 8178 1372
rect 8194 1308 8258 1372
rect 10252 1308 10316 1372
rect 10332 1308 10396 1372
rect 10412 1308 10476 1372
rect 10492 1308 10556 1372
rect 10572 1308 10636 1372
rect 10652 1308 10716 1372
rect 10732 1308 10796 1372
rect 10812 1308 10876 1372
rect 10892 1308 10956 1372
rect 10972 1308 11036 1372
rect 1148 1228 1212 1292
rect 1228 1228 1292 1292
rect 1308 1228 1372 1292
rect 1388 1228 1452 1292
rect 1468 1228 1532 1292
rect 1548 1228 1612 1292
rect 1628 1228 1692 1292
rect 1708 1228 1772 1292
rect 1788 1228 1852 1292
rect 1868 1228 1932 1292
rect 4013 1228 4077 1292
rect 4093 1228 4157 1292
rect 4173 1228 4237 1292
rect 4253 1228 4317 1292
rect 4333 1228 4397 1292
rect 5944 1228 6008 1292
rect 6024 1228 6088 1292
rect 6104 1228 6168 1292
rect 6184 1228 6248 1292
rect 6264 1228 6328 1292
rect 7874 1228 7938 1292
rect 7954 1228 8018 1292
rect 8034 1228 8098 1292
rect 8114 1228 8178 1292
rect 8194 1228 8258 1292
rect 10252 1228 10316 1292
rect 10332 1228 10396 1292
rect 10412 1228 10476 1292
rect 10492 1228 10556 1292
rect 10572 1228 10636 1292
rect 10652 1228 10716 1292
rect 10732 1228 10796 1292
rect 10812 1228 10876 1292
rect 10892 1228 10956 1292
rect 10972 1228 11036 1292
rect 1148 1148 1212 1212
rect 1228 1148 1292 1212
rect 1308 1148 1372 1212
rect 1388 1148 1452 1212
rect 1468 1148 1532 1212
rect 1548 1148 1612 1212
rect 1628 1148 1692 1212
rect 1708 1148 1772 1212
rect 1788 1148 1852 1212
rect 1868 1148 1932 1212
rect 4013 1148 4077 1212
rect 4093 1148 4157 1212
rect 4173 1148 4237 1212
rect 4253 1148 4317 1212
rect 4333 1148 4397 1212
rect 5944 1148 6008 1212
rect 6024 1148 6088 1212
rect 6104 1148 6168 1212
rect 6184 1148 6248 1212
rect 6264 1148 6328 1212
rect 7874 1148 7938 1212
rect 7954 1148 8018 1212
rect 8034 1148 8098 1212
rect 8114 1148 8178 1212
rect 8194 1148 8258 1212
rect 10252 1148 10316 1212
rect 10332 1148 10396 1212
rect 10412 1148 10476 1212
rect 10492 1148 10556 1212
rect 10572 1148 10636 1212
rect 10652 1148 10716 1212
rect 10732 1148 10796 1212
rect 10812 1148 10876 1212
rect 10892 1148 10956 1212
rect 10972 1148 11036 1212
rect 8 728 72 792
rect 88 728 152 792
rect 168 728 232 792
rect 248 728 312 792
rect 328 728 392 792
rect 408 728 472 792
rect 488 728 552 792
rect 568 728 632 792
rect 648 728 712 792
rect 728 728 792 792
rect 4978 728 5042 792
rect 5058 728 5122 792
rect 5138 728 5202 792
rect 5218 728 5282 792
rect 5298 728 5362 792
rect 6909 728 6973 792
rect 6989 728 7053 792
rect 7069 728 7133 792
rect 7149 728 7213 792
rect 7229 728 7293 792
rect 11392 728 11456 792
rect 11472 728 11536 792
rect 11552 728 11616 792
rect 11632 728 11696 792
rect 11712 728 11776 792
rect 11792 728 11856 792
rect 11872 728 11936 792
rect 11952 728 12016 792
rect 12032 728 12096 792
rect 12112 728 12176 792
rect 8 648 72 712
rect 88 648 152 712
rect 168 648 232 712
rect 248 648 312 712
rect 328 648 392 712
rect 408 648 472 712
rect 488 648 552 712
rect 568 648 632 712
rect 648 648 712 712
rect 728 648 792 712
rect 4978 648 5042 712
rect 5058 648 5122 712
rect 5138 648 5202 712
rect 5218 648 5282 712
rect 5298 648 5362 712
rect 6909 648 6973 712
rect 6989 648 7053 712
rect 7069 648 7133 712
rect 7149 648 7213 712
rect 7229 648 7293 712
rect 11392 648 11456 712
rect 11472 648 11536 712
rect 11552 648 11616 712
rect 11632 648 11696 712
rect 11712 648 11776 712
rect 11792 648 11856 712
rect 11872 648 11936 712
rect 11952 648 12016 712
rect 12032 648 12096 712
rect 12112 648 12176 712
rect 8 568 72 632
rect 88 568 152 632
rect 168 568 232 632
rect 248 568 312 632
rect 328 568 392 632
rect 408 568 472 632
rect 488 568 552 632
rect 568 568 632 632
rect 648 568 712 632
rect 728 568 792 632
rect 4978 568 5042 632
rect 5058 568 5122 632
rect 5138 568 5202 632
rect 5218 568 5282 632
rect 5298 568 5362 632
rect 6909 568 6973 632
rect 6989 568 7053 632
rect 7069 568 7133 632
rect 7149 568 7213 632
rect 7229 568 7293 632
rect 11392 568 11456 632
rect 11472 568 11536 632
rect 11552 568 11616 632
rect 11632 568 11696 632
rect 11712 568 11776 632
rect 11792 568 11856 632
rect 11872 568 11936 632
rect 11952 568 12016 632
rect 12032 568 12096 632
rect 12112 568 12176 632
rect 8 488 72 552
rect 88 488 152 552
rect 168 488 232 552
rect 248 488 312 552
rect 328 488 392 552
rect 408 488 472 552
rect 488 488 552 552
rect 568 488 632 552
rect 648 488 712 552
rect 728 488 792 552
rect 4978 488 5042 552
rect 5058 488 5122 552
rect 5138 488 5202 552
rect 5218 488 5282 552
rect 5298 488 5362 552
rect 6909 488 6973 552
rect 6989 488 7053 552
rect 7069 488 7133 552
rect 7149 488 7213 552
rect 7229 488 7293 552
rect 11392 488 11456 552
rect 11472 488 11536 552
rect 11552 488 11616 552
rect 11632 488 11696 552
rect 11712 488 11776 552
rect 11792 488 11856 552
rect 11872 488 11936 552
rect 11952 488 12016 552
rect 12032 488 12096 552
rect 12112 488 12176 552
rect 8 408 72 472
rect 88 408 152 472
rect 168 408 232 472
rect 248 408 312 472
rect 328 408 392 472
rect 408 408 472 472
rect 488 408 552 472
rect 568 408 632 472
rect 648 408 712 472
rect 728 408 792 472
rect 4978 408 5042 472
rect 5058 408 5122 472
rect 5138 408 5202 472
rect 5218 408 5282 472
rect 5298 408 5362 472
rect 6909 408 6973 472
rect 6989 408 7053 472
rect 7069 408 7133 472
rect 7149 408 7213 472
rect 7229 408 7293 472
rect 11392 408 11456 472
rect 11472 408 11536 472
rect 11552 408 11616 472
rect 11632 408 11696 472
rect 11712 408 11776 472
rect 11792 408 11856 472
rect 11872 408 11936 472
rect 11952 408 12016 472
rect 12032 408 12096 472
rect 12112 408 12176 472
rect 8 328 72 392
rect 88 328 152 392
rect 168 328 232 392
rect 248 328 312 392
rect 328 328 392 392
rect 408 328 472 392
rect 488 328 552 392
rect 568 328 632 392
rect 648 328 712 392
rect 728 328 792 392
rect 4978 328 5042 392
rect 5058 328 5122 392
rect 5138 328 5202 392
rect 5218 328 5282 392
rect 5298 328 5362 392
rect 6909 328 6973 392
rect 6989 328 7053 392
rect 7069 328 7133 392
rect 7149 328 7213 392
rect 7229 328 7293 392
rect 11392 328 11456 392
rect 11472 328 11536 392
rect 11552 328 11616 392
rect 11632 328 11696 392
rect 11712 328 11776 392
rect 11792 328 11856 392
rect 11872 328 11936 392
rect 11952 328 12016 392
rect 12032 328 12096 392
rect 12112 328 12176 392
rect 8 248 72 312
rect 88 248 152 312
rect 168 248 232 312
rect 248 248 312 312
rect 328 248 392 312
rect 408 248 472 312
rect 488 248 552 312
rect 568 248 632 312
rect 648 248 712 312
rect 728 248 792 312
rect 4978 248 5042 312
rect 5058 248 5122 312
rect 5138 248 5202 312
rect 5218 248 5282 312
rect 5298 248 5362 312
rect 6909 248 6973 312
rect 6989 248 7053 312
rect 7069 248 7133 312
rect 7149 248 7213 312
rect 7229 248 7293 312
rect 11392 248 11456 312
rect 11472 248 11536 312
rect 11552 248 11616 312
rect 11632 248 11696 312
rect 11712 248 11776 312
rect 11792 248 11856 312
rect 11872 248 11936 312
rect 11952 248 12016 312
rect 12032 248 12096 312
rect 12112 248 12176 312
rect 8 168 72 232
rect 88 168 152 232
rect 168 168 232 232
rect 248 168 312 232
rect 328 168 392 232
rect 408 168 472 232
rect 488 168 552 232
rect 568 168 632 232
rect 648 168 712 232
rect 728 168 792 232
rect 4978 168 5042 232
rect 5058 168 5122 232
rect 5138 168 5202 232
rect 5218 168 5282 232
rect 5298 168 5362 232
rect 6909 168 6973 232
rect 6989 168 7053 232
rect 7069 168 7133 232
rect 7149 168 7213 232
rect 7229 168 7293 232
rect 11392 168 11456 232
rect 11472 168 11536 232
rect 11552 168 11616 232
rect 11632 168 11696 232
rect 11712 168 11776 232
rect 11792 168 11856 232
rect 11872 168 11936 232
rect 11952 168 12016 232
rect 12032 168 12096 232
rect 12112 168 12176 232
rect 8 88 72 152
rect 88 88 152 152
rect 168 88 232 152
rect 248 88 312 152
rect 328 88 392 152
rect 408 88 472 152
rect 488 88 552 152
rect 568 88 632 152
rect 648 88 712 152
rect 728 88 792 152
rect 4978 88 5042 152
rect 5058 88 5122 152
rect 5138 88 5202 152
rect 5218 88 5282 152
rect 5298 88 5362 152
rect 6909 88 6973 152
rect 6989 88 7053 152
rect 7069 88 7133 152
rect 7149 88 7213 152
rect 7229 88 7293 152
rect 11392 88 11456 152
rect 11472 88 11536 152
rect 11552 88 11616 152
rect 11632 88 11696 152
rect 11712 88 11776 152
rect 11792 88 11856 152
rect 11872 88 11936 152
rect 11952 88 12016 152
rect 12032 88 12096 152
rect 12112 88 12176 152
rect 8 8 72 72
rect 88 8 152 72
rect 168 8 232 72
rect 248 8 312 72
rect 328 8 392 72
rect 408 8 472 72
rect 488 8 552 72
rect 568 8 632 72
rect 648 8 712 72
rect 728 8 792 72
rect 4978 8 5042 72
rect 5058 8 5122 72
rect 5138 8 5202 72
rect 5218 8 5282 72
rect 5298 8 5362 72
rect 6909 8 6973 72
rect 6989 8 7053 72
rect 7069 8 7133 72
rect 7149 8 7213 72
rect 7229 8 7293 72
rect 11392 8 11456 72
rect 11472 8 11536 72
rect 11552 8 11616 72
rect 11632 8 11696 72
rect 11712 8 11776 72
rect 11792 8 11856 72
rect 11872 8 11936 72
rect 11952 8 12016 72
rect 12032 8 12096 72
rect 12112 8 12176 72
<< metal4 >>
rect 0 9736 800 9744
rect 0 9672 8 9736
rect 72 9672 88 9736
rect 152 9672 168 9736
rect 232 9672 248 9736
rect 312 9672 328 9736
rect 392 9672 408 9736
rect 472 9672 488 9736
rect 552 9672 568 9736
rect 632 9672 648 9736
rect 712 9672 728 9736
rect 792 9672 800 9736
rect 0 9656 800 9672
rect 0 9592 8 9656
rect 72 9592 88 9656
rect 152 9592 168 9656
rect 232 9592 248 9656
rect 312 9592 328 9656
rect 392 9592 408 9656
rect 472 9592 488 9656
rect 552 9592 568 9656
rect 632 9592 648 9656
rect 712 9592 728 9656
rect 792 9592 800 9656
rect 0 9576 800 9592
rect 0 9512 8 9576
rect 72 9512 88 9576
rect 152 9512 168 9576
rect 232 9512 248 9576
rect 312 9512 328 9576
rect 392 9512 408 9576
rect 472 9512 488 9576
rect 552 9512 568 9576
rect 632 9512 648 9576
rect 712 9512 728 9576
rect 792 9512 800 9576
rect 0 9496 800 9512
rect 0 9432 8 9496
rect 72 9432 88 9496
rect 152 9432 168 9496
rect 232 9432 248 9496
rect 312 9432 328 9496
rect 392 9432 408 9496
rect 472 9432 488 9496
rect 552 9432 568 9496
rect 632 9432 648 9496
rect 712 9432 728 9496
rect 792 9432 800 9496
rect 0 9416 800 9432
rect 0 9352 8 9416
rect 72 9352 88 9416
rect 152 9352 168 9416
rect 232 9352 248 9416
rect 312 9352 328 9416
rect 392 9352 408 9416
rect 472 9352 488 9416
rect 552 9352 568 9416
rect 632 9352 648 9416
rect 712 9352 728 9416
rect 792 9352 800 9416
rect 0 9336 800 9352
rect 0 9272 8 9336
rect 72 9272 88 9336
rect 152 9272 168 9336
rect 232 9272 248 9336
rect 312 9272 328 9336
rect 392 9272 408 9336
rect 472 9272 488 9336
rect 552 9272 568 9336
rect 632 9272 648 9336
rect 712 9272 728 9336
rect 792 9272 800 9336
rect 0 9256 800 9272
rect 0 9192 8 9256
rect 72 9192 88 9256
rect 152 9192 168 9256
rect 232 9192 248 9256
rect 312 9192 328 9256
rect 392 9192 408 9256
rect 472 9192 488 9256
rect 552 9192 568 9256
rect 632 9192 648 9256
rect 712 9192 728 9256
rect 792 9192 800 9256
rect 0 9176 800 9192
rect 0 9112 8 9176
rect 72 9112 88 9176
rect 152 9112 168 9176
rect 232 9112 248 9176
rect 312 9112 328 9176
rect 392 9112 408 9176
rect 472 9112 488 9176
rect 552 9112 568 9176
rect 632 9112 648 9176
rect 712 9112 728 9176
rect 792 9112 800 9176
rect 0 9096 800 9112
rect 0 9032 8 9096
rect 72 9032 88 9096
rect 152 9032 168 9096
rect 232 9032 248 9096
rect 312 9032 328 9096
rect 392 9032 408 9096
rect 472 9032 488 9096
rect 552 9032 568 9096
rect 632 9032 648 9096
rect 712 9032 728 9096
rect 792 9032 800 9096
rect 0 9016 800 9032
rect 0 8952 8 9016
rect 72 8952 88 9016
rect 152 8952 168 9016
rect 232 8952 248 9016
rect 312 8952 328 9016
rect 392 8952 408 9016
rect 472 8952 488 9016
rect 552 8952 568 9016
rect 632 8952 648 9016
rect 712 8952 728 9016
rect 792 8952 800 9016
rect 0 792 800 8952
rect 1140 8596 1940 8604
rect 1140 8532 1148 8596
rect 1212 8532 1228 8596
rect 1292 8532 1308 8596
rect 1372 8532 1388 8596
rect 1452 8532 1468 8596
rect 1532 8532 1548 8596
rect 1612 8532 1628 8596
rect 1692 8532 1708 8596
rect 1772 8532 1788 8596
rect 1852 8532 1868 8596
rect 1932 8532 1940 8596
rect 1140 8516 1940 8532
rect 1140 8452 1148 8516
rect 1212 8452 1228 8516
rect 1292 8452 1308 8516
rect 1372 8452 1388 8516
rect 1452 8452 1468 8516
rect 1532 8452 1548 8516
rect 1612 8452 1628 8516
rect 1692 8452 1708 8516
rect 1772 8452 1788 8516
rect 1852 8452 1868 8516
rect 1932 8452 1940 8516
rect 1140 8436 1940 8452
rect 1140 8372 1148 8436
rect 1212 8372 1228 8436
rect 1292 8372 1308 8436
rect 1372 8372 1388 8436
rect 1452 8372 1468 8436
rect 1532 8372 1548 8436
rect 1612 8372 1628 8436
rect 1692 8372 1708 8436
rect 1772 8372 1788 8436
rect 1852 8372 1868 8436
rect 1932 8372 1940 8436
rect 1140 8356 1940 8372
rect 1140 8292 1148 8356
rect 1212 8292 1228 8356
rect 1292 8292 1308 8356
rect 1372 8292 1388 8356
rect 1452 8292 1468 8356
rect 1532 8292 1548 8356
rect 1612 8292 1628 8356
rect 1692 8292 1708 8356
rect 1772 8292 1788 8356
rect 1852 8292 1868 8356
rect 1932 8292 1940 8356
rect 1140 8276 1940 8292
rect 1140 8212 1148 8276
rect 1212 8212 1228 8276
rect 1292 8212 1308 8276
rect 1372 8212 1388 8276
rect 1452 8212 1468 8276
rect 1532 8212 1548 8276
rect 1612 8212 1628 8276
rect 1692 8212 1708 8276
rect 1772 8212 1788 8276
rect 1852 8212 1868 8276
rect 1932 8212 1940 8276
rect 1140 8196 1940 8212
rect 1140 8132 1148 8196
rect 1212 8132 1228 8196
rect 1292 8132 1308 8196
rect 1372 8132 1388 8196
rect 1452 8132 1468 8196
rect 1532 8132 1548 8196
rect 1612 8132 1628 8196
rect 1692 8132 1708 8196
rect 1772 8132 1788 8196
rect 1852 8132 1868 8196
rect 1932 8132 1940 8196
rect 1140 8116 1940 8132
rect 1140 8052 1148 8116
rect 1212 8052 1228 8116
rect 1292 8052 1308 8116
rect 1372 8052 1388 8116
rect 1452 8052 1468 8116
rect 1532 8052 1548 8116
rect 1612 8052 1628 8116
rect 1692 8052 1708 8116
rect 1772 8052 1788 8116
rect 1852 8052 1868 8116
rect 1932 8052 1940 8116
rect 1140 8036 1940 8052
rect 1140 7972 1148 8036
rect 1212 7972 1228 8036
rect 1292 7972 1308 8036
rect 1372 7972 1388 8036
rect 1452 7972 1468 8036
rect 1532 7972 1548 8036
rect 1612 7972 1628 8036
rect 1692 7972 1708 8036
rect 1772 7972 1788 8036
rect 1852 7972 1868 8036
rect 1932 7972 1940 8036
rect 1140 7956 1940 7972
rect 1140 7892 1148 7956
rect 1212 7892 1228 7956
rect 1292 7892 1308 7956
rect 1372 7892 1388 7956
rect 1452 7892 1468 7956
rect 1532 7892 1548 7956
rect 1612 7892 1628 7956
rect 1692 7892 1708 7956
rect 1772 7892 1788 7956
rect 1852 7892 1868 7956
rect 1932 7892 1940 7956
rect 1140 7876 1940 7892
rect 1140 7812 1148 7876
rect 1212 7812 1228 7876
rect 1292 7812 1308 7876
rect 1372 7812 1388 7876
rect 1452 7812 1468 7876
rect 1532 7812 1548 7876
rect 1612 7812 1628 7876
rect 1692 7812 1708 7876
rect 1772 7812 1788 7876
rect 1852 7812 1868 7876
rect 1932 7812 1940 7876
rect 1140 1932 1940 7812
rect 1140 1868 1148 1932
rect 1212 1868 1228 1932
rect 1292 1868 1308 1932
rect 1372 1868 1388 1932
rect 1452 1868 1468 1932
rect 1532 1868 1548 1932
rect 1612 1868 1628 1932
rect 1692 1868 1708 1932
rect 1772 1868 1788 1932
rect 1852 1868 1868 1932
rect 1932 1868 1940 1932
rect 1140 1852 1940 1868
rect 1140 1788 1148 1852
rect 1212 1788 1228 1852
rect 1292 1788 1308 1852
rect 1372 1788 1388 1852
rect 1452 1788 1468 1852
rect 1532 1788 1548 1852
rect 1612 1788 1628 1852
rect 1692 1788 1708 1852
rect 1772 1788 1788 1852
rect 1852 1788 1868 1852
rect 1932 1788 1940 1852
rect 1140 1772 1940 1788
rect 1140 1708 1148 1772
rect 1212 1708 1228 1772
rect 1292 1708 1308 1772
rect 1372 1708 1388 1772
rect 1452 1708 1468 1772
rect 1532 1708 1548 1772
rect 1612 1708 1628 1772
rect 1692 1708 1708 1772
rect 1772 1708 1788 1772
rect 1852 1708 1868 1772
rect 1932 1708 1940 1772
rect 1140 1692 1940 1708
rect 1140 1628 1148 1692
rect 1212 1628 1228 1692
rect 1292 1628 1308 1692
rect 1372 1628 1388 1692
rect 1452 1628 1468 1692
rect 1532 1628 1548 1692
rect 1612 1628 1628 1692
rect 1692 1628 1708 1692
rect 1772 1628 1788 1692
rect 1852 1628 1868 1692
rect 1932 1628 1940 1692
rect 1140 1612 1940 1628
rect 1140 1548 1148 1612
rect 1212 1548 1228 1612
rect 1292 1548 1308 1612
rect 1372 1548 1388 1612
rect 1452 1548 1468 1612
rect 1532 1548 1548 1612
rect 1612 1548 1628 1612
rect 1692 1548 1708 1612
rect 1772 1548 1788 1612
rect 1852 1548 1868 1612
rect 1932 1548 1940 1612
rect 1140 1532 1940 1548
rect 1140 1468 1148 1532
rect 1212 1468 1228 1532
rect 1292 1468 1308 1532
rect 1372 1468 1388 1532
rect 1452 1468 1468 1532
rect 1532 1468 1548 1532
rect 1612 1468 1628 1532
rect 1692 1468 1708 1532
rect 1772 1468 1788 1532
rect 1852 1468 1868 1532
rect 1932 1468 1940 1532
rect 1140 1452 1940 1468
rect 1140 1388 1148 1452
rect 1212 1388 1228 1452
rect 1292 1388 1308 1452
rect 1372 1388 1388 1452
rect 1452 1388 1468 1452
rect 1532 1388 1548 1452
rect 1612 1388 1628 1452
rect 1692 1388 1708 1452
rect 1772 1388 1788 1452
rect 1852 1388 1868 1452
rect 1932 1388 1940 1452
rect 1140 1372 1940 1388
rect 1140 1308 1148 1372
rect 1212 1308 1228 1372
rect 1292 1308 1308 1372
rect 1372 1308 1388 1372
rect 1452 1308 1468 1372
rect 1532 1308 1548 1372
rect 1612 1308 1628 1372
rect 1692 1308 1708 1372
rect 1772 1308 1788 1372
rect 1852 1308 1868 1372
rect 1932 1308 1940 1372
rect 1140 1292 1940 1308
rect 1140 1228 1148 1292
rect 1212 1228 1228 1292
rect 1292 1228 1308 1292
rect 1372 1228 1388 1292
rect 1452 1228 1468 1292
rect 1532 1228 1548 1292
rect 1612 1228 1628 1292
rect 1692 1228 1708 1292
rect 1772 1228 1788 1292
rect 1852 1228 1868 1292
rect 1932 1228 1940 1292
rect 1140 1212 1940 1228
rect 1140 1148 1148 1212
rect 1212 1148 1228 1212
rect 1292 1148 1308 1212
rect 1372 1148 1388 1212
rect 1452 1148 1468 1212
rect 1532 1148 1548 1212
rect 1612 1148 1628 1212
rect 1692 1148 1708 1212
rect 1772 1148 1788 1212
rect 1852 1148 1868 1212
rect 1932 1148 1940 1212
rect 1140 1140 1940 1148
rect 3995 8596 4415 9744
rect 3995 8532 4013 8596
rect 4077 8532 4093 8596
rect 4157 8532 4173 8596
rect 4237 8532 4253 8596
rect 4317 8532 4333 8596
rect 4397 8532 4415 8596
rect 3995 8516 4415 8532
rect 3995 8452 4013 8516
rect 4077 8452 4093 8516
rect 4157 8452 4173 8516
rect 4237 8452 4253 8516
rect 4317 8452 4333 8516
rect 4397 8452 4415 8516
rect 3995 8436 4415 8452
rect 3995 8372 4013 8436
rect 4077 8372 4093 8436
rect 4157 8372 4173 8436
rect 4237 8372 4253 8436
rect 4317 8372 4333 8436
rect 4397 8372 4415 8436
rect 3995 8356 4415 8372
rect 3995 8292 4013 8356
rect 4077 8292 4093 8356
rect 4157 8292 4173 8356
rect 4237 8292 4253 8356
rect 4317 8292 4333 8356
rect 4397 8292 4415 8356
rect 3995 8276 4415 8292
rect 3995 8212 4013 8276
rect 4077 8212 4093 8276
rect 4157 8212 4173 8276
rect 4237 8212 4253 8276
rect 4317 8212 4333 8276
rect 4397 8212 4415 8276
rect 3995 8196 4415 8212
rect 3995 8132 4013 8196
rect 4077 8132 4093 8196
rect 4157 8132 4173 8196
rect 4237 8132 4253 8196
rect 4317 8132 4333 8196
rect 4397 8132 4415 8196
rect 3995 8116 4415 8132
rect 3995 8052 4013 8116
rect 4077 8052 4093 8116
rect 4157 8052 4173 8116
rect 4237 8052 4253 8116
rect 4317 8052 4333 8116
rect 4397 8052 4415 8116
rect 3995 8036 4415 8052
rect 3995 7972 4013 8036
rect 4077 7972 4093 8036
rect 4157 7972 4173 8036
rect 4237 7972 4253 8036
rect 4317 7972 4333 8036
rect 4397 7972 4415 8036
rect 3995 7956 4415 7972
rect 3995 7892 4013 7956
rect 4077 7892 4093 7956
rect 4157 7892 4173 7956
rect 4237 7892 4253 7956
rect 4317 7892 4333 7956
rect 4397 7892 4415 7956
rect 3995 7876 4415 7892
rect 3995 7812 4013 7876
rect 4077 7812 4093 7876
rect 4157 7812 4173 7876
rect 4237 7812 4253 7876
rect 4317 7812 4333 7876
rect 4397 7812 4415 7876
rect 3995 6536 4415 7812
rect 3995 6472 4013 6536
rect 4077 6472 4093 6536
rect 4157 6472 4173 6536
rect 4237 6472 4253 6536
rect 4317 6472 4333 6536
rect 4397 6472 4415 6536
rect 3995 5448 4415 6472
rect 3995 5384 4013 5448
rect 4077 5384 4093 5448
rect 4157 5384 4173 5448
rect 4237 5384 4253 5448
rect 4317 5384 4333 5448
rect 4397 5384 4415 5448
rect 3995 4360 4415 5384
rect 3995 4296 4013 4360
rect 4077 4296 4093 4360
rect 4157 4296 4173 4360
rect 4237 4296 4253 4360
rect 4317 4296 4333 4360
rect 4397 4296 4415 4360
rect 3995 3272 4415 4296
rect 3995 3208 4013 3272
rect 4077 3208 4093 3272
rect 4157 3208 4173 3272
rect 4237 3208 4253 3272
rect 4317 3208 4333 3272
rect 4397 3208 4415 3272
rect 3995 1932 4415 3208
rect 3995 1868 4013 1932
rect 4077 1868 4093 1932
rect 4157 1868 4173 1932
rect 4237 1868 4253 1932
rect 4317 1868 4333 1932
rect 4397 1868 4415 1932
rect 3995 1852 4415 1868
rect 3995 1788 4013 1852
rect 4077 1788 4093 1852
rect 4157 1788 4173 1852
rect 4237 1788 4253 1852
rect 4317 1788 4333 1852
rect 4397 1788 4415 1852
rect 3995 1772 4415 1788
rect 3995 1708 4013 1772
rect 4077 1708 4093 1772
rect 4157 1708 4173 1772
rect 4237 1708 4253 1772
rect 4317 1708 4333 1772
rect 4397 1708 4415 1772
rect 3995 1692 4415 1708
rect 3995 1628 4013 1692
rect 4077 1628 4093 1692
rect 4157 1628 4173 1692
rect 4237 1628 4253 1692
rect 4317 1628 4333 1692
rect 4397 1628 4415 1692
rect 3995 1612 4415 1628
rect 3995 1548 4013 1612
rect 4077 1548 4093 1612
rect 4157 1548 4173 1612
rect 4237 1548 4253 1612
rect 4317 1548 4333 1612
rect 4397 1548 4415 1612
rect 3995 1532 4415 1548
rect 3995 1468 4013 1532
rect 4077 1468 4093 1532
rect 4157 1468 4173 1532
rect 4237 1468 4253 1532
rect 4317 1468 4333 1532
rect 4397 1468 4415 1532
rect 3995 1452 4415 1468
rect 3995 1388 4013 1452
rect 4077 1388 4093 1452
rect 4157 1388 4173 1452
rect 4237 1388 4253 1452
rect 4317 1388 4333 1452
rect 4397 1388 4415 1452
rect 3995 1372 4415 1388
rect 3995 1308 4013 1372
rect 4077 1308 4093 1372
rect 4157 1308 4173 1372
rect 4237 1308 4253 1372
rect 4317 1308 4333 1372
rect 4397 1308 4415 1372
rect 3995 1292 4415 1308
rect 3995 1228 4013 1292
rect 4077 1228 4093 1292
rect 4157 1228 4173 1292
rect 4237 1228 4253 1292
rect 4317 1228 4333 1292
rect 4397 1228 4415 1292
rect 3995 1212 4415 1228
rect 3995 1148 4013 1212
rect 4077 1148 4093 1212
rect 4157 1148 4173 1212
rect 4237 1148 4253 1212
rect 4317 1148 4333 1212
rect 4397 1148 4415 1212
rect 0 728 8 792
rect 72 728 88 792
rect 152 728 168 792
rect 232 728 248 792
rect 312 728 328 792
rect 392 728 408 792
rect 472 728 488 792
rect 552 728 568 792
rect 632 728 648 792
rect 712 728 728 792
rect 792 728 800 792
rect 0 712 800 728
rect 0 648 8 712
rect 72 648 88 712
rect 152 648 168 712
rect 232 648 248 712
rect 312 648 328 712
rect 392 648 408 712
rect 472 648 488 712
rect 552 648 568 712
rect 632 648 648 712
rect 712 648 728 712
rect 792 648 800 712
rect 0 632 800 648
rect 0 568 8 632
rect 72 568 88 632
rect 152 568 168 632
rect 232 568 248 632
rect 312 568 328 632
rect 392 568 408 632
rect 472 568 488 632
rect 552 568 568 632
rect 632 568 648 632
rect 712 568 728 632
rect 792 568 800 632
rect 0 552 800 568
rect 0 488 8 552
rect 72 488 88 552
rect 152 488 168 552
rect 232 488 248 552
rect 312 488 328 552
rect 392 488 408 552
rect 472 488 488 552
rect 552 488 568 552
rect 632 488 648 552
rect 712 488 728 552
rect 792 488 800 552
rect 0 472 800 488
rect 0 408 8 472
rect 72 408 88 472
rect 152 408 168 472
rect 232 408 248 472
rect 312 408 328 472
rect 392 408 408 472
rect 472 408 488 472
rect 552 408 568 472
rect 632 408 648 472
rect 712 408 728 472
rect 792 408 800 472
rect 0 392 800 408
rect 0 328 8 392
rect 72 328 88 392
rect 152 328 168 392
rect 232 328 248 392
rect 312 328 328 392
rect 392 328 408 392
rect 472 328 488 392
rect 552 328 568 392
rect 632 328 648 392
rect 712 328 728 392
rect 792 328 800 392
rect 0 312 800 328
rect 0 248 8 312
rect 72 248 88 312
rect 152 248 168 312
rect 232 248 248 312
rect 312 248 328 312
rect 392 248 408 312
rect 472 248 488 312
rect 552 248 568 312
rect 632 248 648 312
rect 712 248 728 312
rect 792 248 800 312
rect 0 232 800 248
rect 0 168 8 232
rect 72 168 88 232
rect 152 168 168 232
rect 232 168 248 232
rect 312 168 328 232
rect 392 168 408 232
rect 472 168 488 232
rect 552 168 568 232
rect 632 168 648 232
rect 712 168 728 232
rect 792 168 800 232
rect 0 152 800 168
rect 0 88 8 152
rect 72 88 88 152
rect 152 88 168 152
rect 232 88 248 152
rect 312 88 328 152
rect 392 88 408 152
rect 472 88 488 152
rect 552 88 568 152
rect 632 88 648 152
rect 712 88 728 152
rect 792 88 800 152
rect 0 72 800 88
rect 0 8 8 72
rect 72 8 88 72
rect 152 8 168 72
rect 232 8 248 72
rect 312 8 328 72
rect 392 8 408 72
rect 472 8 488 72
rect 552 8 568 72
rect 632 8 648 72
rect 712 8 728 72
rect 792 8 800 72
rect 0 0 800 8
rect 3995 0 4415 1148
rect 4960 9736 5381 9744
rect 4960 9672 4978 9736
rect 5042 9672 5058 9736
rect 5122 9672 5138 9736
rect 5202 9672 5218 9736
rect 5282 9672 5298 9736
rect 5362 9672 5381 9736
rect 4960 9656 5381 9672
rect 4960 9592 4978 9656
rect 5042 9592 5058 9656
rect 5122 9592 5138 9656
rect 5202 9592 5218 9656
rect 5282 9592 5298 9656
rect 5362 9592 5381 9656
rect 4960 9576 5381 9592
rect 4960 9512 4978 9576
rect 5042 9512 5058 9576
rect 5122 9512 5138 9576
rect 5202 9512 5218 9576
rect 5282 9512 5298 9576
rect 5362 9512 5381 9576
rect 4960 9496 5381 9512
rect 4960 9432 4978 9496
rect 5042 9432 5058 9496
rect 5122 9432 5138 9496
rect 5202 9432 5218 9496
rect 5282 9432 5298 9496
rect 5362 9432 5381 9496
rect 4960 9416 5381 9432
rect 4960 9352 4978 9416
rect 5042 9352 5058 9416
rect 5122 9352 5138 9416
rect 5202 9352 5218 9416
rect 5282 9352 5298 9416
rect 5362 9352 5381 9416
rect 4960 9336 5381 9352
rect 4960 9272 4978 9336
rect 5042 9272 5058 9336
rect 5122 9272 5138 9336
rect 5202 9272 5218 9336
rect 5282 9272 5298 9336
rect 5362 9272 5381 9336
rect 4960 9256 5381 9272
rect 4960 9192 4978 9256
rect 5042 9192 5058 9256
rect 5122 9192 5138 9256
rect 5202 9192 5218 9256
rect 5282 9192 5298 9256
rect 5362 9192 5381 9256
rect 4960 9176 5381 9192
rect 4960 9112 4978 9176
rect 5042 9112 5058 9176
rect 5122 9112 5138 9176
rect 5202 9112 5218 9176
rect 5282 9112 5298 9176
rect 5362 9112 5381 9176
rect 4960 9096 5381 9112
rect 4960 9032 4978 9096
rect 5042 9032 5058 9096
rect 5122 9032 5138 9096
rect 5202 9032 5218 9096
rect 5282 9032 5298 9096
rect 5362 9032 5381 9096
rect 4960 9016 5381 9032
rect 4960 8952 4978 9016
rect 5042 8952 5058 9016
rect 5122 8952 5138 9016
rect 5202 8952 5218 9016
rect 5282 8952 5298 9016
rect 5362 8952 5381 9016
rect 4960 5992 5381 8952
rect 4960 5928 4978 5992
rect 5042 5928 5058 5992
rect 5122 5928 5138 5992
rect 5202 5928 5218 5992
rect 5282 5928 5298 5992
rect 5362 5928 5381 5992
rect 4960 4904 5381 5928
rect 4960 4840 4978 4904
rect 5042 4840 5058 4904
rect 5122 4840 5138 4904
rect 5202 4840 5218 4904
rect 5282 4840 5298 4904
rect 5362 4840 5381 4904
rect 4960 3816 5381 4840
rect 4960 3752 4978 3816
rect 5042 3752 5058 3816
rect 5122 3752 5138 3816
rect 5202 3752 5218 3816
rect 5282 3752 5298 3816
rect 5362 3752 5381 3816
rect 4960 792 5381 3752
rect 4960 728 4978 792
rect 5042 728 5058 792
rect 5122 728 5138 792
rect 5202 728 5218 792
rect 5282 728 5298 792
rect 5362 728 5381 792
rect 4960 712 5381 728
rect 4960 648 4978 712
rect 5042 648 5058 712
rect 5122 648 5138 712
rect 5202 648 5218 712
rect 5282 648 5298 712
rect 5362 648 5381 712
rect 4960 632 5381 648
rect 4960 568 4978 632
rect 5042 568 5058 632
rect 5122 568 5138 632
rect 5202 568 5218 632
rect 5282 568 5298 632
rect 5362 568 5381 632
rect 4960 552 5381 568
rect 4960 488 4978 552
rect 5042 488 5058 552
rect 5122 488 5138 552
rect 5202 488 5218 552
rect 5282 488 5298 552
rect 5362 488 5381 552
rect 4960 472 5381 488
rect 4960 408 4978 472
rect 5042 408 5058 472
rect 5122 408 5138 472
rect 5202 408 5218 472
rect 5282 408 5298 472
rect 5362 408 5381 472
rect 4960 392 5381 408
rect 4960 328 4978 392
rect 5042 328 5058 392
rect 5122 328 5138 392
rect 5202 328 5218 392
rect 5282 328 5298 392
rect 5362 328 5381 392
rect 4960 312 5381 328
rect 4960 248 4978 312
rect 5042 248 5058 312
rect 5122 248 5138 312
rect 5202 248 5218 312
rect 5282 248 5298 312
rect 5362 248 5381 312
rect 4960 232 5381 248
rect 4960 168 4978 232
rect 5042 168 5058 232
rect 5122 168 5138 232
rect 5202 168 5218 232
rect 5282 168 5298 232
rect 5362 168 5381 232
rect 4960 152 5381 168
rect 4960 88 4978 152
rect 5042 88 5058 152
rect 5122 88 5138 152
rect 5202 88 5218 152
rect 5282 88 5298 152
rect 5362 88 5381 152
rect 4960 72 5381 88
rect 4960 8 4978 72
rect 5042 8 5058 72
rect 5122 8 5138 72
rect 5202 8 5218 72
rect 5282 8 5298 72
rect 5362 8 5381 72
rect 4960 0 5381 8
rect 5926 8596 6346 9744
rect 5926 8532 5944 8596
rect 6008 8532 6024 8596
rect 6088 8532 6104 8596
rect 6168 8532 6184 8596
rect 6248 8532 6264 8596
rect 6328 8532 6346 8596
rect 5926 8516 6346 8532
rect 5926 8452 5944 8516
rect 6008 8452 6024 8516
rect 6088 8452 6104 8516
rect 6168 8452 6184 8516
rect 6248 8452 6264 8516
rect 6328 8452 6346 8516
rect 5926 8436 6346 8452
rect 5926 8372 5944 8436
rect 6008 8372 6024 8436
rect 6088 8372 6104 8436
rect 6168 8372 6184 8436
rect 6248 8372 6264 8436
rect 6328 8372 6346 8436
rect 5926 8356 6346 8372
rect 5926 8292 5944 8356
rect 6008 8292 6024 8356
rect 6088 8292 6104 8356
rect 6168 8292 6184 8356
rect 6248 8292 6264 8356
rect 6328 8292 6346 8356
rect 5926 8276 6346 8292
rect 5926 8212 5944 8276
rect 6008 8212 6024 8276
rect 6088 8212 6104 8276
rect 6168 8212 6184 8276
rect 6248 8212 6264 8276
rect 6328 8212 6346 8276
rect 5926 8196 6346 8212
rect 5926 8132 5944 8196
rect 6008 8132 6024 8196
rect 6088 8132 6104 8196
rect 6168 8132 6184 8196
rect 6248 8132 6264 8196
rect 6328 8132 6346 8196
rect 5926 8116 6346 8132
rect 5926 8052 5944 8116
rect 6008 8052 6024 8116
rect 6088 8052 6104 8116
rect 6168 8052 6184 8116
rect 6248 8052 6264 8116
rect 6328 8052 6346 8116
rect 5926 8036 6346 8052
rect 5926 7972 5944 8036
rect 6008 7972 6024 8036
rect 6088 7972 6104 8036
rect 6168 7972 6184 8036
rect 6248 7972 6264 8036
rect 6328 7972 6346 8036
rect 5926 7956 6346 7972
rect 5926 7892 5944 7956
rect 6008 7892 6024 7956
rect 6088 7892 6104 7956
rect 6168 7892 6184 7956
rect 6248 7892 6264 7956
rect 6328 7892 6346 7956
rect 5926 7876 6346 7892
rect 5926 7812 5944 7876
rect 6008 7812 6024 7876
rect 6088 7812 6104 7876
rect 6168 7812 6184 7876
rect 6248 7812 6264 7876
rect 6328 7812 6346 7876
rect 5926 6536 6346 7812
rect 5926 6472 5944 6536
rect 6008 6472 6024 6536
rect 6088 6472 6104 6536
rect 6168 6472 6184 6536
rect 6248 6472 6264 6536
rect 6328 6472 6346 6536
rect 5926 5448 6346 6472
rect 5926 5384 5944 5448
rect 6008 5384 6024 5448
rect 6088 5384 6104 5448
rect 6168 5384 6184 5448
rect 6248 5384 6264 5448
rect 6328 5384 6346 5448
rect 5926 4360 6346 5384
rect 5926 4296 5944 4360
rect 6008 4296 6024 4360
rect 6088 4296 6104 4360
rect 6168 4296 6184 4360
rect 6248 4296 6264 4360
rect 6328 4296 6346 4360
rect 5926 3272 6346 4296
rect 5926 3208 5944 3272
rect 6008 3208 6024 3272
rect 6088 3208 6104 3272
rect 6168 3208 6184 3272
rect 6248 3208 6264 3272
rect 6328 3208 6346 3272
rect 5926 1932 6346 3208
rect 5926 1868 5944 1932
rect 6008 1868 6024 1932
rect 6088 1868 6104 1932
rect 6168 1868 6184 1932
rect 6248 1868 6264 1932
rect 6328 1868 6346 1932
rect 5926 1852 6346 1868
rect 5926 1788 5944 1852
rect 6008 1788 6024 1852
rect 6088 1788 6104 1852
rect 6168 1788 6184 1852
rect 6248 1788 6264 1852
rect 6328 1788 6346 1852
rect 5926 1772 6346 1788
rect 5926 1708 5944 1772
rect 6008 1708 6024 1772
rect 6088 1708 6104 1772
rect 6168 1708 6184 1772
rect 6248 1708 6264 1772
rect 6328 1708 6346 1772
rect 5926 1692 6346 1708
rect 5926 1628 5944 1692
rect 6008 1628 6024 1692
rect 6088 1628 6104 1692
rect 6168 1628 6184 1692
rect 6248 1628 6264 1692
rect 6328 1628 6346 1692
rect 5926 1612 6346 1628
rect 5926 1548 5944 1612
rect 6008 1548 6024 1612
rect 6088 1548 6104 1612
rect 6168 1548 6184 1612
rect 6248 1548 6264 1612
rect 6328 1548 6346 1612
rect 5926 1532 6346 1548
rect 5926 1468 5944 1532
rect 6008 1468 6024 1532
rect 6088 1468 6104 1532
rect 6168 1468 6184 1532
rect 6248 1468 6264 1532
rect 6328 1468 6346 1532
rect 5926 1452 6346 1468
rect 5926 1388 5944 1452
rect 6008 1388 6024 1452
rect 6088 1388 6104 1452
rect 6168 1388 6184 1452
rect 6248 1388 6264 1452
rect 6328 1388 6346 1452
rect 5926 1372 6346 1388
rect 5926 1308 5944 1372
rect 6008 1308 6024 1372
rect 6088 1308 6104 1372
rect 6168 1308 6184 1372
rect 6248 1308 6264 1372
rect 6328 1308 6346 1372
rect 5926 1292 6346 1308
rect 5926 1228 5944 1292
rect 6008 1228 6024 1292
rect 6088 1228 6104 1292
rect 6168 1228 6184 1292
rect 6248 1228 6264 1292
rect 6328 1228 6346 1292
rect 5926 1212 6346 1228
rect 5926 1148 5944 1212
rect 6008 1148 6024 1212
rect 6088 1148 6104 1212
rect 6168 1148 6184 1212
rect 6248 1148 6264 1212
rect 6328 1148 6346 1212
rect 5926 0 6346 1148
rect 6891 9736 7311 9744
rect 6891 9672 6909 9736
rect 6973 9672 6989 9736
rect 7053 9672 7069 9736
rect 7133 9672 7149 9736
rect 7213 9672 7229 9736
rect 7293 9672 7311 9736
rect 6891 9656 7311 9672
rect 6891 9592 6909 9656
rect 6973 9592 6989 9656
rect 7053 9592 7069 9656
rect 7133 9592 7149 9656
rect 7213 9592 7229 9656
rect 7293 9592 7311 9656
rect 6891 9576 7311 9592
rect 6891 9512 6909 9576
rect 6973 9512 6989 9576
rect 7053 9512 7069 9576
rect 7133 9512 7149 9576
rect 7213 9512 7229 9576
rect 7293 9512 7311 9576
rect 6891 9496 7311 9512
rect 6891 9432 6909 9496
rect 6973 9432 6989 9496
rect 7053 9432 7069 9496
rect 7133 9432 7149 9496
rect 7213 9432 7229 9496
rect 7293 9432 7311 9496
rect 6891 9416 7311 9432
rect 6891 9352 6909 9416
rect 6973 9352 6989 9416
rect 7053 9352 7069 9416
rect 7133 9352 7149 9416
rect 7213 9352 7229 9416
rect 7293 9352 7311 9416
rect 6891 9336 7311 9352
rect 6891 9272 6909 9336
rect 6973 9272 6989 9336
rect 7053 9272 7069 9336
rect 7133 9272 7149 9336
rect 7213 9272 7229 9336
rect 7293 9272 7311 9336
rect 6891 9256 7311 9272
rect 6891 9192 6909 9256
rect 6973 9192 6989 9256
rect 7053 9192 7069 9256
rect 7133 9192 7149 9256
rect 7213 9192 7229 9256
rect 7293 9192 7311 9256
rect 6891 9176 7311 9192
rect 6891 9112 6909 9176
rect 6973 9112 6989 9176
rect 7053 9112 7069 9176
rect 7133 9112 7149 9176
rect 7213 9112 7229 9176
rect 7293 9112 7311 9176
rect 6891 9096 7311 9112
rect 6891 9032 6909 9096
rect 6973 9032 6989 9096
rect 7053 9032 7069 9096
rect 7133 9032 7149 9096
rect 7213 9032 7229 9096
rect 7293 9032 7311 9096
rect 6891 9016 7311 9032
rect 6891 8952 6909 9016
rect 6973 8952 6989 9016
rect 7053 8952 7069 9016
rect 7133 8952 7149 9016
rect 7213 8952 7229 9016
rect 7293 8952 7311 9016
rect 6891 5992 7311 8952
rect 6891 5928 6909 5992
rect 6973 5928 6989 5992
rect 7053 5928 7069 5992
rect 7133 5928 7149 5992
rect 7213 5928 7229 5992
rect 7293 5928 7311 5992
rect 6891 4904 7311 5928
rect 6891 4840 6909 4904
rect 6973 4840 6989 4904
rect 7053 4840 7069 4904
rect 7133 4840 7149 4904
rect 7213 4840 7229 4904
rect 7293 4840 7311 4904
rect 6891 3816 7311 4840
rect 6891 3752 6909 3816
rect 6973 3752 6989 3816
rect 7053 3752 7069 3816
rect 7133 3752 7149 3816
rect 7213 3752 7229 3816
rect 7293 3752 7311 3816
rect 6891 792 7311 3752
rect 6891 728 6909 792
rect 6973 728 6989 792
rect 7053 728 7069 792
rect 7133 728 7149 792
rect 7213 728 7229 792
rect 7293 728 7311 792
rect 6891 712 7311 728
rect 6891 648 6909 712
rect 6973 648 6989 712
rect 7053 648 7069 712
rect 7133 648 7149 712
rect 7213 648 7229 712
rect 7293 648 7311 712
rect 6891 632 7311 648
rect 6891 568 6909 632
rect 6973 568 6989 632
rect 7053 568 7069 632
rect 7133 568 7149 632
rect 7213 568 7229 632
rect 7293 568 7311 632
rect 6891 552 7311 568
rect 6891 488 6909 552
rect 6973 488 6989 552
rect 7053 488 7069 552
rect 7133 488 7149 552
rect 7213 488 7229 552
rect 7293 488 7311 552
rect 6891 472 7311 488
rect 6891 408 6909 472
rect 6973 408 6989 472
rect 7053 408 7069 472
rect 7133 408 7149 472
rect 7213 408 7229 472
rect 7293 408 7311 472
rect 6891 392 7311 408
rect 6891 328 6909 392
rect 6973 328 6989 392
rect 7053 328 7069 392
rect 7133 328 7149 392
rect 7213 328 7229 392
rect 7293 328 7311 392
rect 6891 312 7311 328
rect 6891 248 6909 312
rect 6973 248 6989 312
rect 7053 248 7069 312
rect 7133 248 7149 312
rect 7213 248 7229 312
rect 7293 248 7311 312
rect 6891 232 7311 248
rect 6891 168 6909 232
rect 6973 168 6989 232
rect 7053 168 7069 232
rect 7133 168 7149 232
rect 7213 168 7229 232
rect 7293 168 7311 232
rect 6891 152 7311 168
rect 6891 88 6909 152
rect 6973 88 6989 152
rect 7053 88 7069 152
rect 7133 88 7149 152
rect 7213 88 7229 152
rect 7293 88 7311 152
rect 6891 72 7311 88
rect 6891 8 6909 72
rect 6973 8 6989 72
rect 7053 8 7069 72
rect 7133 8 7149 72
rect 7213 8 7229 72
rect 7293 8 7311 72
rect 6891 0 7311 8
rect 7856 8596 8277 9744
rect 11384 9736 12184 9744
rect 11384 9672 11392 9736
rect 11456 9672 11472 9736
rect 11536 9672 11552 9736
rect 11616 9672 11632 9736
rect 11696 9672 11712 9736
rect 11776 9672 11792 9736
rect 11856 9672 11872 9736
rect 11936 9672 11952 9736
rect 12016 9672 12032 9736
rect 12096 9672 12112 9736
rect 12176 9672 12184 9736
rect 11384 9656 12184 9672
rect 11384 9592 11392 9656
rect 11456 9592 11472 9656
rect 11536 9592 11552 9656
rect 11616 9592 11632 9656
rect 11696 9592 11712 9656
rect 11776 9592 11792 9656
rect 11856 9592 11872 9656
rect 11936 9592 11952 9656
rect 12016 9592 12032 9656
rect 12096 9592 12112 9656
rect 12176 9592 12184 9656
rect 11384 9576 12184 9592
rect 11384 9512 11392 9576
rect 11456 9512 11472 9576
rect 11536 9512 11552 9576
rect 11616 9512 11632 9576
rect 11696 9512 11712 9576
rect 11776 9512 11792 9576
rect 11856 9512 11872 9576
rect 11936 9512 11952 9576
rect 12016 9512 12032 9576
rect 12096 9512 12112 9576
rect 12176 9512 12184 9576
rect 11384 9496 12184 9512
rect 11384 9432 11392 9496
rect 11456 9432 11472 9496
rect 11536 9432 11552 9496
rect 11616 9432 11632 9496
rect 11696 9432 11712 9496
rect 11776 9432 11792 9496
rect 11856 9432 11872 9496
rect 11936 9432 11952 9496
rect 12016 9432 12032 9496
rect 12096 9432 12112 9496
rect 12176 9432 12184 9496
rect 11384 9416 12184 9432
rect 11384 9352 11392 9416
rect 11456 9352 11472 9416
rect 11536 9352 11552 9416
rect 11616 9352 11632 9416
rect 11696 9352 11712 9416
rect 11776 9352 11792 9416
rect 11856 9352 11872 9416
rect 11936 9352 11952 9416
rect 12016 9352 12032 9416
rect 12096 9352 12112 9416
rect 12176 9352 12184 9416
rect 11384 9336 12184 9352
rect 11384 9272 11392 9336
rect 11456 9272 11472 9336
rect 11536 9272 11552 9336
rect 11616 9272 11632 9336
rect 11696 9272 11712 9336
rect 11776 9272 11792 9336
rect 11856 9272 11872 9336
rect 11936 9272 11952 9336
rect 12016 9272 12032 9336
rect 12096 9272 12112 9336
rect 12176 9272 12184 9336
rect 11384 9256 12184 9272
rect 11384 9192 11392 9256
rect 11456 9192 11472 9256
rect 11536 9192 11552 9256
rect 11616 9192 11632 9256
rect 11696 9192 11712 9256
rect 11776 9192 11792 9256
rect 11856 9192 11872 9256
rect 11936 9192 11952 9256
rect 12016 9192 12032 9256
rect 12096 9192 12112 9256
rect 12176 9192 12184 9256
rect 11384 9176 12184 9192
rect 11384 9112 11392 9176
rect 11456 9112 11472 9176
rect 11536 9112 11552 9176
rect 11616 9112 11632 9176
rect 11696 9112 11712 9176
rect 11776 9112 11792 9176
rect 11856 9112 11872 9176
rect 11936 9112 11952 9176
rect 12016 9112 12032 9176
rect 12096 9112 12112 9176
rect 12176 9112 12184 9176
rect 11384 9096 12184 9112
rect 11384 9032 11392 9096
rect 11456 9032 11472 9096
rect 11536 9032 11552 9096
rect 11616 9032 11632 9096
rect 11696 9032 11712 9096
rect 11776 9032 11792 9096
rect 11856 9032 11872 9096
rect 11936 9032 11952 9096
rect 12016 9032 12032 9096
rect 12096 9032 12112 9096
rect 12176 9032 12184 9096
rect 11384 9016 12184 9032
rect 11384 8952 11392 9016
rect 11456 8952 11472 9016
rect 11536 8952 11552 9016
rect 11616 8952 11632 9016
rect 11696 8952 11712 9016
rect 11776 8952 11792 9016
rect 11856 8952 11872 9016
rect 11936 8952 11952 9016
rect 12016 8952 12032 9016
rect 12096 8952 12112 9016
rect 12176 8952 12184 9016
rect 7856 8532 7874 8596
rect 7938 8532 7954 8596
rect 8018 8532 8034 8596
rect 8098 8532 8114 8596
rect 8178 8532 8194 8596
rect 8258 8532 8277 8596
rect 7856 8516 8277 8532
rect 7856 8452 7874 8516
rect 7938 8452 7954 8516
rect 8018 8452 8034 8516
rect 8098 8452 8114 8516
rect 8178 8452 8194 8516
rect 8258 8452 8277 8516
rect 7856 8436 8277 8452
rect 7856 8372 7874 8436
rect 7938 8372 7954 8436
rect 8018 8372 8034 8436
rect 8098 8372 8114 8436
rect 8178 8372 8194 8436
rect 8258 8372 8277 8436
rect 7856 8356 8277 8372
rect 7856 8292 7874 8356
rect 7938 8292 7954 8356
rect 8018 8292 8034 8356
rect 8098 8292 8114 8356
rect 8178 8292 8194 8356
rect 8258 8292 8277 8356
rect 7856 8276 8277 8292
rect 7856 8212 7874 8276
rect 7938 8212 7954 8276
rect 8018 8212 8034 8276
rect 8098 8212 8114 8276
rect 8178 8212 8194 8276
rect 8258 8212 8277 8276
rect 7856 8196 8277 8212
rect 7856 8132 7874 8196
rect 7938 8132 7954 8196
rect 8018 8132 8034 8196
rect 8098 8132 8114 8196
rect 8178 8132 8194 8196
rect 8258 8132 8277 8196
rect 7856 8116 8277 8132
rect 7856 8052 7874 8116
rect 7938 8052 7954 8116
rect 8018 8052 8034 8116
rect 8098 8052 8114 8116
rect 8178 8052 8194 8116
rect 8258 8052 8277 8116
rect 7856 8036 8277 8052
rect 7856 7972 7874 8036
rect 7938 7972 7954 8036
rect 8018 7972 8034 8036
rect 8098 7972 8114 8036
rect 8178 7972 8194 8036
rect 8258 7972 8277 8036
rect 7856 7956 8277 7972
rect 7856 7892 7874 7956
rect 7938 7892 7954 7956
rect 8018 7892 8034 7956
rect 8098 7892 8114 7956
rect 8178 7892 8194 7956
rect 8258 7892 8277 7956
rect 7856 7876 8277 7892
rect 7856 7812 7874 7876
rect 7938 7812 7954 7876
rect 8018 7812 8034 7876
rect 8098 7812 8114 7876
rect 8178 7812 8194 7876
rect 8258 7812 8277 7876
rect 7856 6536 8277 7812
rect 7856 6472 7874 6536
rect 7938 6472 7954 6536
rect 8018 6472 8034 6536
rect 8098 6472 8114 6536
rect 8178 6472 8194 6536
rect 8258 6472 8277 6536
rect 7856 5448 8277 6472
rect 7856 5384 7874 5448
rect 7938 5384 7954 5448
rect 8018 5384 8034 5448
rect 8098 5384 8114 5448
rect 8178 5384 8194 5448
rect 8258 5384 8277 5448
rect 7856 4360 8277 5384
rect 7856 4296 7874 4360
rect 7938 4296 7954 4360
rect 8018 4296 8034 4360
rect 8098 4296 8114 4360
rect 8178 4296 8194 4360
rect 8258 4296 8277 4360
rect 7856 3272 8277 4296
rect 7856 3208 7874 3272
rect 7938 3208 7954 3272
rect 8018 3208 8034 3272
rect 8098 3208 8114 3272
rect 8178 3208 8194 3272
rect 8258 3208 8277 3272
rect 7856 1932 8277 3208
rect 7856 1868 7874 1932
rect 7938 1868 7954 1932
rect 8018 1868 8034 1932
rect 8098 1868 8114 1932
rect 8178 1868 8194 1932
rect 8258 1868 8277 1932
rect 7856 1852 8277 1868
rect 7856 1788 7874 1852
rect 7938 1788 7954 1852
rect 8018 1788 8034 1852
rect 8098 1788 8114 1852
rect 8178 1788 8194 1852
rect 8258 1788 8277 1852
rect 7856 1772 8277 1788
rect 7856 1708 7874 1772
rect 7938 1708 7954 1772
rect 8018 1708 8034 1772
rect 8098 1708 8114 1772
rect 8178 1708 8194 1772
rect 8258 1708 8277 1772
rect 7856 1692 8277 1708
rect 7856 1628 7874 1692
rect 7938 1628 7954 1692
rect 8018 1628 8034 1692
rect 8098 1628 8114 1692
rect 8178 1628 8194 1692
rect 8258 1628 8277 1692
rect 7856 1612 8277 1628
rect 7856 1548 7874 1612
rect 7938 1548 7954 1612
rect 8018 1548 8034 1612
rect 8098 1548 8114 1612
rect 8178 1548 8194 1612
rect 8258 1548 8277 1612
rect 7856 1532 8277 1548
rect 7856 1468 7874 1532
rect 7938 1468 7954 1532
rect 8018 1468 8034 1532
rect 8098 1468 8114 1532
rect 8178 1468 8194 1532
rect 8258 1468 8277 1532
rect 7856 1452 8277 1468
rect 7856 1388 7874 1452
rect 7938 1388 7954 1452
rect 8018 1388 8034 1452
rect 8098 1388 8114 1452
rect 8178 1388 8194 1452
rect 8258 1388 8277 1452
rect 7856 1372 8277 1388
rect 7856 1308 7874 1372
rect 7938 1308 7954 1372
rect 8018 1308 8034 1372
rect 8098 1308 8114 1372
rect 8178 1308 8194 1372
rect 8258 1308 8277 1372
rect 7856 1292 8277 1308
rect 7856 1228 7874 1292
rect 7938 1228 7954 1292
rect 8018 1228 8034 1292
rect 8098 1228 8114 1292
rect 8178 1228 8194 1292
rect 8258 1228 8277 1292
rect 7856 1212 8277 1228
rect 7856 1148 7874 1212
rect 7938 1148 7954 1212
rect 8018 1148 8034 1212
rect 8098 1148 8114 1212
rect 8178 1148 8194 1212
rect 8258 1148 8277 1212
rect 7856 0 8277 1148
rect 10244 8596 11044 8604
rect 10244 8532 10252 8596
rect 10316 8532 10332 8596
rect 10396 8532 10412 8596
rect 10476 8532 10492 8596
rect 10556 8532 10572 8596
rect 10636 8532 10652 8596
rect 10716 8532 10732 8596
rect 10796 8532 10812 8596
rect 10876 8532 10892 8596
rect 10956 8532 10972 8596
rect 11036 8532 11044 8596
rect 10244 8516 11044 8532
rect 10244 8452 10252 8516
rect 10316 8452 10332 8516
rect 10396 8452 10412 8516
rect 10476 8452 10492 8516
rect 10556 8452 10572 8516
rect 10636 8452 10652 8516
rect 10716 8452 10732 8516
rect 10796 8452 10812 8516
rect 10876 8452 10892 8516
rect 10956 8452 10972 8516
rect 11036 8452 11044 8516
rect 10244 8436 11044 8452
rect 10244 8372 10252 8436
rect 10316 8372 10332 8436
rect 10396 8372 10412 8436
rect 10476 8372 10492 8436
rect 10556 8372 10572 8436
rect 10636 8372 10652 8436
rect 10716 8372 10732 8436
rect 10796 8372 10812 8436
rect 10876 8372 10892 8436
rect 10956 8372 10972 8436
rect 11036 8372 11044 8436
rect 10244 8356 11044 8372
rect 10244 8292 10252 8356
rect 10316 8292 10332 8356
rect 10396 8292 10412 8356
rect 10476 8292 10492 8356
rect 10556 8292 10572 8356
rect 10636 8292 10652 8356
rect 10716 8292 10732 8356
rect 10796 8292 10812 8356
rect 10876 8292 10892 8356
rect 10956 8292 10972 8356
rect 11036 8292 11044 8356
rect 10244 8276 11044 8292
rect 10244 8212 10252 8276
rect 10316 8212 10332 8276
rect 10396 8212 10412 8276
rect 10476 8212 10492 8276
rect 10556 8212 10572 8276
rect 10636 8212 10652 8276
rect 10716 8212 10732 8276
rect 10796 8212 10812 8276
rect 10876 8212 10892 8276
rect 10956 8212 10972 8276
rect 11036 8212 11044 8276
rect 10244 8196 11044 8212
rect 10244 8132 10252 8196
rect 10316 8132 10332 8196
rect 10396 8132 10412 8196
rect 10476 8132 10492 8196
rect 10556 8132 10572 8196
rect 10636 8132 10652 8196
rect 10716 8132 10732 8196
rect 10796 8132 10812 8196
rect 10876 8132 10892 8196
rect 10956 8132 10972 8196
rect 11036 8132 11044 8196
rect 10244 8116 11044 8132
rect 10244 8052 10252 8116
rect 10316 8052 10332 8116
rect 10396 8052 10412 8116
rect 10476 8052 10492 8116
rect 10556 8052 10572 8116
rect 10636 8052 10652 8116
rect 10716 8052 10732 8116
rect 10796 8052 10812 8116
rect 10876 8052 10892 8116
rect 10956 8052 10972 8116
rect 11036 8052 11044 8116
rect 10244 8036 11044 8052
rect 10244 7972 10252 8036
rect 10316 7972 10332 8036
rect 10396 7972 10412 8036
rect 10476 7972 10492 8036
rect 10556 7972 10572 8036
rect 10636 7972 10652 8036
rect 10716 7972 10732 8036
rect 10796 7972 10812 8036
rect 10876 7972 10892 8036
rect 10956 7972 10972 8036
rect 11036 7972 11044 8036
rect 10244 7956 11044 7972
rect 10244 7892 10252 7956
rect 10316 7892 10332 7956
rect 10396 7892 10412 7956
rect 10476 7892 10492 7956
rect 10556 7892 10572 7956
rect 10636 7892 10652 7956
rect 10716 7892 10732 7956
rect 10796 7892 10812 7956
rect 10876 7892 10892 7956
rect 10956 7892 10972 7956
rect 11036 7892 11044 7956
rect 10244 7876 11044 7892
rect 10244 7812 10252 7876
rect 10316 7812 10332 7876
rect 10396 7812 10412 7876
rect 10476 7812 10492 7876
rect 10556 7812 10572 7876
rect 10636 7812 10652 7876
rect 10716 7812 10732 7876
rect 10796 7812 10812 7876
rect 10876 7812 10892 7876
rect 10956 7812 10972 7876
rect 11036 7812 11044 7876
rect 10244 1932 11044 7812
rect 10244 1868 10252 1932
rect 10316 1868 10332 1932
rect 10396 1868 10412 1932
rect 10476 1868 10492 1932
rect 10556 1868 10572 1932
rect 10636 1868 10652 1932
rect 10716 1868 10732 1932
rect 10796 1868 10812 1932
rect 10876 1868 10892 1932
rect 10956 1868 10972 1932
rect 11036 1868 11044 1932
rect 10244 1852 11044 1868
rect 10244 1788 10252 1852
rect 10316 1788 10332 1852
rect 10396 1788 10412 1852
rect 10476 1788 10492 1852
rect 10556 1788 10572 1852
rect 10636 1788 10652 1852
rect 10716 1788 10732 1852
rect 10796 1788 10812 1852
rect 10876 1788 10892 1852
rect 10956 1788 10972 1852
rect 11036 1788 11044 1852
rect 10244 1772 11044 1788
rect 10244 1708 10252 1772
rect 10316 1708 10332 1772
rect 10396 1708 10412 1772
rect 10476 1708 10492 1772
rect 10556 1708 10572 1772
rect 10636 1708 10652 1772
rect 10716 1708 10732 1772
rect 10796 1708 10812 1772
rect 10876 1708 10892 1772
rect 10956 1708 10972 1772
rect 11036 1708 11044 1772
rect 10244 1692 11044 1708
rect 10244 1628 10252 1692
rect 10316 1628 10332 1692
rect 10396 1628 10412 1692
rect 10476 1628 10492 1692
rect 10556 1628 10572 1692
rect 10636 1628 10652 1692
rect 10716 1628 10732 1692
rect 10796 1628 10812 1692
rect 10876 1628 10892 1692
rect 10956 1628 10972 1692
rect 11036 1628 11044 1692
rect 10244 1612 11044 1628
rect 10244 1548 10252 1612
rect 10316 1548 10332 1612
rect 10396 1548 10412 1612
rect 10476 1548 10492 1612
rect 10556 1548 10572 1612
rect 10636 1548 10652 1612
rect 10716 1548 10732 1612
rect 10796 1548 10812 1612
rect 10876 1548 10892 1612
rect 10956 1548 10972 1612
rect 11036 1548 11044 1612
rect 10244 1532 11044 1548
rect 10244 1468 10252 1532
rect 10316 1468 10332 1532
rect 10396 1468 10412 1532
rect 10476 1468 10492 1532
rect 10556 1468 10572 1532
rect 10636 1468 10652 1532
rect 10716 1468 10732 1532
rect 10796 1468 10812 1532
rect 10876 1468 10892 1532
rect 10956 1468 10972 1532
rect 11036 1468 11044 1532
rect 10244 1452 11044 1468
rect 10244 1388 10252 1452
rect 10316 1388 10332 1452
rect 10396 1388 10412 1452
rect 10476 1388 10492 1452
rect 10556 1388 10572 1452
rect 10636 1388 10652 1452
rect 10716 1388 10732 1452
rect 10796 1388 10812 1452
rect 10876 1388 10892 1452
rect 10956 1388 10972 1452
rect 11036 1388 11044 1452
rect 10244 1372 11044 1388
rect 10244 1308 10252 1372
rect 10316 1308 10332 1372
rect 10396 1308 10412 1372
rect 10476 1308 10492 1372
rect 10556 1308 10572 1372
rect 10636 1308 10652 1372
rect 10716 1308 10732 1372
rect 10796 1308 10812 1372
rect 10876 1308 10892 1372
rect 10956 1308 10972 1372
rect 11036 1308 11044 1372
rect 10244 1292 11044 1308
rect 10244 1228 10252 1292
rect 10316 1228 10332 1292
rect 10396 1228 10412 1292
rect 10476 1228 10492 1292
rect 10556 1228 10572 1292
rect 10636 1228 10652 1292
rect 10716 1228 10732 1292
rect 10796 1228 10812 1292
rect 10876 1228 10892 1292
rect 10956 1228 10972 1292
rect 11036 1228 11044 1292
rect 10244 1212 11044 1228
rect 10244 1148 10252 1212
rect 10316 1148 10332 1212
rect 10396 1148 10412 1212
rect 10476 1148 10492 1212
rect 10556 1148 10572 1212
rect 10636 1148 10652 1212
rect 10716 1148 10732 1212
rect 10796 1148 10812 1212
rect 10876 1148 10892 1212
rect 10956 1148 10972 1212
rect 11036 1148 11044 1212
rect 10244 1140 11044 1148
rect 11384 792 12184 8952
rect 11384 728 11392 792
rect 11456 728 11472 792
rect 11536 728 11552 792
rect 11616 728 11632 792
rect 11696 728 11712 792
rect 11776 728 11792 792
rect 11856 728 11872 792
rect 11936 728 11952 792
rect 12016 728 12032 792
rect 12096 728 12112 792
rect 12176 728 12184 792
rect 11384 712 12184 728
rect 11384 648 11392 712
rect 11456 648 11472 712
rect 11536 648 11552 712
rect 11616 648 11632 712
rect 11696 648 11712 712
rect 11776 648 11792 712
rect 11856 648 11872 712
rect 11936 648 11952 712
rect 12016 648 12032 712
rect 12096 648 12112 712
rect 12176 648 12184 712
rect 11384 632 12184 648
rect 11384 568 11392 632
rect 11456 568 11472 632
rect 11536 568 11552 632
rect 11616 568 11632 632
rect 11696 568 11712 632
rect 11776 568 11792 632
rect 11856 568 11872 632
rect 11936 568 11952 632
rect 12016 568 12032 632
rect 12096 568 12112 632
rect 12176 568 12184 632
rect 11384 552 12184 568
rect 11384 488 11392 552
rect 11456 488 11472 552
rect 11536 488 11552 552
rect 11616 488 11632 552
rect 11696 488 11712 552
rect 11776 488 11792 552
rect 11856 488 11872 552
rect 11936 488 11952 552
rect 12016 488 12032 552
rect 12096 488 12112 552
rect 12176 488 12184 552
rect 11384 472 12184 488
rect 11384 408 11392 472
rect 11456 408 11472 472
rect 11536 408 11552 472
rect 11616 408 11632 472
rect 11696 408 11712 472
rect 11776 408 11792 472
rect 11856 408 11872 472
rect 11936 408 11952 472
rect 12016 408 12032 472
rect 12096 408 12112 472
rect 12176 408 12184 472
rect 11384 392 12184 408
rect 11384 328 11392 392
rect 11456 328 11472 392
rect 11536 328 11552 392
rect 11616 328 11632 392
rect 11696 328 11712 392
rect 11776 328 11792 392
rect 11856 328 11872 392
rect 11936 328 11952 392
rect 12016 328 12032 392
rect 12096 328 12112 392
rect 12176 328 12184 392
rect 11384 312 12184 328
rect 11384 248 11392 312
rect 11456 248 11472 312
rect 11536 248 11552 312
rect 11616 248 11632 312
rect 11696 248 11712 312
rect 11776 248 11792 312
rect 11856 248 11872 312
rect 11936 248 11952 312
rect 12016 248 12032 312
rect 12096 248 12112 312
rect 12176 248 12184 312
rect 11384 232 12184 248
rect 11384 168 11392 232
rect 11456 168 11472 232
rect 11536 168 11552 232
rect 11616 168 11632 232
rect 11696 168 11712 232
rect 11776 168 11792 232
rect 11856 168 11872 232
rect 11936 168 11952 232
rect 12016 168 12032 232
rect 12096 168 12112 232
rect 12176 168 12184 232
rect 11384 152 12184 168
rect 11384 88 11392 152
rect 11456 88 11472 152
rect 11536 88 11552 152
rect 11616 88 11632 152
rect 11696 88 11712 152
rect 11776 88 11792 152
rect 11856 88 11872 152
rect 11936 88 11952 152
rect 12016 88 12032 152
rect 12096 88 12112 152
rect 12176 88 12184 152
rect 11384 72 12184 88
rect 11384 8 11392 72
rect 11456 8 11472 72
rect 11536 8 11552 72
rect 11616 8 11632 72
rect 11696 8 11712 72
rect 11776 8 11792 72
rect 11856 8 11872 72
rect 11936 8 11952 72
rect 12016 8 12032 72
rect 12096 8 12112 72
rect 12176 8 12184 72
rect 11384 0 12184 8
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3516 0 1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1624635492
transform 1 0 3516 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3240 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 3240 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5540 0 1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4620 0 1 3784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1624635492
transform 1 0 4620 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x9_B1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5356 0 1 3784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1624635492
transform 1 0 6000 0 1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6736 0 -1 3784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6368 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1624635492
transform 1 0 6000 0 -1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5724 0 -1 3784
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5908 0 1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12
timestamp 1624635492
transform 1 0 5908 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  x9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6368 0 1 3784
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6460 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1624635492
transform 1 0 7656 0 1 3784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1624635492
transform 1 0 7012 0 1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1624635492
transform 1 0 7564 0 -1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44
timestamp 1624635492
transform 1 0 7288 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 7564 0 -1 3784
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8208 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1624635492
transform 1 0 7380 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_56
timestamp 1624635492
transform 1 0 8392 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1624635492
transform 1 0 8208 0 -1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1624635492
transform 1 0 8576 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 8944 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 8944 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624635492
transform 1 0 3516 0 -1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 3240 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_21
timestamp 1624635492
transform 1 0 5172 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1624635492
transform 1 0 4620 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x6_B1
timestamp 1624635492
transform 1 0 4988 0 -1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__inv_1  x15
timestamp 1624635492
transform 1 0 5540 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_28
timestamp 1624635492
transform 1 0 5816 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  x6
timestamp 1624635492
transform 1 0 6184 0 -1 4872
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_50
timestamp 1624635492
transform 1 0 7840 0 -1 4872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1624635492
transform 1 0 6828 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7196 0 -1 4872
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_2_58
timestamp 1624635492
transform 1 0 8576 0 -1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1624635492
transform 1 0 8392 0 -1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1624635492
transform 1 0 8484 0 -1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 8944 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_12
timestamp 1624635492
transform 1 0 4344 0 1 4872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1624635492
transform 1 0 3792 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 4344 0 1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3792 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 3240 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1624635492
transform 1 0 5540 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_20
timestamp 1624635492
transform 1 0 5080 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x15_A
timestamp 1624635492
transform -1 0 5540 0 1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1624635492
transform 1 0 6000 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16
timestamp 1624635492
transform 1 0 5908 0 1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__a221oi_1  x8
timestamp 1624635492
transform 1 0 6368 0 1 4872
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_49
timestamp 1624635492
transform 1 0 7748 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_41
timestamp 1624635492
transform 1 0 7012 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7380 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_55
timestamp 1624635492
transform 1 0 8300 0 1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform 1 0 8116 0 1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 8944 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 3516 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 3240 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 4620 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1624635492
transform 1 0 6460 0 -1 5960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_27
timestamp 1624635492
transform 1 0 5724 0 -1 5960
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  x11
timestamp 1624635492
transform 1 0 6644 0 -1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp 1624635492
transform 1 0 7748 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1624635492
transform 1 0 7012 0 -1 5960
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform -1 0 8116 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1624635492
transform 1 0 8576 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1624635492
transform 1 0 8116 0 -1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1624635492
transform 1 0 8484 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 8944 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_12
timestamp 1624635492
transform 1 0 4344 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1624635492
transform 1 0 3792 0 1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 4344 0 1 5960
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 3516 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 3240 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1624635492
transform 1 0 5448 0 1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1624635492
transform 1 0 6000 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_28
timestamp 1624635492
transform 1 0 5816 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18
timestamp 1624635492
transform 1 0 5908 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_50
timestamp 1624635492
transform 1 0 7840 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_42
timestamp 1624635492
transform 1 0 7104 0 1 5960
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1624635492
transform 1 0 7932 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_54
timestamp 1624635492
transform 1 0 8208 0 1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1624635492
transform 1 0 8576 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 8944 0 1 5960
box -38 -48 314 592
<< labels >>
rlabel metal2 s 9336 4954 10136 5178 6 INN
port 0 nsew signal input
rlabel metal2 s 9336 2286 10136 2510 6 INP
port 1 nsew signal input
rlabel metal2 s 9336 7622 10136 7846 6 Q
port 2 nsew signal tristate
rlabel metal2 s 2136 7622 2936 7846 6 VDD
port 3 nsew signal input
rlabel metal2 s 2136 4954 2936 5178 6 VSS
port 4 nsew signal input
rlabel metal2 s 2136 2286 2936 2510 6 clk
port 5 nsew signal input
rlabel metal3 s 1140 7804 11044 8604 6 vccd2
port 6 nsew power bidirectional
rlabel metal3 s 1140 1140 11044 1940 6 vccd2
port 7 nsew power bidirectional
rlabel metal4 s 7857 0 8277 9744 6 vccd2
port 8 nsew power bidirectional
rlabel metal4 s 5926 0 6346 9744 6 vccd2
port 9 nsew power bidirectional
rlabel metal4 s 3995 0 4415 9744 6 vccd2
port 10 nsew power bidirectional
rlabel metal4 s 10244 1140 11044 8604 6 vccd2
port 11 nsew power bidirectional
rlabel metal4 s 1140 1140 1940 8604 4 vccd2
port 12 nsew power bidirectional
rlabel metal3 s 0 8944 12184 9744 6 vssd2
port 13 nsew ground bidirectional
rlabel metal3 s 0 0 12184 800 8 vssd2
port 14 nsew ground bidirectional
rlabel metal4 s 11384 0 12184 9744 6 vssd2
port 15 nsew ground bidirectional
rlabel metal4 s 6891 0 7311 9744 6 vssd2
port 16 nsew ground bidirectional
rlabel metal4 s 4961 0 5381 9744 6 vssd2
port 17 nsew ground bidirectional
rlabel metal4 s 0 0 800 9744 4 vssd2
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12184 9744
<< end >>
