magic
tech sky130A
magscale 1 2
timestamp 1626450099
<< checkpaint >>
rect -1266 -7308 14774 6984
<< locali >>
rect 232 5402 290 5482
rect 13190 3488 13240 3490
rect 10096 3434 13240 3488
rect 10096 3428 12540 3434
rect 7408 2028 7508 3300
rect 7408 1994 7442 2028
rect 7476 1994 7508 2028
rect 7408 1962 7508 1994
rect 3880 1546 3940 1602
rect 3880 1420 3948 1546
rect 7398 1424 7500 1478
rect 3880 1414 3952 1420
rect 3884 1069 3952 1414
rect 3884 1035 3896 1069
rect 3930 1035 3952 1069
rect 3884 1022 3952 1035
rect 7398 1390 7432 1424
rect 7466 1390 7500 1424
rect 7398 1034 7500 1390
rect 7390 862 7500 1034
rect 3880 741 3948 764
rect 800 468 844 736
rect 3880 707 3898 741
rect 3932 707 3948 741
rect 788 464 852 468
rect 788 430 805 464
rect 839 430 852 464
rect 788 424 852 430
rect 3880 386 3948 707
rect 794 226 858 234
rect 794 192 808 226
rect 842 192 858 226
rect 794 186 858 192
rect 20 0 316 46
rect 266 -280 316 0
rect 800 -296 846 186
rect 788 -306 864 -296
rect 788 -317 866 -306
rect 788 -351 809 -317
rect 843 -351 866 -317
rect 40 -572 90 -358
rect 788 -360 866 -351
rect 790 -370 866 -360
rect 786 -539 860 -518
rect 40 -622 282 -572
rect 786 -573 806 -539
rect 840 -573 860 -539
rect 786 -592 860 -573
rect 798 -754 844 -592
rect 3880 -602 3950 386
rect 7390 -32 7492 862
rect 13190 806 13242 3434
rect 13188 782 13242 806
rect 13188 556 13240 782
rect 13358 272 13514 284
rect 13358 238 13370 272
rect 13404 238 13514 272
rect 13358 224 13514 238
rect 10958 64 11044 158
rect 7390 -120 7498 -32
rect 3878 -621 3956 -602
rect 3878 -655 3898 -621
rect 3932 -655 3956 -621
rect 3878 -676 3956 -655
rect 796 -1042 846 -754
rect 796 -1070 872 -1042
rect 798 -1106 872 -1070
rect 3884 -1071 3954 -1052
rect 3884 -1105 3900 -1071
rect 3934 -1105 3954 -1071
rect 3884 -1584 3954 -1105
rect 7396 -1152 7498 -120
rect 7396 -1186 7428 -1152
rect 7462 -1186 7498 -1152
rect 7396 -1222 7498 -1186
rect 7398 -1678 7492 -1626
rect 7398 -1712 7422 -1678
rect 7456 -1712 7492 -1678
rect 7398 -2702 7492 -1712
rect 13196 -2524 13258 -194
rect 9972 -2584 13266 -2524
rect 10 -6048 72 -5968
<< viali >>
rect 7442 1994 7476 2028
rect 3896 1035 3930 1069
rect 7432 1390 7466 1424
rect 3898 707 3932 741
rect 805 430 839 464
rect 808 192 842 226
rect 809 -351 843 -317
rect 806 -573 840 -539
rect 13370 238 13404 272
rect 3898 -655 3932 -621
rect 3900 -1105 3934 -1071
rect 7428 -1186 7462 -1152
rect 7422 -1712 7456 -1678
<< metal1 >>
rect 7392 2028 7506 2070
rect 7392 1994 7442 2028
rect 7476 1994 7506 2028
rect 7392 1424 7506 1994
rect 7392 1390 7432 1424
rect 7466 1390 7506 1424
rect 7392 1356 7506 1390
rect 3884 1084 3930 1130
rect 3880 1069 3948 1084
rect 3880 1035 3896 1069
rect 3930 1035 3948 1069
rect 3880 741 3948 1035
rect 3880 707 3898 741
rect 3932 707 3948 741
rect 3880 686 3948 707
rect 11832 591 11926 606
rect 11832 539 11859 591
rect 11911 539 11926 591
rect 11832 528 11926 539
rect 798 470 844 502
rect 798 468 846 470
rect 788 464 852 468
rect 788 430 805 464
rect 839 430 852 464
rect 788 424 852 430
rect 800 234 846 424
rect 13368 238 13370 272
rect 13404 238 13406 272
rect 794 226 858 234
rect 794 192 808 226
rect 842 192 858 226
rect 794 186 858 192
rect 11092 -208 11208 -132
rect 11092 -260 11096 -208
rect 11148 -260 11208 -208
rect 11092 -278 11208 -260
rect 788 -306 864 -296
rect 788 -317 866 -306
rect 788 -351 809 -317
rect 843 -351 866 -317
rect 788 -360 866 -351
rect 790 -370 866 -360
rect 800 -518 846 -370
rect 786 -539 860 -518
rect 786 -573 806 -539
rect 840 -573 860 -539
rect 786 -592 860 -573
rect 3882 -602 3952 -596
rect 3878 -621 3956 -602
rect 3878 -655 3898 -621
rect 3932 -655 3956 -621
rect 3878 -676 3956 -655
rect 3882 -1071 3952 -676
rect 3882 -1105 3900 -1071
rect 3934 -1105 3952 -1071
rect 3882 -1128 3952 -1105
rect 7396 -1134 7500 -1118
rect 7390 -1152 7500 -1134
rect 7390 -1186 7428 -1152
rect 7462 -1186 7500 -1152
rect 7390 -1218 7500 -1186
rect 7390 -1678 7492 -1218
rect 7390 -1712 7422 -1678
rect 7456 -1712 7492 -1678
rect 7390 -1750 7492 -1712
<< via1 >>
rect 11859 539 11911 591
rect 11096 -260 11148 -208
<< metal2 >>
rect 11848 687 11924 702
rect 11848 631 11860 687
rect 11916 631 11924 687
rect 11848 591 11924 631
rect 11848 539 11859 591
rect 11911 539 11924 591
rect 11848 530 11924 539
rect 6532 -216 6570 218
rect 11090 -208 11164 -192
rect 11090 -216 11096 -208
rect 6532 -260 11096 -216
rect 11148 -260 11164 -208
rect 6532 -264 11164 -260
rect 6532 -5868 6570 -264
<< via2 >>
rect 11860 631 11916 687
<< metal3 >>
rect 11850 826 11926 840
rect 11850 772 11860 826
rect 11848 762 11860 772
rect 11924 762 11926 826
rect 11848 687 11926 762
rect 11848 631 11860 687
rect 11916 631 11926 687
rect 11848 620 11926 631
<< via3 >>
rect 11860 762 11924 826
<< metal4 >>
rect 6842 962 6920 3000
rect 6820 884 11926 962
rect 6842 -774 6920 884
rect 11850 826 11926 884
rect 11850 762 11860 826
rect 11924 762 11926 826
rect 11850 750 11926 762
use switch_layout  switch_layout_0
timestamp 1626450099
transform 1 0 10954 0 1 -454
box 40 154 2460 1180
use res250_layout  res250_layout_0
timestamp 1626450099
transform 0 -1 -48 1 0 -668
box 202 -342 510 -90
use 3bitdac_layout  3bitdac_layout_0
timestamp 1626450099
transform 1 0 54 0 1 3060
box -54 -3060 10120 2664
use 3bitdac_layout  3bitdac_layout_1
timestamp 1626450099
transform 1 0 48 0 1 -2954
box -54 -3060 10120 2664
<< labels >>
rlabel locali s 10594 3462 10594 3462 4 x1_out_v
port 1 nsew
rlabel locali s 10334 -2560 10334 -2560 4 x2_out_v
port 2 nsew
rlabel locali s 254 5442 254 5442 4 inp1
port 3 nsew
rlabel locali s 40 -6024 40 -6024 4 inp2
port 4 nsew
rlabel locali s 292 -138 292 -138 4 x1_vref5
port 5 nsew
rlabel locali s 202 -604 202 -604 4 x2_vref1
port 6 nsew
rlabel locali s 818 -52 818 -52 4 d0
port 7 nsew
rlabel locali s 3908 -10 3908 -10 4 d1
port 8 nsew
rlabel locali s 7436 126 7436 126 4 d2
port 9 nsew
rlabel locali s 10976 102 10976 102 4 d3
port 10 nsew
rlabel locali s 13434 248 13434 248 4 out_v
port 11 nsew
rlabel metal2 s 10968 -246 10968 -246 4 gnd!
port 12 nsew
rlabel metal4 s 11590 914 11590 914 4 vdd!
port 13 nsew
<< properties >>
string GDS_FILE gds/adc_wrapper.gds
string GDS_END 36634
string GDS_START 29978
<< end >>
