magic
tech sky130A
magscale 1 2
timestamp 1626375338
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 1104 2128 68816 67504
<< metal2 >>
rect 17498 69200 17554 70000
rect 52458 69200 52514 70000
rect 17498 0 17554 800
rect 52458 0 52514 800
<< obsm2 >>
rect 1398 69144 17442 69200
rect 17610 69144 52402 69200
rect 52570 69144 68154 69200
rect 1398 856 68154 69144
rect 1398 800 17442 856
rect 17610 800 52402 856
rect 52570 800 68154 856
<< metal3 >>
rect 0 66376 800 66496
rect 0 59440 800 59560
rect 69200 58216 70000 58336
rect 0 52368 800 52488
rect 0 45432 800 45552
rect 0 38360 800 38480
rect 69200 34824 70000 34944
rect 0 31424 800 31544
rect 0 24352 800 24472
rect 0 17416 800 17536
rect 69200 11568 70000 11688
rect 0 10344 800 10464
rect 0 3408 800 3528
<< obsm3 >>
rect 800 66576 69200 67489
rect 880 66296 69200 66576
rect 800 59640 69200 66296
rect 880 59360 69200 59640
rect 800 58416 69200 59360
rect 800 58136 69120 58416
rect 800 52568 69200 58136
rect 880 52288 69200 52568
rect 800 45632 69200 52288
rect 880 45352 69200 45632
rect 800 38560 69200 45352
rect 880 38280 69200 38560
rect 800 35024 69200 38280
rect 800 34744 69120 35024
rect 800 31624 69200 34744
rect 880 31344 69200 31624
rect 800 24552 69200 31344
rect 880 24272 69200 24552
rect 800 17616 69200 24272
rect 880 17336 69200 17616
rect 800 11768 69200 17336
rect 800 11488 69120 11768
rect 800 10544 69200 11488
rect 880 10264 69200 10544
rect 800 3608 69200 10264
rect 880 3328 69200 3608
rect 800 2000 69200 3328
<< metal4 >>
rect 4018 2128 4718 67504
rect 5058 2176 5758 67456
rect 8518 2128 9218 67504
rect 9558 2176 10258 67456
rect 13018 2128 13718 67504
rect 14058 2176 14758 67456
rect 17518 2128 18218 67504
rect 18558 2176 19258 67456
rect 22018 2176 22718 67504
rect 23058 2176 23758 67456
rect 26518 2176 27218 67504
rect 27558 2176 28258 67456
rect 31018 2176 31718 67504
rect 32058 2176 32758 67456
rect 35518 2176 36218 67504
rect 36558 2176 37258 67456
rect 40018 2128 40718 67504
rect 41058 2176 41758 67456
rect 44518 2128 45218 67504
rect 45558 2176 46258 67456
rect 49018 2128 49718 67504
rect 50058 2176 50758 67456
rect 53518 2128 54218 67504
rect 54558 2176 55258 67456
rect 58018 2128 58718 67504
rect 59058 2176 59758 67456
rect 62518 2128 63218 67504
rect 63558 2176 64258 67456
rect 67018 2128 67718 67504
<< metal5 >>
rect -2236 70476 72156 70796
rect -1576 69816 71496 70136
rect -916 69156 70836 69476
rect -256 68496 70176 68816
rect -916 66570 70836 66890
rect -2236 51960 72156 52280
rect -916 51252 70836 51572
rect -2236 36642 72156 36962
rect -916 35934 70836 36254
rect -2236 21324 72156 21644
rect -916 20616 70836 20936
rect -2236 6006 72156 6326
rect -916 5298 70836 5618
rect -256 816 70176 1136
rect -916 156 70836 476
rect -1576 -504 71496 -184
rect -2236 -1164 72156 -844
<< labels >>
rlabel metal3 s 69200 34824 70000 34944 6 INN
port 1 nsew signal input
rlabel metal3 s 69200 11568 70000 11688 6 INP
port 2 nsew signal input
rlabel metal3 s 69200 58216 70000 58336 6 Q
port 3 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 clk
port 4 nsew signal input
rlabel metal2 s 52458 69200 52514 70000 6 cmp
port 5 nsew signal input
rlabel metal2 s 17498 69200 17554 70000 6 cmp_sel
port 6 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 data[0]
port 7 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 data[1]
port 8 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 data[2]
port 9 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 data[3]
port 10 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 data[4]
port 11 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 data[5]
port 12 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 data[6]
port 13 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 data[7]
port 14 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 done
port 15 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 rstn
port 16 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 start
port 17 nsew signal input
rlabel metal4 s 67018 2128 67718 67504 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 58018 2128 58718 67504 6 vccd1
port 19 nsew power bidirectional
rlabel metal4 s 49018 2128 49718 67504 6 vccd1
port 20 nsew power bidirectional
rlabel metal4 s 40018 2128 40718 67504 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 31018 2176 31718 67504 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 22018 2176 22718 67504 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 13018 2128 13718 67504 6 vccd1
port 24 nsew power bidirectional
rlabel metal4 s 4018 2128 4718 67504 6 vccd1
port 25 nsew power bidirectional
rlabel metal5 s -256 68496 70176 68816 6 vccd1
port 26 nsew power bidirectional
rlabel metal5 s -916 66570 70836 66890 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -916 35934 70836 36254 6 vccd1
port 28 nsew power bidirectional
rlabel metal5 s -916 5298 70836 5618 6 vccd1
port 29 nsew power bidirectional
rlabel metal5 s -256 816 70176 1136 6 vccd1
port 30 nsew power bidirectional
rlabel metal4 s 62518 2128 63218 67504 6 vssd1
port 31 nsew ground bidirectional
rlabel metal4 s 53518 2128 54218 67504 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 44518 2128 45218 67504 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 35518 2176 36218 67504 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 26518 2176 27218 67504 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 17518 2128 18218 67504 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 8518 2128 9218 67504 6 vssd1
port 37 nsew ground bidirectional
rlabel metal5 s -916 69156 70836 69476 6 vssd1
port 38 nsew ground bidirectional
rlabel metal5 s -916 51252 70836 51572 6 vssd1
port 39 nsew ground bidirectional
rlabel metal5 s -916 20616 70836 20936 6 vssd1
port 40 nsew ground bidirectional
rlabel metal5 s -916 156 70836 476 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 59058 2176 59758 67456 6 vccd2
port 42 nsew power bidirectional
rlabel metal4 s 50058 2176 50758 67456 6 vccd2
port 43 nsew power bidirectional
rlabel metal4 s 41058 2176 41758 67456 6 vccd2
port 44 nsew power bidirectional
rlabel metal4 s 32058 2176 32758 67456 6 vccd2
port 45 nsew power bidirectional
rlabel metal4 s 23058 2176 23758 67456 6 vccd2
port 46 nsew power bidirectional
rlabel metal4 s 14058 2176 14758 67456 6 vccd2
port 47 nsew power bidirectional
rlabel metal4 s 5058 2176 5758 67456 6 vccd2
port 48 nsew power bidirectional
rlabel metal5 s -1576 69816 71496 70136 6 vccd2
port 49 nsew power bidirectional
rlabel metal5 s -2236 36642 72156 36962 6 vccd2
port 50 nsew power bidirectional
rlabel metal5 s -2236 6006 72156 6326 6 vccd2
port 51 nsew power bidirectional
rlabel metal5 s -1576 -504 71496 -184 8 vccd2
port 52 nsew power bidirectional
rlabel metal4 s 63558 2176 64258 67456 6 vssd2
port 53 nsew ground bidirectional
rlabel metal4 s 54558 2176 55258 67456 6 vssd2
port 54 nsew ground bidirectional
rlabel metal4 s 45558 2176 46258 67456 6 vssd2
port 55 nsew ground bidirectional
rlabel metal4 s 36558 2176 37258 67456 6 vssd2
port 56 nsew ground bidirectional
rlabel metal4 s 27558 2176 28258 67456 6 vssd2
port 57 nsew ground bidirectional
rlabel metal4 s 18558 2176 19258 67456 6 vssd2
port 58 nsew ground bidirectional
rlabel metal4 s 9558 2176 10258 67456 6 vssd2
port 59 nsew ground bidirectional
rlabel metal5 s -2236 70476 72156 70796 6 vssd2
port 60 nsew ground bidirectional
rlabel metal5 s -2236 51960 72156 52280 6 vssd2
port 61 nsew ground bidirectional
rlabel metal5 s -2236 21324 72156 21644 6 vssd2
port 62 nsew ground bidirectional
rlabel metal5 s -2236 -1164 72156 -844 8 vssd2
port 63 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 70000 70000
string LEFview TRUE
string GDS_FILE /project/openlane/ACMP_SAR/runs/ACMP_SAR/results/magic/ACMP_SAR.gds
string GDS_END 3180786
string GDS_START 489608
<< end >>

