module ACMP_HVL (INN,
    INP,
    Q,
    clk,
    vccd2,
    vssd2);
 input INN;
 input INP;
 output Q;
 input clk;
 input vccd2;
 input vssd2;

 sky130_fd_sc_hvl__inv_1 x0 (.A(clk),
    .Y(\x2.CLK ),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__nand3_1 \x1.x1  (.A(clk),
    .B(INP),
    .C(\x1.Q0 ),
    .Y(\x1.Q0b ),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__nand3_1 \x1.x2  (.A(clk),
    .B(INN),
    .C(\x1.Q0b ),
    .Y(\x1.Q0 ),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__inv_4 \x1.x3  (.A(\x1.Q0 ),
    .Y(\x1.Qb ),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__inv_4 \x1.x4  (.A(\x1.Q0b ),
    .Y(\x1.Q ),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__nor3_1 \x2.x1  (.A(\x2.CLK ),
    .B(INP),
    .C(\x2.Q ),
    .Y(\x2.Qb ),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__nor3_1 \x2.x2  (.A(\x2.CLK ),
    .B(INN),
    .C(\x2.Qb ),
    .Y(\x2.Q ),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__nor3_1 x5 (.A(\x1.Qb ),
    .B(\x2.Qb ),
    .C(Qb),
    .Y(Q),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__nor3_1 x6 (.A(\x1.Q ),
    .B(\x2.Q ),
    .C(Q),
    .Y(Qb),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__diode_2 \ANTENNA_x2.x2_B  (.DIODE(INN),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__diode_2 \ANTENNA_x1.x2_B  (.DIODE(INN),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__diode_2 \ANTENNA_x2.x1_B  (.DIODE(INP),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__diode_2 \ANTENNA_x1.x1_B  (.DIODE(INP),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__diode_2 \ANTENNA_x1.x2_A  (.DIODE(clk),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__diode_2 \ANTENNA_x1.x1_A  (.DIODE(clk),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__diode_2 ANTENNA_x0_A (.DIODE(clk),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_0_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_0_116 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_0_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_0_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_0_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_1 FILLER_1_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_1_107 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_1_118 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_124 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_1_132 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_1_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_2_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_2_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_2_100 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_2_107 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_2_118 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_2_129 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_2_135 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_2_139 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_1 FILLER_2_141 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_3_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_3_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_3_100 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_3_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_3_108 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_3_118 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_3_129 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_3_135 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_3_139 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_1 FILLER_3_141 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_4_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_4_108 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_4_118 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_4_129 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_4_137 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_1 FILLER_4_141 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_1 FILLER_5_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_5_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_5_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_5_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_6_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_6_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_6_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_7_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_7_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_7_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_8_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_8_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_8_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_9_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_9_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_9_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_10_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_10_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_10_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_11_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_11_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_11_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_12_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_12_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_12_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_13_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_13_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_13_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_14_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_14_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_14_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_56 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_64 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_72 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_80 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_96 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_104 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_120 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_8 FILLER_15_128 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__decap_4 FILLER_15_136 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hvl__fill_2 FILLER_15_140 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
endmodule
