magic
tech sky130A
magscale 1 2
timestamp 1626450099
<< checkpaint >>
rect -1298 -1308 3230 1852
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 201 773 203
rect 1747 201 1931 203
rect 1 21 1931 201
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 762 47 792 175
rect 851 47 881 175
rect 935 47 965 175
rect 1175 47 1205 175
rect 1272 47 1302 175
rect 1399 47 1429 175
rect 1483 47 1513 175
rect 1723 47 1753 175
rect 1823 47 1853 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 762 297 792 497
rect 1007 297 1037 497
rect 1091 297 1121 497
rect 1175 297 1205 497
rect 1272 297 1302 497
rect 1555 297 1585 497
rect 1639 297 1669 497
rect 1723 297 1753 497
rect 1823 297 1853 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 163 177
rect 109 67 119 101
rect 153 67 163 101
rect 109 47 163 67
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 109 331 177
rect 277 75 287 109
rect 321 75 331 109
rect 277 47 331 75
rect 361 93 415 177
rect 361 59 371 93
rect 405 59 415 93
rect 361 47 415 59
rect 445 101 499 177
rect 445 67 455 101
rect 489 67 499 101
rect 445 47 499 67
rect 529 93 583 177
rect 529 59 539 93
rect 573 59 583 93
rect 529 47 583 59
rect 613 109 667 177
rect 613 75 623 109
rect 657 75 667 109
rect 613 47 667 75
rect 697 175 747 177
rect 1773 175 1823 177
rect 697 93 762 175
rect 697 59 707 93
rect 741 59 762 93
rect 697 47 762 59
rect 792 93 851 175
rect 792 59 807 93
rect 841 59 851 93
rect 792 47 851 59
rect 881 161 935 175
rect 881 127 891 161
rect 925 127 935 161
rect 881 47 935 127
rect 965 93 1175 175
rect 965 59 975 93
rect 1009 59 1175 93
rect 965 47 1175 59
rect 1205 93 1272 175
rect 1205 59 1228 93
rect 1262 59 1272 93
rect 1205 47 1272 59
rect 1302 93 1399 175
rect 1302 59 1331 93
rect 1365 59 1399 93
rect 1302 47 1399 59
rect 1429 161 1483 175
rect 1429 127 1439 161
rect 1473 127 1483 161
rect 1429 47 1483 127
rect 1513 93 1723 175
rect 1513 59 1523 93
rect 1557 59 1723 93
rect 1513 47 1723 59
rect 1753 93 1823 175
rect 1753 59 1779 93
rect 1813 59 1823 93
rect 1753 47 1823 59
rect 1853 109 1905 177
rect 1853 75 1863 109
rect 1897 75 1905 109
rect 1853 47 1905 75
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 297 79 383
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 477 499 497
rect 445 443 455 477
rect 489 443 499 477
rect 445 409 499 443
rect 445 375 455 409
rect 489 375 499 409
rect 445 297 499 375
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 477 667 497
rect 613 443 623 477
rect 657 443 667 477
rect 613 409 667 443
rect 613 375 623 409
rect 657 375 667 409
rect 613 297 667 375
rect 697 485 762 497
rect 697 451 707 485
rect 741 451 762 485
rect 697 297 762 451
rect 792 485 1007 497
rect 792 451 807 485
rect 841 451 1007 485
rect 792 297 1007 451
rect 1037 401 1091 497
rect 1037 367 1047 401
rect 1081 367 1091 401
rect 1037 297 1091 367
rect 1121 485 1175 497
rect 1121 451 1131 485
rect 1165 451 1175 485
rect 1121 297 1175 451
rect 1205 485 1272 497
rect 1205 451 1215 485
rect 1249 451 1272 485
rect 1205 297 1272 451
rect 1302 485 1555 497
rect 1302 451 1312 485
rect 1346 451 1555 485
rect 1302 297 1555 451
rect 1585 401 1639 497
rect 1585 367 1595 401
rect 1629 367 1639 401
rect 1585 297 1639 367
rect 1669 485 1723 497
rect 1669 451 1679 485
rect 1713 451 1723 485
rect 1669 297 1723 451
rect 1753 485 1823 497
rect 1753 451 1779 485
rect 1813 451 1823 485
rect 1753 297 1823 451
rect 1853 477 1905 497
rect 1853 443 1863 477
rect 1897 443 1905 477
rect 1853 409 1905 443
rect 1853 375 1863 409
rect 1897 375 1905 409
rect 1853 297 1905 375
<< ndiffc >>
rect 35 59 69 93
rect 119 67 153 101
rect 203 59 237 93
rect 287 75 321 109
rect 371 59 405 93
rect 455 67 489 101
rect 539 59 573 93
rect 623 75 657 109
rect 707 59 741 93
rect 807 59 841 93
rect 891 127 925 161
rect 975 59 1009 93
rect 1228 59 1262 93
rect 1331 59 1365 93
rect 1439 127 1473 161
rect 1523 59 1557 93
rect 1779 59 1813 93
rect 1863 75 1897 109
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 119 443 153 477
rect 119 375 153 409
rect 203 451 237 485
rect 203 383 237 417
rect 287 443 321 477
rect 287 375 321 409
rect 371 451 405 485
rect 371 383 405 417
rect 455 443 489 477
rect 455 375 489 409
rect 539 451 573 485
rect 539 383 573 417
rect 623 443 657 477
rect 623 375 657 409
rect 707 451 741 485
rect 807 451 841 485
rect 1047 367 1081 401
rect 1131 451 1165 485
rect 1215 451 1249 485
rect 1312 451 1346 485
rect 1595 367 1629 401
rect 1679 451 1713 485
rect 1779 451 1813 485
rect 1863 443 1897 477
rect 1863 375 1897 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 762 497 792 523
rect 1007 497 1037 523
rect 1091 497 1121 523
rect 1175 497 1205 523
rect 1272 497 1302 523
rect 1555 497 1585 523
rect 1639 497 1669 523
rect 1723 497 1753 523
rect 1823 497 1853 523
rect 79 269 109 297
rect 163 269 193 297
rect 247 269 277 297
rect 331 269 361 297
rect 415 269 445 297
rect 499 269 529 297
rect 583 269 613 297
rect 667 269 697 297
rect 79 249 697 269
rect 762 265 792 297
rect 1007 282 1037 297
rect 1091 282 1121 297
rect 79 215 213 249
rect 247 215 281 249
rect 315 215 349 249
rect 383 215 417 249
rect 451 215 485 249
rect 519 215 553 249
rect 587 215 621 249
rect 655 215 697 249
rect 79 199 697 215
rect 749 249 804 265
rect 749 215 759 249
rect 793 215 804 249
rect 749 199 804 215
rect 851 249 965 265
rect 851 215 861 249
rect 895 215 965 249
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 762 175 792 199
rect 851 192 965 215
rect 1007 249 1121 282
rect 1175 265 1205 297
rect 1272 265 1302 297
rect 1555 282 1585 297
rect 1639 282 1669 297
rect 1007 215 1036 249
rect 1070 215 1121 249
rect 1007 199 1121 215
rect 1163 249 1217 265
rect 1163 215 1173 249
rect 1207 215 1217 249
rect 1163 199 1217 215
rect 1259 249 1326 265
rect 1259 215 1269 249
rect 1303 215 1326 249
rect 1259 199 1326 215
rect 1395 249 1513 265
rect 1395 215 1405 249
rect 1439 215 1513 249
rect 1395 199 1513 215
rect 1555 249 1669 282
rect 1555 215 1615 249
rect 1649 215 1669 249
rect 1555 199 1669 215
rect 1723 265 1753 297
rect 1823 265 1853 297
rect 1723 249 1781 265
rect 1723 215 1737 249
rect 1771 215 1781 249
rect 1723 199 1781 215
rect 1823 249 1887 265
rect 1823 215 1843 249
rect 1877 215 1887 249
rect 1823 199 1887 215
rect 851 175 881 192
rect 935 175 965 192
rect 1175 175 1205 199
rect 1272 175 1302 199
rect 1399 192 1513 199
rect 1399 175 1429 192
rect 1483 175 1513 192
rect 1723 175 1753 199
rect 1823 177 1853 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 762 21 792 47
rect 851 21 881 47
rect 935 21 965 47
rect 1175 21 1205 47
rect 1272 21 1302 47
rect 1399 21 1429 47
rect 1483 21 1513 47
rect 1723 21 1753 47
rect 1823 21 1853 47
<< polycont >>
rect 213 215 247 249
rect 281 215 315 249
rect 349 215 383 249
rect 417 215 451 249
rect 485 215 519 249
rect 553 215 587 249
rect 621 215 655 249
rect 759 215 793 249
rect 861 215 895 249
rect 1036 215 1070 249
rect 1173 215 1207 249
rect 1269 215 1303 249
rect 1405 215 1439 249
rect 1615 215 1649 249
rect 1737 215 1771 249
rect 1843 215 1877 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 119 477 153 493
rect 119 409 153 443
rect 187 485 253 527
rect 187 451 203 485
rect 237 451 253 485
rect 187 417 253 451
rect 187 383 203 417
rect 237 383 253 417
rect 287 477 321 493
rect 287 409 321 443
rect 119 349 153 375
rect 355 485 421 527
rect 355 451 371 485
rect 405 451 421 485
rect 355 417 421 451
rect 355 383 371 417
rect 405 383 421 417
rect 455 477 489 493
rect 455 409 489 443
rect 287 349 321 375
rect 523 485 589 527
rect 523 451 539 485
rect 573 451 589 485
rect 523 417 589 451
rect 523 383 539 417
rect 573 383 589 417
rect 623 477 657 493
rect 691 485 757 527
rect 1215 485 1249 527
rect 1763 485 1829 527
rect 691 451 707 485
rect 741 451 757 485
rect 791 451 807 485
rect 841 451 1131 485
rect 1165 451 1181 485
rect 1296 451 1312 485
rect 1346 451 1679 485
rect 1713 451 1729 485
rect 1763 451 1779 485
rect 1813 451 1829 485
rect 1863 477 1897 493
rect 623 409 657 443
rect 1215 435 1249 451
rect 1863 417 1897 443
rect 455 349 489 375
rect 1737 409 1897 417
rect 623 349 657 375
rect 119 315 657 349
rect 691 367 1047 401
rect 1081 367 1595 401
rect 1629 367 1645 401
rect 1737 383 1863 409
rect 119 161 163 315
rect 691 249 725 367
rect 1737 333 1771 383
rect 1863 359 1897 375
rect 197 215 213 249
rect 247 215 281 249
rect 315 215 349 249
rect 383 215 417 249
rect 451 215 485 249
rect 519 215 553 249
rect 587 215 621 249
rect 655 215 725 249
rect 691 161 725 215
rect 759 323 1207 333
rect 759 299 1134 323
rect 759 249 793 299
rect 1168 289 1207 323
rect 861 255 895 265
rect 892 249 895 255
rect 759 199 793 215
rect 861 199 895 215
rect 1036 249 1070 265
rect 119 127 657 161
rect 691 127 891 161
rect 925 153 950 161
rect 925 127 984 153
rect 1036 163 1070 215
rect 1134 249 1207 289
rect 1134 215 1173 249
rect 1134 199 1207 215
rect 1269 299 1771 333
rect 1269 249 1303 299
rect 1405 249 1439 265
rect 1269 199 1303 215
rect 1345 215 1405 233
rect 1345 199 1439 215
rect 1592 255 1649 265
rect 1626 249 1649 255
rect 1592 215 1615 221
rect 1592 199 1649 215
rect 1737 249 1771 299
rect 1345 163 1379 199
rect 1036 129 1379 163
rect 119 101 153 127
rect 18 59 35 93
rect 69 59 85 93
rect 18 17 85 59
rect 287 109 321 127
rect 119 51 153 67
rect 187 59 203 93
rect 237 59 253 93
rect 455 101 489 127
rect 287 59 321 75
rect 355 59 371 93
rect 405 59 421 93
rect 187 17 253 59
rect 355 17 421 59
rect 623 109 657 127
rect 455 51 489 67
rect 523 59 539 93
rect 573 59 589 93
rect 623 59 657 75
rect 691 59 707 93
rect 741 59 757 93
rect 791 59 807 93
rect 841 59 975 93
rect 1009 59 1025 93
rect 1061 85 1178 129
rect 1423 127 1439 161
rect 1473 153 1500 161
rect 1473 127 1534 153
rect 1737 163 1771 215
rect 1843 289 1868 323
rect 1843 249 1902 289
rect 1877 215 1902 249
rect 1843 199 1902 215
rect 1737 129 1897 163
rect 1863 109 1897 129
rect 1212 59 1228 93
rect 1262 59 1278 93
rect 1315 59 1331 93
rect 1365 59 1523 93
rect 1557 59 1573 93
rect 1763 59 1779 93
rect 1813 59 1829 93
rect 1863 59 1897 75
rect 523 17 589 59
rect 691 17 757 59
rect 1212 17 1278 59
rect 1763 17 1829 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1134 289 1168 323
rect 858 249 892 255
rect 858 221 861 249
rect 861 221 892 249
rect 950 153 984 187
rect 1592 249 1626 255
rect 1592 221 1615 249
rect 1615 221 1626 249
rect 1500 153 1534 187
rect 1868 289 1902 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 1122 323 1180 329
rect 1122 289 1134 323
rect 1168 320 1180 323
rect 1856 323 1914 329
rect 1856 320 1868 323
rect 1168 292 1868 320
rect 1168 289 1180 292
rect 1122 283 1180 289
rect 1856 289 1868 292
rect 1902 289 1914 323
rect 1856 283 1914 289
rect 846 255 904 261
rect 846 221 858 255
rect 892 252 904 255
rect 1580 255 1638 261
rect 1580 252 1592 255
rect 892 224 1592 252
rect 892 221 904 224
rect 846 215 904 221
rect 1580 221 1592 224
rect 1626 221 1638 255
rect 1580 215 1638 221
rect 938 187 996 193
rect 938 153 950 187
rect 984 184 996 187
rect 1488 187 1546 193
rect 1488 184 1500 187
rect 984 156 1500 184
rect 984 153 996 156
rect 938 147 996 153
rect 1488 153 1500 156
rect 1534 153 1546 187
rect 1488 147 1546 153
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel metal1 s 1868 289 1902 323 0 FreeSans 200 0 0 0 S
flabel metal1 s 1592 221 1626 255 0 FreeSans 200 0 0 0 A1
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
flabel locali s 1134 85 1168 119 0 FreeSans 200 0 0 0 A0
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 X
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 mux2_8
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE gds/adc_wrapper.gds
string GDS_END 157794
string GDS_START 145122
string path 0.000 2.720 9.660 2.720 
<< end >>
