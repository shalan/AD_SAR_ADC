VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ACMP
  CLASS BLOCK ;
  FOREIGN ACMP ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.920 BY 48.720 ;
  PIN INN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.680 24.770 50.680 25.890 ;
    END
  END INN
  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.680 11.430 50.680 12.550 ;
    END
  END INP
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.680 38.110 50.680 39.230 ;
    END
  END Q
  PIN VDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.680 38.110 14.680 39.230 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.680 24.770 14.680 25.890 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.680 11.430 14.680 12.550 ;
    END
  END clk
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.700 39.020 55.220 43.020 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.700 5.700 55.220 9.700 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 39.285 0.000 41.385 48.720 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.630 0.000 31.730 48.720 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.975 0.000 22.075 48.720 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 51.220 5.700 55.220 43.020 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.700 5.700 9.700 43.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.720 60.920 48.720 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 60.920 4.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 56.920 0.000 60.920 48.720 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.455 0.000 36.555 48.720 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.805 0.000 26.905 48.720 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 4.000 48.720 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 16.200 16.115 44.720 32.605 ;
      LAYER met1 ;
        RECT 15.810 15.960 46.030 32.760 ;
      LAYER met2 ;
        RECT 14.960 37.830 46.400 38.740 ;
        RECT 14.680 26.170 46.680 37.830 ;
        RECT 14.960 24.490 46.400 26.170 ;
        RECT 14.680 12.830 46.680 24.490 ;
        RECT 14.960 11.920 46.400 12.830 ;
      LAYER met3 ;
        RECT 19.975 16.035 41.380 32.685 ;
      LAYER met4 ;
        RECT 27.305 0.000 29.230 48.720 ;
        RECT 32.130 0.000 34.055 48.720 ;
        RECT 36.955 0.000 38.885 48.720 ;
  END
END ACMP
END LIBRARY

