* NGSPICE file created from adc_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for ACMP abstract view
.subckt ACMP INN INP Q VDD VSS clk VPWR VGND
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

.subckt adc_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12] analog_io[13]
+ analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18] analog_io[19]
+ analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23] analog_io[24]
+ analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2] analog_io[3]
+ analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ VPWR VGND
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input127_A la_data_in[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_294_ VGND VGND VPWR VPWR _294_/HI _294_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input92_A la_data_in[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput401 _109_/LO VGND VGND VPWR VPWR io_oeb[5] sky130_fd_sc_hd__clkbuf_2
Xoutput412 _154_/LO VGND VGND VPWR VPWR io_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput423 _164_/LO VGND VGND VPWR VPWR io_out[25] sky130_fd_sc_hd__clkbuf_2
Xoutput434 _340_/Q VGND VGND VPWR VPWR io_out[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput478 _182_/LO VGND VGND VPWR VPWR la_data_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput445 _267_/LO VGND VGND VPWR VPWR la_data_out[100] sky130_fd_sc_hd__clkbuf_2
Xoutput456 _277_/LO VGND VGND VPWR VPWR la_data_out[110] sky130_fd_sc_hd__clkbuf_2
Xoutput467 _287_/LO VGND VGND VPWR VPWR la_data_out[120] sky130_fd_sc_hd__clkbuf_2
Xoutput489 _192_/LO VGND VGND VPWR VPWR la_data_out[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input244_A la_oenb[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_346_ _349_/CLK _346_/D VGND VGND VPWR VPWR _346_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_277_ VGND VGND VPWR VPWR _277_/HI _277_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output463_A _284_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_200_ VGND VGND VPWR VPWR _200_/HI _200_/LO sky130_fd_sc_hd__conb_1
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_131_ VGND VGND VPWR VPWR _131_/HI _131_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input194_A la_oenb[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_062_ _062_/A VGND VGND VPWR VPWR _069_/A sky130_fd_sc_hd__buf_4
XANTENNA_input361_A wbs_dat_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input55_A la_data_in[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output580_A _312_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ VGND VGND VPWR VPWR _329_/HI _329_/LO sky130_fd_sc_hd__conb_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input207_A la_oenb[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ VGND VGND VPWR VPWR _114_/HI _114_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output426_A _166_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__080__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput301 wbs_adr_i[13] VGND VGND VPWR VPWR input301/X sky130_fd_sc_hd__buf_1
Xinput312 wbs_adr_i[23] VGND VGND VPWR VPWR input312/X sky130_fd_sc_hd__buf_1
XANTENNA_input157_A la_data_in[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput345 wbs_dat_i[23] VGND VGND VPWR VPWR input345/X sky130_fd_sc_hd__buf_1
Xinput323 wbs_adr_i[4] VGND VGND VPWR VPWR input323/X sky130_fd_sc_hd__buf_1
Xinput334 wbs_dat_i[13] VGND VGND VPWR VPWR input334/X sky130_fd_sc_hd__buf_1
XFILLER_102_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput356 wbs_dat_i[4] VGND VGND VPWR VPWR input356/X sky130_fd_sc_hd__buf_1
XANTENNA_input324_A wbs_adr_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput367 wbs_we_i VGND VGND VPWR VPWR input367/X sky130_fd_sc_hd__buf_1
XANTENNA_input18_A io_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output543_A _241_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input274_A la_oenb[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput120 la_data_in[58] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__buf_1
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput142 la_data_in[78] VGND VGND VPWR VPWR input142/X sky130_fd_sc_hd__buf_1
Xinput131 la_data_in[68] VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__buf_1
Xinput153 la_data_in[88] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__buf_1
XFILLER_64_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput164 la_data_in[98] VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_1
Xinput175 la_oenb[107] VGND VGND VPWR VPWR input175/X sky130_fd_sc_hd__buf_1
Xinput186 la_oenb[117] VGND VGND VPWR VPWR input186/X sky130_fd_sc_hd__buf_1
Xinput197 la_oenb[127] VGND VGND VPWR VPWR input197/X sky130_fd_sc_hd__buf_1
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output493_A _196_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput605 _306_/LO VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ VGND VGND VPWR VPWR _293_/HI _293_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input85_A la_data_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output506_A _207_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput402 _110_/LO VGND VGND VPWR VPWR io_oeb[6] sky130_fd_sc_hd__clkbuf_2
Xoutput413 _155_/LO VGND VGND VPWR VPWR io_out[16] sky130_fd_sc_hd__clkbuf_2
Xoutput424 _165_/LO VGND VGND VPWR VPWR io_out[26] sky130_fd_sc_hd__clkbuf_2
Xoutput435 _341_/Q VGND VGND VPWR VPWR io_out[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput446 _268_/LO VGND VGND VPWR VPWR la_data_out[101] sky130_fd_sc_hd__clkbuf_2
Xoutput457 _278_/LO VGND VGND VPWR VPWR la_data_out[111] sky130_fd_sc_hd__clkbuf_2
Xoutput468 _288_/LO VGND VGND VPWR VPWR la_data_out[121] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput479 _183_/LO VGND VGND VPWR VPWR la_data_out[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input237_A la_oenb[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_345_ _350_/CLK _345_/D VGND VGND VPWR VPWR _345_/Q sky130_fd_sc_hd__dfxtp_4
X_276_ VGND VGND VPWR VPWR _276_/HI _276_/LO sky130_fd_sc_hd__conb_1
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output456_A _277_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__050__A _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_130_ VGND VGND VPWR VPWR _130_/HI _130_/LO sky130_fd_sc_hd__conb_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_061_ _350_/Q VGND VGND VPWR VPWR _063_/A sky130_fd_sc_hd__clkinv_4
XANTENNA_input187_A la_oenb[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input354_A wbs_dat_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input48_A la_data_in[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_328_ VGND VGND VPWR VPWR _328_/HI _328_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output573_A _296_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_259_ VGND VGND VPWR VPWR _259_/HI _259_/LO sky130_fd_sc_hd__conb_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input102_A la_data_in[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ VGND VGND VPWR VPWR _113_/HI _113_/LO sky130_fd_sc_hd__conb_1
XFILLER_50_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output419_A _160_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__080__A2 _094_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput302 wbs_adr_i[14] VGND VGND VPWR VPWR input302/X sky130_fd_sc_hd__buf_1
XFILLER_102_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput324 wbs_adr_i[5] VGND VGND VPWR VPWR input324/X sky130_fd_sc_hd__buf_1
Xinput335 wbs_dat_i[14] VGND VGND VPWR VPWR input335/X sky130_fd_sc_hd__buf_1
Xinput313 wbs_adr_i[24] VGND VGND VPWR VPWR input313/X sky130_fd_sc_hd__buf_1
Xinput346 wbs_dat_i[24] VGND VGND VPWR VPWR input346/X sky130_fd_sc_hd__buf_1
Xinput357 wbs_dat_i[5] VGND VGND VPWR VPWR input357/X sky130_fd_sc_hd__buf_1
XFILLER_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input317_A wbs_adr_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output536_A _235_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__341__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__334__RESET_B hold1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input267_A la_oenb[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 la_data_in[49] VGND VGND VPWR VPWR input110/X sky130_fd_sc_hd__buf_1
XFILLER_76_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input30_A io_in[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput143 la_data_in[79] VGND VGND VPWR VPWR input143/X sky130_fd_sc_hd__buf_1
Xinput121 la_data_in[59] VGND VGND VPWR VPWR input121/X sky130_fd_sc_hd__buf_1
Xinput132 la_data_in[69] VGND VGND VPWR VPWR input132/X sky130_fd_sc_hd__buf_1
Xinput154 la_data_in[89] VGND VGND VPWR VPWR input154/X sky130_fd_sc_hd__buf_1
XFILLER_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput165 la_data_in[99] VGND VGND VPWR VPWR input165/X sky130_fd_sc_hd__buf_1
Xinput176 la_oenb[108] VGND VGND VPWR VPWR input176/X sky130_fd_sc_hd__buf_1
Xinput187 la_oenb[118] VGND VGND VPWR VPWR input187/X sky130_fd_sc_hd__buf_1
XFILLER_91_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput198 la_oenb[12] VGND VGND VPWR VPWR input198/X sky130_fd_sc_hd__buf_1
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output486_A _189_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput606 _307_/LO VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__053__A _334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_292_ VGND VGND VPWR VPWR _292_/HI _292_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input78_A la_data_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output401_A _109_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput414 _156_/LO VGND VGND VPWR VPWR io_out[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput425 _331_/X VGND VGND VPWR VPWR io_out[27] sky130_fd_sc_hd__clkbuf_2
Xoutput403 _101_/HI VGND VGND VPWR VPWR io_oeb[7] sky130_fd_sc_hd__clkbuf_2
Xoutput436 _342_/Q VGND VGND VPWR VPWR io_out[37] sky130_fd_sc_hd__clkbuf_2
Xoutput447 _269_/LO VGND VGND VPWR VPWR la_data_out[102] sky130_fd_sc_hd__clkbuf_2
Xoutput458 _279_/LO VGND VGND VPWR VPWR la_data_out[112] sky130_fd_sc_hd__clkbuf_2
Xoutput469 _289_/LO VGND VGND VPWR VPWR la_data_out[122] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input132_A la_data_in[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_344_ _350_/CLK _344_/D VGND VGND VPWR VPWR _344_/Q sky130_fd_sc_hd__dfxtp_4
X_275_ VGND VGND VPWR VPWR _275_/HI _275_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output449_A _271_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__331__A _331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__050__B _333_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_060_ _344_/Q _052_/A _343_/Q _334_/Q VGND VGND VPWR VPWR _343_/D sky130_fd_sc_hd__a22o_2
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input347_A wbs_dat_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_327_ VGND VGND VPWR VPWR _327_/HI _327_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output399_A _107_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_258_ VGND VGND VPWR VPWR _258_/HI _258_/LO sky130_fd_sc_hd__conb_1
X_189_ VGND VGND VPWR VPWR _189_/HI _189_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output566_A _262_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__B1 _335_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__061__A _350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__083__B1 _338_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input297_A wbs_adr_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_112_ VGND VGND VPWR VPWR _112_/HI _112_/LO sky130_fd_sc_hd__conb_1
XFILLER_50_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input60_A la_data_in[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__074__B1 _341_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__080__A3 _348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput303 wbs_adr_i[15] VGND VGND VPWR VPWR input303/X sky130_fd_sc_hd__buf_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput325 wbs_adr_i[6] VGND VGND VPWR VPWR input325/X sky130_fd_sc_hd__buf_1
Xinput336 wbs_dat_i[15] VGND VGND VPWR VPWR input336/X sky130_fd_sc_hd__buf_1
Xinput314 wbs_adr_i[25] VGND VGND VPWR VPWR input314/X sky130_fd_sc_hd__buf_1
Xinput347 wbs_dat_i[25] VGND VGND VPWR VPWR input347/X sky130_fd_sc_hd__buf_1
Xinput358 wbs_dat_i[6] VGND VGND VPWR VPWR input358/X sky130_fd_sc_hd__buf_1
XANTENNA__056__B1 _347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input212_A la_oenb[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output529_A _228_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output431_A _337_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input162_A la_data_in[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput100 la_data_in[3] VGND VGND VPWR VPWR input100/X sky130_fd_sc_hd__buf_1
Xinput111 la_data_in[4] VGND VGND VPWR VPWR input111/X sky130_fd_sc_hd__buf_1
XFILLER_88_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput144 la_data_in[7] VGND VGND VPWR VPWR input144/X sky130_fd_sc_hd__buf_1
Xinput122 la_data_in[5] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__buf_1
Xinput133 la_data_in[6] VGND VGND VPWR VPWR input133/X sky130_fd_sc_hd__buf_1
XFILLER_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput166 la_data_in[9] VGND VGND VPWR VPWR input166/X sky130_fd_sc_hd__buf_1
Xinput155 la_data_in[8] VGND VGND VPWR VPWR input155/X sky130_fd_sc_hd__buf_1
Xinput177 la_oenb[109] VGND VGND VPWR VPWR input177/X sky130_fd_sc_hd__buf_1
XANTENNA_input23_A io_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput199 la_oenb[13] VGND VGND VPWR VPWR input199/X sky130_fd_sc_hd__buf_1
Xinput188 la_oenb[119] VGND VGND VPWR VPWR input188/X sky130_fd_sc_hd__buf_1
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output381_A _123_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output479_A _183_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput607 _308_/LO VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_291_ VGND VGND VPWR VPWR _291_/HI _291_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output596_A _327_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput415 _157_/LO VGND VGND VPWR VPWR io_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput426 _166_/LO VGND VGND VPWR VPWR io_out[28] sky130_fd_sc_hd__clkbuf_2
Xoutput404 _102_/HI VGND VGND VPWR VPWR io_oeb[8] sky130_fd_sc_hd__clkbuf_2
Xoutput448 _270_/LO VGND VGND VPWR VPWR la_data_out[103] sky130_fd_sc_hd__clkbuf_2
Xoutput459 _280_/LO VGND VGND VPWR VPWR la_data_out[113] sky130_fd_sc_hd__clkbuf_2
Xoutput437 _142_/LO VGND VGND VPWR VPWR io_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__064__A _333_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input125_A la_data_in[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_343_ _350_/CLK _343_/D VGND VGND VPWR VPWR _343_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input90_A la_data_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_274_ VGND VGND VPWR VPWR _274_/HI _274_/LO sky130_fd_sc_hd__conb_1
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output511_A _212_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input242_A la_oenb[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_326_ VGND VGND VPWR VPWR _326_/HI _326_/LO sky130_fd_sc_hd__conb_1
XFILLER_30_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_257_ VGND VGND VPWR VPWR _257_/HI _257_/LO sky130_fd_sc_hd__conb_1
X_188_ VGND VGND VPWR VPWR _188_/HI _188_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output461_A _282_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output559_A _256_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__A1 _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__083__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_111_ VGND VGND VPWR VPWR _111_/HI _111_/LO sky130_fd_sc_hd__conb_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input192_A la_oenb[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input53_A la_data_in[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__074__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_309_ VGND VGND VPWR VPWR _309_/HI _309_/LO sky130_fd_sc_hd__conb_1
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__072__A _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput304 wbs_adr_i[16] VGND VGND VPWR VPWR input304/X sky130_fd_sc_hd__buf_1
Xinput326 wbs_adr_i[7] VGND VGND VPWR VPWR input326/X sky130_fd_sc_hd__buf_1
Xinput315 wbs_adr_i[26] VGND VGND VPWR VPWR input315/X sky130_fd_sc_hd__buf_1
Xinput348 wbs_dat_i[26] VGND VGND VPWR VPWR input348/X sky130_fd_sc_hd__buf_1
Xinput359 wbs_dat_i[7] VGND VGND VPWR VPWR input359/X sky130_fd_sc_hd__buf_1
Xinput337 wbs_dat_i[16] VGND VGND VPWR VPWR input337/X sky130_fd_sc_hd__buf_1
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__056__A1 _348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__056__B2 _053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input205_A la_oenb[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output424_A _165_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput101 la_data_in[40] VGND VGND VPWR VPWR input101/X sky130_fd_sc_hd__buf_1
XANTENNA_input155_A la_data_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput145 la_data_in[80] VGND VGND VPWR VPWR input145/X sky130_fd_sc_hd__buf_1
Xinput134 la_data_in[70] VGND VGND VPWR VPWR input134/X sky130_fd_sc_hd__buf_1
Xinput123 la_data_in[60] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__buf_1
Xinput112 la_data_in[50] VGND VGND VPWR VPWR input112/X sky130_fd_sc_hd__buf_1
Xinput178 la_oenb[10] VGND VGND VPWR VPWR input178/X sky130_fd_sc_hd__buf_1
Xinput167 la_oenb[0] VGND VGND VPWR VPWR input167/X sky130_fd_sc_hd__buf_1
XANTENNA_input322_A wbs_adr_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput156 la_data_in[90] VGND VGND VPWR VPWR input156/X sky130_fd_sc_hd__buf_1
XFILLER_48_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input16_A io_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput189 la_oenb[11] VGND VGND VPWR VPWR input189/X sky130_fd_sc_hd__buf_1
XFILLER_56_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output374_A _117_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output541_A _239_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input8_A io_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_290_ VGND VGND VPWR VPWR _290_/HI _290_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input272_A la_oenb[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output491_A _194_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output589_A _320_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput416 _158_/LO VGND VGND VPWR VPWR io_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput405 _111_/LO VGND VGND VPWR VPWR io_oeb[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput449 _271_/LO VGND VGND VPWR VPWR la_data_out[104] sky130_fd_sc_hd__clkbuf_2
Xoutput438 _143_/LO VGND VGND VPWR VPWR io_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput427 _332_/X VGND VGND VPWR VPWR io_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input118_A la_data_in[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_342_ _350_/CLK _342_/D VGND VGND VPWR VPWR _342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_273_ VGND VGND VPWR VPWR _273_/HI _273_/LO sky130_fd_sc_hd__conb_1
XFILLER_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input83_A la_data_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output504_A _206_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input235_A la_oenb[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_325_ VGND VGND VPWR VPWR _325_/HI _325_/LO sky130_fd_sc_hd__conb_1
X_256_ VGND VGND VPWR VPWR _256_/HI _256_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_187_ VGND VGND VPWR VPWR _187_/HI _187_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output454_A _276_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__A2 _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__344__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__083__A2 _094_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_110_ VGND VGND VPWR VPWR _110_/HI _110_/LO sky130_fd_sc_hd__conb_1
XFILLER_8_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input185_A la_oenb[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input352_A wbs_dat_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input46_A la_data_in[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__074__A2 _094_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output571_A _176_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ VGND VGND VPWR VPWR _308_/HI _308_/LO sky130_fd_sc_hd__conb_1
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_239_ VGND VGND VPWR VPWR _239_/HI _239_/LO sky130_fd_sc_hd__conb_1
XFILLER_115_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput316 wbs_adr_i[27] VGND VGND VPWR VPWR input316/X sky130_fd_sc_hd__buf_1
Xinput327 wbs_adr_i[8] VGND VGND VPWR VPWR input327/X sky130_fd_sc_hd__buf_1
Xinput305 wbs_adr_i[17] VGND VGND VPWR VPWR input305/X sky130_fd_sc_hd__buf_1
XFILLER_48_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput349 wbs_dat_i[27] VGND VGND VPWR VPWR input349/X sky130_fd_sc_hd__buf_1
Xinput338 wbs_dat_i[17] VGND VGND VPWR VPWR input338/X sky130_fd_sc_hd__buf_1
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__056__A2 _052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input100_A la_data_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output417_A _140_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput102 la_data_in[41] VGND VGND VPWR VPWR input102/X sky130_fd_sc_hd__buf_1
XFILLER_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput113 la_data_in[51] VGND VGND VPWR VPWR input113/X sky130_fd_sc_hd__buf_1
Xinput124 la_data_in[61] VGND VGND VPWR VPWR input124/X sky130_fd_sc_hd__buf_1
Xinput135 la_data_in[71] VGND VGND VPWR VPWR input135/X sky130_fd_sc_hd__buf_1
XANTENNA_input148_A la_data_in[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput146 la_data_in[81] VGND VGND VPWR VPWR input146/X sky130_fd_sc_hd__buf_1
Xinput168 la_oenb[100] VGND VGND VPWR VPWR input168/X sky130_fd_sc_hd__buf_1
Xinput157 la_data_in[91] VGND VGND VPWR VPWR input157/X sky130_fd_sc_hd__buf_1
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput179 la_oenb[110] VGND VGND VPWR VPWR input179/X sky130_fd_sc_hd__buf_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input315_A wbs_adr_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output534_A _233_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input265_A la_oenb[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output484_A _187_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput406 _139_/LO VGND VGND VPWR VPWR io_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput417 _140_/LO VGND VGND VPWR VPWR io_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput428 _141_/LO VGND VGND VPWR VPWR io_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput439 _144_/LO VGND VGND VPWR VPWR io_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_341_ _350_/CLK _341_/D VGND VGND VPWR VPWR _341_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_272_ VGND VGND VPWR VPWR _272_/HI _272_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input76_A la_data_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__091__A _343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__086__B1 _337_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input130_A la_data_in[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input228_A la_oenb[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_324_ VGND VGND VPWR VPWR _324_/HI _324_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_255_ VGND VGND VPWR VPWR _255_/HI _255_/LO sky130_fd_sc_hd__conb_1
X_186_ VGND VGND VPWR VPWR _186_/HI _186_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output447_A _269_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__077__B1 _340_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__092__A3 _344_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__083__A3 _347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input178_A la_oenb[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input345_A wbs_dat_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__059__B1 _344_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input39_A la_data_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__074__A3 _350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output397_A _137_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_307_ VGND VGND VPWR VPWR _307_/HI _307_/LO sky130_fd_sc_hd__conb_1
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_238_ VGND VGND VPWR VPWR _238_/HI _238_/LO sky130_fd_sc_hd__conb_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_169_ VGND VGND VPWR VPWR _169_/HI _169_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output564_A _260_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput317 wbs_adr_i[28] VGND VGND VPWR VPWR input317/X sky130_fd_sc_hd__buf_1
Xinput306 wbs_adr_i[18] VGND VGND VPWR VPWR input306/X sky130_fd_sc_hd__buf_1
Xinput328 wbs_adr_i[9] VGND VGND VPWR VPWR input328/X sky130_fd_sc_hd__buf_1
Xinput339 wbs_dat_i[18] VGND VGND VPWR VPWR input339/X sky130_fd_sc_hd__buf_1
XFILLER_56_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input295_A user_clock2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__334__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput136 la_data_in[72] VGND VGND VPWR VPWR input136/X sky130_fd_sc_hd__buf_1
Xinput125 la_data_in[62] VGND VGND VPWR VPWR input125/X sky130_fd_sc_hd__buf_1
Xinput114 la_data_in[52] VGND VGND VPWR VPWR input114/X sky130_fd_sc_hd__buf_1
Xinput103 la_data_in[42] VGND VGND VPWR VPWR input103/X sky130_fd_sc_hd__buf_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput147 la_data_in[82] VGND VGND VPWR VPWR input147/X sky130_fd_sc_hd__buf_1
Xinput158 la_data_in[92] VGND VGND VPWR VPWR input158/X sky130_fd_sc_hd__buf_1
Xinput169 la_oenb[101] VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__buf_1
XFILLER_56_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input210_A la_oenb[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input308_A wbs_adr_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output527_A _172_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__334__D _334_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__094__A _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input258_A la_oenb[67] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input160_A la_data_in[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input21_A io_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output477_A _181_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput407 _149_/LO VGND VGND VPWR VPWR io_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput418 _159_/LO VGND VGND VPWR VPWR io_out[20] sky130_fd_sc_hd__clkbuf_2
Xoutput429 _335_/Q VGND VGND VPWR VPWR io_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_340_ _350_/CLK _340_/D VGND VGND VPWR VPWR _340_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_271_ VGND VGND VPWR VPWR _271_/HI _271_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input69_A la_data_in[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__086__A1 _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input123_A la_data_in[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_323_ VGND VGND VPWR VPWR _323_/HI _323_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_254_ VGND VGND VPWR VPWR _254_/HI _254_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_185_ VGND VGND VPWR VPWR _185_/HI _185_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__077__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output607_A _308_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__342__D _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput590 _321_/LO VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__clkbuf_2
XANTENNA__059__B2 _334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__059__A1 _345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input338_A wbs_dat_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input240_A la_oenb[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_306_ VGND VGND VPWR VPWR _306_/HI _306_/LO sky130_fd_sc_hd__conb_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_237_ VGND VGND VPWR VPWR _237_/HI _237_/LO sky130_fd_sc_hd__conb_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_168_ VGND VGND VPWR VPWR _168_/HI _168_/LO sky130_fd_sc_hd__conb_1
XFILLER_115_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output557_A _254_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ _099_/A _099_/B VGND VGND VPWR VPWR _334_/D sky130_fd_sc_hd__nor2_8
XFILLER_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__337__D _337_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput307 wbs_adr_i[19] VGND VGND VPWR VPWR input307/X sky130_fd_sc_hd__buf_1
Xinput318 wbs_adr_i[29] VGND VGND VPWR VPWR input318/X sky130_fd_sc_hd__buf_1
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput329 wbs_cyc_i VGND VGND VPWR VPWR input329/X sky130_fd_sc_hd__buf_1
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__097__A _346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input190_A la_oenb[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input288_A la_oenb[94] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input51_A la_data_in[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput104 la_data_in[43] VGND VGND VPWR VPWR input104/X sky130_fd_sc_hd__buf_1
Xinput126 la_data_in[63] VGND VGND VPWR VPWR input126/X sky130_fd_sc_hd__buf_1
Xinput115 la_data_in[53] VGND VGND VPWR VPWR input115/X sky130_fd_sc_hd__buf_1
Xinput148 la_data_in[83] VGND VGND VPWR VPWR input148/X sky130_fd_sc_hd__buf_1
Xinput137 la_data_in[73] VGND VGND VPWR VPWR input137/X sky130_fd_sc_hd__buf_1
Xinput159 la_data_in[93] VGND VGND VPWR VPWR input159/X sky130_fd_sc_hd__buf_1
XFILLER_17_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input203_A la_oenb[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A la_data_in[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output422_A _163_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__350__D _350_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__094__B _094_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input153_A la_data_in[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input320_A wbs_adr_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input14_A io_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output372_A _115_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput408 _150_/LO VGND VGND VPWR VPWR io_out[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput419 _160_/LO VGND VGND VPWR VPWR io_out[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__347__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__345__D _345_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input6_A io_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ VGND VGND VPWR VPWR _270_/HI _270_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input270_A la_oenb[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output587_A _300_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__086__A2 _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input116_A la_data_in[54] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_322_ VGND VGND VPWR VPWR _322_/HI _322_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_253_ VGND VGND VPWR VPWR _253_/HI _253_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input81_A la_data_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_184_ VGND VGND VPWR VPWR _184_/HI _184_/LO sky130_fd_sc_hd__conb_1
XFILLER_108_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__077__A2 _094_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output502_A _204_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput580 _312_/LO VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__clkbuf_2
XANTENNA__059__A2 _052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput591 _322_/LO VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input233_A la_oenb[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305_ VGND VGND VPWR VPWR _305_/HI _305_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_236_ VGND VGND VPWR VPWR _236_/HI _236_/LO sky130_fd_sc_hd__conb_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_167_ VGND VGND VPWR VPWR _167_/HI _167_/LO sky130_fd_sc_hd__conb_1
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_098_ _052_/X _099_/B _098_/B1 _066_/Y VGND VGND VPWR VPWR _333_/D sky130_fd_sc_hd__a22o_2
XANTENNA_output452_A _274_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput308 wbs_adr_i[1] VGND VGND VPWR VPWR input308/X sky130_fd_sc_hd__buf_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput319 wbs_adr_i[2] VGND VGND VPWR VPWR input319/X sky130_fd_sc_hd__buf_1
XFILLER_96_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__097__B _345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input183_A la_oenb[114] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input350_A wbs_dat_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input44_A la_data_in[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_219_ VGND VGND VPWR VPWR _219_/HI _219_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__348__D _348_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput116 la_data_in[54] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__buf_1
Xinput127 la_data_in[64] VGND VGND VPWR VPWR input127/X sky130_fd_sc_hd__buf_1
Xinput105 la_data_in[44] VGND VGND VPWR VPWR input105/X sky130_fd_sc_hd__buf_1
XFILLER_49_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput138 la_data_in[74] VGND VGND VPWR VPWR input138/X sky130_fd_sc_hd__buf_1
Xinput149 la_data_in[84] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__buf_1
XFILLER_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output415_A _157_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input146_A la_data_in[81] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input313_A wbs_adr_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput409 _151_/LO VGND VGND VPWR VPWR io_out[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_79_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _350_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__098__B1 _098_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input263_A la_oenb[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__089__B1 _336_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output482_A _186_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__086__A3 _346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_321_ VGND VGND VPWR VPWR _321_/HI _321_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input109_A la_data_in[48] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_252_ VGND VGND VPWR VPWR _252_/HI _252_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_183_ VGND VGND VPWR VPWR _183_/HI _183_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input74_A la_data_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__337__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__077__A3 _349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput581 _313_/LO VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput570 _266_/LO VGND VGND VPWR VPWR la_data_out[99] sky130_fd_sc_hd__clkbuf_2
Xoutput592 _323_/LO VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input226_A la_oenb[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_304_ VGND VGND VPWR VPWR _304_/HI _304_/LO sky130_fd_sc_hd__conb_1
X_235_ VGND VGND VPWR VPWR _235_/HI _235_/LO sky130_fd_sc_hd__conb_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_166_ VGND VGND VPWR VPWR _166_/HI _166_/LO sky130_fd_sc_hd__conb_1
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_097_ _346_/Q _345_/Q _097_/C _097_/D VGND VGND VPWR VPWR _099_/B sky130_fd_sc_hd__or4_4
XFILLER_97_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output445_A _267_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput309 wbs_adr_i[20] VGND VGND VPWR VPWR input309/X sky130_fd_sc_hd__buf_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__097__C _097_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input176_A la_oenb[108] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input343_A wbs_dat_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input37_A io_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output395_A _135_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_218_ VGND VGND VPWR VPWR _218_/HI _218_/LO sky130_fd_sc_hd__conb_1
X_149_ VGND VGND VPWR VPWR _149_/HI _149_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output562_A _258_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput106 la_data_in[45] VGND VGND VPWR VPWR input106/X sky130_fd_sc_hd__buf_1
Xinput117 la_data_in[55] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__buf_1
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput128 la_data_in[65] VGND VGND VPWR VPWR input128/X sky130_fd_sc_hd__buf_1
Xinput139 la_data_in[75] VGND VGND VPWR VPWR input139/X sky130_fd_sc_hd__buf_1
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input293_A la_oenb[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output408_A _150_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input139_A la_data_in[75] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input306_A wbs_adr_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output525_A _225_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__098__B2 _066_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__098__A1 _052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__089__A1 _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input256_A la_oenb[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output475_A _179_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_320_ VGND VGND VPWR VPWR _320_/HI _320_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_251_ VGND VGND VPWR VPWR _251_/HI _251_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_182_ VGND VGND VPWR VPWR _182_/HI _182_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input67_A la_data_in[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output592_A _323_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput571 _176_/LO VGND VGND VPWR VPWR la_data_out[9] sky130_fd_sc_hd__clkbuf_2
Xoutput560 _175_/LO VGND VGND VPWR VPWR la_data_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput582 _314_/LO VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput593 _324_/LO VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input121_A la_data_in[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input219_A la_oenb[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_303_ VGND VGND VPWR VPWR _303_/HI _303_/LO sky130_fd_sc_hd__conb_1
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_234_ VGND VGND VPWR VPWR _234_/HI _234_/LO sky130_fd_sc_hd__conb_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_165_ VGND VGND VPWR VPWR _165_/HI _165_/LO sky130_fd_sc_hd__conb_1
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_096_ _350_/Q _349_/Q _348_/Q _347_/Q VGND VGND VPWR VPWR _097_/D sky130_fd_sc_hd__or4_4
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output438_A _143_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output605_A _306_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__097__D _097_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input169_A la_oenb[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput390 _106_/LO VGND VGND VPWR VPWR io_oeb[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input336_A wbs_dat_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_217_ VGND VGND VPWR VPWR _217_/HI _217_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output388_A _103_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_148_ VGND VGND VPWR VPWR _148_/HI _148_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output555_A _252_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ _347_/Q VGND VGND VPWR VPWR _079_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput107 la_data_in[46] VGND VGND VPWR VPWR input107/X sky130_fd_sc_hd__buf_1
Xinput118 la_data_in[56] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__buf_1
XFILLER_102_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput129 la_data_in[66] VGND VGND VPWR VPWR input129/X sky130_fd_sc_hd__buf_1
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input286_A la_oenb[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input201_A la_oenb[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input97_A la_data_in[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output420_A _161_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output518_A _218_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__098__A2 _099_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__089__A2 _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input151_A la_data_in[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input249_A la_oenb[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input12_A io_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output370_A _113_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output468_A _288_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput290 la_oenb[96] VGND VGND VPWR VPWR input290/X sky130_fd_sc_hd__buf_1
XFILLER_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input4_A io_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ VGND VGND VPWR VPWR _250_/HI _250_/LO sky130_fd_sc_hd__conb_1
X_181_ VGND VGND VPWR VPWR _181_/HI _181_/LO sky130_fd_sc_hd__conb_1
XFILLER_50_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input199_A la_oenb[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input366_A wbs_stb_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output585_A _317_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput550 _247_/LO VGND VGND VPWR VPWR la_data_out[80] sky130_fd_sc_hd__clkbuf_2
Xoutput561 _257_/LO VGND VGND VPWR VPWR la_data_out[90] sky130_fd_sc_hd__clkbuf_2
Xoutput572 _295_/LO VGND VGND VPWR VPWR user_irq[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput583 _315_/LO VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__clkbuf_2
Xoutput594 _325_/LO VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input114_A la_data_in[52] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_302_ VGND VGND VPWR VPWR _302_/HI _302_/LO sky130_fd_sc_hd__conb_1
X_233_ VGND VGND VPWR VPWR _233_/HI _233_/LO sky130_fd_sc_hd__conb_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_164_ VGND VGND VPWR VPWR _164_/HI _164_/LO sky130_fd_sc_hd__conb_1
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_095_ _344_/Q _095_/B VGND VGND VPWR VPWR _097_/C sky130_fd_sc_hd__or2_2
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output500_A _202_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput380 _122_/LO VGND VGND VPWR VPWR io_oeb[20] sky130_fd_sc_hd__clkbuf_2
Xoutput391 _131_/LO VGND VGND VPWR VPWR io_oeb[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input231_A la_oenb[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input329_A wbs_cyc_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ VGND VGND VPWR VPWR _216_/HI _216_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_147_ VGND VGND VPWR VPWR _147_/HI _147_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output548_A _246_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output450_A _272_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ _076_/Y _099_/A _070_/X _071_/X _077_/X VGND VGND VPWR VPWR _340_/D sky130_fd_sc_hd__o311a_1
XFILLER_112_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput108 la_data_in[47] VGND VGND VPWR VPWR input108/X sky130_fd_sc_hd__buf_1
XFILLER_102_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput119 la_data_in[57] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__buf_1
XFILLER_69_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input279_A la_oenb[86] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input181_A la_oenb[112] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input42_A la_data_in[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output498_A _200_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput90 la_data_in[30] VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__buf_1
XFILLER_103_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output413_A _155_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__089__A3 _345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input144_A la_data_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input311_A wbs_adr_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output530_A _229_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput280 la_oenb[87] VGND VGND VPWR VPWR input280/X sky130_fd_sc_hd__buf_1
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput291 la_oenb[97] VGND VGND VPWR VPWR input291/X sky130_fd_sc_hd__buf_1
XFILLER_48_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_180_ VGND VGND VPWR VPWR _180_/HI _180_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input261_A la_oenb[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input359_A wbs_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _349_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output480_A _184_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output578_A _310_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput551 _248_/LO VGND VGND VPWR VPWR la_data_out[81] sky130_fd_sc_hd__clkbuf_2
Xoutput540 _238_/LO VGND VGND VPWR VPWR la_data_out[71] sky130_fd_sc_hd__clkbuf_2
Xoutput562 _258_/LO VGND VGND VPWR VPWR la_data_out[91] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput584 _316_/LO VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__clkbuf_2
Xoutput595 _326_/LO VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput573 _296_/LO VGND VGND VPWR VPWR user_irq[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input107_A la_data_in[46] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_301_ VGND VGND VPWR VPWR _301_/HI _301_/LO sky130_fd_sc_hd__conb_1
X_232_ VGND VGND VPWR VPWR _232_/HI _232_/LO sky130_fd_sc_hd__conb_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_163_ VGND VGND VPWR VPWR _163_/HI _163_/LO sky130_fd_sc_hd__conb_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input72_A la_data_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_094_ _094_/A _094_/B VGND VGND VPWR VPWR _332_/A sky130_fd_sc_hd__nor2_1
XFILLER_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__350__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput370 _113_/LO VGND VGND VPWR VPWR io_oeb[11] sky130_fd_sc_hd__clkbuf_2
Xoutput381 _123_/LO VGND VGND VPWR VPWR io_oeb[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput392 _132_/LO VGND VGND VPWR VPWR io_oeb[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input224_A la_oenb[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ VGND VGND VPWR VPWR _215_/HI _215_/LO sky130_fd_sc_hd__conb_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_146_ VGND VGND VPWR VPWR _146_/HI _146_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_077_ _094_/A _094_/B _349_/Q _340_/Q VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__a31o_2
XANTENNA_output443_A _148_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput109 la_data_in[48] VGND VGND VPWR VPWR input109/X sky130_fd_sc_hd__buf_1
XFILLER_69_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input174_A la_oenb[106] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input341_A wbs_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input35_A io_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output393_A _133_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output560_A _175_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_129_ VGND VGND VPWR VPWR _129_/HI _129_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput80 la_data_in[21] VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_1
Xinput91 la_data_in[31] VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__buf_1
XFILLER_89_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input291_A la_oenb[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output406_A _139_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input137_A la_data_in[73] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input304_A wbs_adr_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output523_A _223_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput270 la_oenb[78] VGND VGND VPWR VPWR input270/X sky130_fd_sc_hd__buf_1
Xinput281 la_oenb[88] VGND VGND VPWR VPWR input281/X sky130_fd_sc_hd__buf_1
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput292 la_oenb[98] VGND VGND VPWR VPWR input292/X sky130_fd_sc_hd__buf_1
XFILLER_48_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input254_A la_oenb[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output473_A _293_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput530 _229_/LO VGND VGND VPWR VPWR la_data_out[62] sky130_fd_sc_hd__clkbuf_2
Xoutput552 _249_/LO VGND VGND VPWR VPWR la_data_out[82] sky130_fd_sc_hd__clkbuf_2
Xoutput541 _239_/LO VGND VGND VPWR VPWR la_data_out[72] sky130_fd_sc_hd__clkbuf_2
Xoutput563 _259_/LO VGND VGND VPWR VPWR la_data_out[92] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput596 _327_/LO VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput585 _317_/LO VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput574 _297_/LO VGND VGND VPWR VPWR user_irq[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_300_ VGND VGND VPWR VPWR _300_/HI _300_/LO sky130_fd_sc_hd__conb_1
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_231_ VGND VGND VPWR VPWR _231_/HI _231_/LO sky130_fd_sc_hd__conb_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_162_ VGND VGND VPWR VPWR _162_/HI _162_/LO sky130_fd_sc_hd__conb_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_093_ _095_/B _331_/A _099_/A _071_/A _092_/X VGND VGND VPWR VPWR _335_/D sky130_fd_sc_hd__o311a_4
XANTENNA_input65_A la_data_in[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__333__RESET_B hold1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output590_A _321_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput1 io_in[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_1
XFILLER_37_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput371 _114_/LO VGND VGND VPWR VPWR io_oeb[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput382 _124_/LO VGND VGND VPWR VPWR io_oeb[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput393 _133_/LO VGND VGND VPWR VPWR io_oeb[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input217_A la_oenb[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ VGND VGND VPWR VPWR _214_/HI _214_/LO sky130_fd_sc_hd__conb_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_145_ VGND VGND VPWR VPWR _145_/HI _145_/LO sky130_fd_sc_hd__conb_1
X_076_ _348_/Q VGND VGND VPWR VPWR _076_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output436_A _342_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output603_A _304_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__340__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input167_A la_oenb[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input334_A wbs_dat_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input28_A io_in[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output386_A _128_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_128_ VGND VGND VPWR VPWR _128_/HI _128_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output553_A _250_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_059_ _345_/Q _052_/A _344_/Q _334_/Q VGND VGND VPWR VPWR _344_/D sky130_fd_sc_hd__a22o_1
XFILLER_98_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput81 la_data_in[22] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_1
Xinput70 la_data_in[12] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__buf_1
XFILLER_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput92 la_data_in[32] VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__buf_1
XFILLER_103_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input284_A la_oenb[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input95_A la_data_in[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output516_A _171_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput260 la_oenb[69] VGND VGND VPWR VPWR input260/X sky130_fd_sc_hd__buf_1
Xinput271 la_oenb[79] VGND VGND VPWR VPWR input271/X sky130_fd_sc_hd__buf_1
XFILLER_63_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput293 la_oenb[99] VGND VGND VPWR VPWR input293/X sky130_fd_sc_hd__buf_1
Xinput282 la_oenb[89] VGND VGND VPWR VPWR input282/X sky130_fd_sc_hd__buf_1
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input247_A la_oenb[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input10_A io_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output466_A _178_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput520 _220_/LO VGND VGND VPWR VPWR la_data_out[53] sky130_fd_sc_hd__clkbuf_2
Xoutput542 _240_/LO VGND VGND VPWR VPWR la_data_out[73] sky130_fd_sc_hd__clkbuf_2
Xoutput531 _230_/LO VGND VGND VPWR VPWR la_data_out[63] sky130_fd_sc_hd__clkbuf_2
Xoutput553 _250_/LO VGND VGND VPWR VPWR la_data_out[83] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput586 _318_/LO VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput575 _298_/LO VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__clkbuf_2
Xoutput564 _260_/LO VGND VGND VPWR VPWR la_data_out[93] sky130_fd_sc_hd__clkbuf_2
XANTENNA__051__A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput597 _328_/LO VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A io_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_230_ VGND VGND VPWR VPWR _230_/HI _230_/LO sky130_fd_sc_hd__conb_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_161_ VGND VGND VPWR VPWR _161_/HI _161_/LO sky130_fd_sc_hd__conb_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input197_A la_oenb[127] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_092_ _072_/A _073_/A _344_/Q _335_/Q VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__a31o_2
XFILLER_40_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input364_A wbs_sel_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_A la_data_in[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output583_A _315_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 io_in[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_1
XFILLER_110_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput372 _115_/LO VGND VGND VPWR VPWR io_oeb[13] sky130_fd_sc_hd__clkbuf_2
Xoutput383 _125_/LO VGND VGND VPWR VPWR io_oeb[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput394 _134_/LO VGND VGND VPWR VPWR io_oeb[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__055__B1 _348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input112_A la_data_in[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_213_ VGND VGND VPWR VPWR _213_/HI _213_/LO sky130_fd_sc_hd__conb_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_144_ VGND VGND VPWR VPWR _144_/HI _144_/LO sky130_fd_sc_hd__conb_1
X_075_ _068_/Y _099_/A _070_/X _071_/X _074_/X VGND VGND VPWR VPWR _341_/D sky130_fd_sc_hd__o311a_2
XFILLER_111_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output429_A _335_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input327_A wbs_adr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output379_A _105_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_127_ VGND VGND VPWR VPWR _127_/HI _127_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output546_A _244_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_058_ _346_/Q _052_/A _345_/Q _053_/X VGND VGND VPWR VPWR _345_/D sky130_fd_sc_hd__a22o_2
XFILLER_98_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput82 la_data_in[23] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_1
Xinput71 la_data_in[13] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_1
Xinput60 la_data_in[119] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_1
XFILLER_115_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput93 la_data_in[33] VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_1
XFILLER_89_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input277_A la_oenb[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A la_data_in[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output496_A _198_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input88_A la_data_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput261 la_oenb[6] VGND VGND VPWR VPWR input261/X sky130_fd_sc_hd__buf_1
Xinput250 la_oenb[5] VGND VGND VPWR VPWR input250/X sky130_fd_sc_hd__buf_1
Xinput272 la_oenb[7] VGND VGND VPWR VPWR input272/X sky130_fd_sc_hd__buf_1
XANTENNA_output411_A _153_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput294 la_oenb[9] VGND VGND VPWR VPWR input294/X sky130_fd_sc_hd__buf_1
Xinput283 la_oenb[8] VGND VGND VPWR VPWR input283/X sky130_fd_sc_hd__buf_1
XANTENNA_output509_A _210_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__049__A _334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input142_A la_data_in[78] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output459_A _280_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput510 _211_/LO VGND VGND VPWR VPWR la_data_out[44] sky130_fd_sc_hd__clkbuf_2
Xoutput543 _241_/LO VGND VGND VPWR VPWR la_data_out[74] sky130_fd_sc_hd__clkbuf_2
Xoutput521 _221_/LO VGND VGND VPWR VPWR la_data_out[54] sky130_fd_sc_hd__clkbuf_2
Xoutput532 _231_/LO VGND VGND VPWR VPWR la_data_out[64] sky130_fd_sc_hd__clkbuf_2
Xoutput554 _251_/LO VGND VGND VPWR VPWR la_data_out[84] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput587 _300_/LO VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput576 _299_/LO VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput565 _261_/LO VGND VGND VPWR VPWR la_data_out[94] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput598 _301_/LO VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_160_ VGND VGND VPWR VPWR _160_/HI _160_/LO sky130_fd_sc_hd__conb_1
XFILLER_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ _343_/Q VGND VGND VPWR VPWR _095_/B sky130_fd_sc_hd__clkinv_4
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input357_A wbs_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output576_A _299_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ VGND VGND VPWR VPWR _289_/HI _289_/LO sky130_fd_sc_hd__conb_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput3 io_in[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_1
XFILLER_49_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__062__A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput373 _116_/LO VGND VGND VPWR VPWR io_oeb[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput384 _126_/LO VGND VGND VPWR VPWR io_oeb[24] sky130_fd_sc_hd__clkbuf_2
Xoutput395 _135_/LO VGND VGND VPWR VPWR io_oeb[34] sky130_fd_sc_hd__clkbuf_2
XANTENNA__055__A1 _349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__055__B2 _053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A la_data_in[44] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ VGND VGND VPWR VPWR _212_/HI _212_/LO sky130_fd_sc_hd__conb_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_143_ VGND VGND VPWR VPWR _143_/HI _143_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input70_A la_data_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ _094_/A _094_/B _350_/Q _341_/Q VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__a31o_2
XFILLER_3_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input222_A la_oenb[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_126_ VGND VGND VPWR VPWR _126_/HI _126_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_057_ _347_/Q _052_/A _346_/Q _053_/X VGND VGND VPWR VPWR _346_/D sky130_fd_sc_hd__a22o_2
XFILLER_97_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output539_A _237_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput72 la_data_in[14] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__buf_1
Xinput61 la_data_in[11] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_1
Xinput50 la_data_in[10] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_1
Xinput83 la_data_in[24] VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_1
Xinput94 la_data_in[34] VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__buf_1
XFILLER_115_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input172_A la_oenb[104] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input33_A io_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output489_A _192_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output391_A _131_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_109_ VGND VGND VPWR VPWR _109_/HI _109_/LO sky130_fd_sc_hd__conb_1
XFILLER_112_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__070__A _331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__100__B1 _071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput262 la_oenb[70] VGND VGND VPWR VPWR input262/X sky130_fd_sc_hd__buf_1
Xinput240 la_oenb[50] VGND VGND VPWR VPWR input240/X sky130_fd_sc_hd__buf_1
Xinput251 la_oenb[60] VGND VGND VPWR VPWR input251/X sky130_fd_sc_hd__buf_1
XFILLER_76_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput273 la_oenb[80] VGND VGND VPWR VPWR input273/X sky130_fd_sc_hd__buf_1
Xinput284 la_oenb[90] VGND VGND VPWR VPWR input284/X sky130_fd_sc_hd__buf_1
Xinput295 user_clock2 VGND VGND VPWR VPWR input295/X sky130_fd_sc_hd__buf_1
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__065__A _334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input135_A la_data_in[71] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input302_A wbs_adr_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output521_A _221_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput511 _212_/LO VGND VGND VPWR VPWR la_data_out[45] sky130_fd_sc_hd__clkbuf_2
Xoutput500 _202_/LO VGND VGND VPWR VPWR la_data_out[35] sky130_fd_sc_hd__clkbuf_2
Xoutput533 _232_/LO VGND VGND VPWR VPWR la_data_out[65] sky130_fd_sc_hd__clkbuf_2
Xoutput522 _222_/LO VGND VGND VPWR VPWR la_data_out[55] sky130_fd_sc_hd__clkbuf_2
Xoutput544 _242_/LO VGND VGND VPWR VPWR la_data_out[75] sky130_fd_sc_hd__clkbuf_2
Xoutput577 _309_/LO VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput555 _252_/LO VGND VGND VPWR VPWR la_data_out[85] sky130_fd_sc_hd__clkbuf_2
Xoutput566 _262_/LO VGND VGND VPWR VPWR la_data_out[95] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput599 _329_/LO VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__clkbuf_2
Xoutput588 _319_/LO VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_74_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_090_ _088_/Y _069_/A _331_/A _071_/A _089_/X VGND VGND VPWR VPWR _336_/D sky130_fd_sc_hd__o311a_2
XANTENNA__343__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input252_A la_oenb[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_288_ VGND VGND VPWR VPWR _288_/HI _288_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output569_A _265_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output471_A _291_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput4 io_in[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
XFILLER_49_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput374 _117_/LO VGND VGND VPWR VPWR io_oeb[15] sky130_fd_sc_hd__clkbuf_2
Xoutput385 _127_/LO VGND VGND VPWR VPWR io_oeb[25] sky130_fd_sc_hd__clkbuf_2
Xoutput396 _136_/LO VGND VGND VPWR VPWR io_oeb[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__055__A2 _052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ VGND VGND VPWR VPWR _211_/HI _211_/LO sky130_fd_sc_hd__conb_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_142_ VGND VGND VPWR VPWR _142_/HI _142_/LO sky130_fd_sc_hd__conb_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_073_ _073_/A VGND VGND VPWR VPWR _094_/B sky130_fd_sc_hd__buf_8
XANTENNA_input63_A la_data_in[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__073__A _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input215_A la_oenb[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_125_ VGND VGND VPWR VPWR _125_/HI _125_/LO sky130_fd_sc_hd__conb_1
X_056_ _348_/Q _052_/X _347_/Q _053_/X VGND VGND VPWR VPWR _347_/D sky130_fd_sc_hd__a22o_2
XFILLER_3_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output434_A _340_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output601_A _302_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput40 la_data_in[100] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__buf_1
Xinput73 la_data_in[15] VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__buf_1
Xinput51 la_data_in[110] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_1
Xinput62 la_data_in[120] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_1
Xinput84 la_data_in[25] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_1
Xinput95 la_data_in[35] VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__buf_1
XFILLER_115_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__068__A _349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input165_A la_data_in[99] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input332_A wbs_dat_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input26_A io_in[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output384_A _126_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ VGND VGND VPWR VPWR _108_/HI _108_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output551_A _248_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__100__A1 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input282_A la_oenb[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput230 la_oenb[41] VGND VGND VPWR VPWR input230/X sky130_fd_sc_hd__buf_1
Xinput263 la_oenb[71] VGND VGND VPWR VPWR input263/X sky130_fd_sc_hd__buf_1
Xinput252 la_oenb[61] VGND VGND VPWR VPWR input252/X sky130_fd_sc_hd__buf_1
Xinput241 la_oenb[51] VGND VGND VPWR VPWR input241/X sky130_fd_sc_hd__buf_1
Xinput296 wb_rst_i VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__buf_6
Xinput274 la_oenb[81] VGND VGND VPWR VPWR input274/X sky130_fd_sc_hd__buf_1
Xinput285 la_oenb[91] VGND VGND VPWR VPWR input285/X sky130_fd_sc_hd__buf_1
XFILLER_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output599_A _329_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__065__B _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input128_A la_data_in[65] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input93_A la_data_in[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output514_A _215_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput501 _203_/LO VGND VGND VPWR VPWR la_data_out[36] sky130_fd_sc_hd__clkbuf_2
Xoutput512 _213_/LO VGND VGND VPWR VPWR la_data_out[46] sky130_fd_sc_hd__clkbuf_2
Xoutput545 _243_/LO VGND VGND VPWR VPWR la_data_out[76] sky130_fd_sc_hd__clkbuf_2
Xoutput534 _233_/LO VGND VGND VPWR VPWR la_data_out[66] sky130_fd_sc_hd__clkbuf_2
Xoutput523 _223_/LO VGND VGND VPWR VPWR la_data_out[56] sky130_fd_sc_hd__clkbuf_2
Xoutput578 _310_/LO VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput556 _253_/LO VGND VGND VPWR VPWR la_data_out[86] sky130_fd_sc_hd__clkbuf_2
Xoutput567 _263_/LO VGND VGND VPWR VPWR la_data_out[96] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput589 _320_/LO VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__067__B1 _066_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__076__A _348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input245_A la_oenb[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__058__B1 _345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_287_ VGND VGND VPWR VPWR _287_/HI _287_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output464_A _285_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 io_in[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_1
XFILLER_64_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput375 _118_/LO VGND VGND VPWR VPWR io_oeb[16] sky130_fd_sc_hd__clkbuf_2
Xoutput386 _128_/LO VGND VGND VPWR VPWR io_oeb[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput397 _137_/LO VGND VGND VPWR VPWR io_oeb[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ VGND VGND VPWR VPWR _210_/HI _210_/LO sky130_fd_sc_hd__conb_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ VGND VGND VPWR VPWR _141_/HI _141_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input195_A la_oenb[125] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_072_ _072_/A VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__buf_8
XANTENNA_input362_A wbs_sel_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input56_A la_data_in[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output581_A _313_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_339_ _349_/CLK _339_/D VGND VGND VPWR VPWR _339_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__333__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input208_A la_oenb[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_in[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_124_ VGND VGND VPWR VPWR _124_/HI _124_/LO sky130_fd_sc_hd__conb_1
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_055_ _349_/Q _052_/X _348_/Q _053_/X VGND VGND VPWR VPWR _348_/D sky130_fd_sc_hd__a22o_2
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output427_A _332_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput30 io_in[36] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__buf_1
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput41 la_data_in[101] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__buf_1
Xinput52 la_data_in[111] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__buf_1
Xinput63 la_data_in[121] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__buf_1
Xinput85 la_data_in[26] VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_1
Xinput74 la_data_in[16] VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__buf_1
Xinput96 la_data_in[36] VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_1
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input158_A la_data_in[92] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input325_A wbs_adr_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input19_A io_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output377_A _120_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ VGND VGND VPWR VPWR _107_/HI _107_/LO sky130_fd_sc_hd__conb_1
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output544_A _242_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__100__A2 _052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__079__A _347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input275_A la_oenb[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput220 la_oenb[32] VGND VGND VPWR VPWR input220/X sky130_fd_sc_hd__buf_1
Xinput242 la_oenb[52] VGND VGND VPWR VPWR input242/X sky130_fd_sc_hd__buf_1
Xinput253 la_oenb[62] VGND VGND VPWR VPWR input253/X sky130_fd_sc_hd__buf_1
Xinput231 la_oenb[42] VGND VGND VPWR VPWR input231/X sky130_fd_sc_hd__buf_1
XFILLER_48_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput297 wbs_adr_i[0] VGND VGND VPWR VPWR input297/X sky130_fd_sc_hd__buf_1
Xinput264 la_oenb[72] VGND VGND VPWR VPWR input264/X sky130_fd_sc_hd__buf_1
Xinput275 la_oenb[82] VGND VGND VPWR VPWR input275/X sky130_fd_sc_hd__buf_1
Xinput286 la_oenb[92] VGND VGND VPWR VPWR input286/X sky130_fd_sc_hd__buf_1
XFILLER_90_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output494_A _169_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input86_A la_data_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output507_A _208_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput502 _204_/LO VGND VGND VPWR VPWR la_data_out[37] sky130_fd_sc_hd__clkbuf_2
Xoutput535 _234_/LO VGND VGND VPWR VPWR la_data_out[67] sky130_fd_sc_hd__clkbuf_2
Xoutput513 _214_/LO VGND VGND VPWR VPWR la_data_out[47] sky130_fd_sc_hd__clkbuf_2
Xoutput524 _224_/LO VGND VGND VPWR VPWR la_data_out[57] sky130_fd_sc_hd__clkbuf_2
Xoutput546 _244_/LO VGND VGND VPWR VPWR la_data_out[77] sky130_fd_sc_hd__clkbuf_2
Xoutput557 _254_/LO VGND VGND VPWR VPWR la_data_out[87] sky130_fd_sc_hd__clkbuf_2
Xoutput568 _264_/LO VGND VGND VPWR VPWR la_data_out[97] sky130_fd_sc_hd__clkbuf_2
Xoutput579 _311_/LO VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__067__A1 _342_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__058__A1 _346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input238_A la_oenb[49] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input140_A la_data_in[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__058__B2 _053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_286_ VGND VGND VPWR VPWR _286_/HI _286_/LO sky130_fd_sc_hd__conb_1
XFILLER_115_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output457_A _278_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput6 io_in[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__buf_1
XFILLER_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput376 _119_/LO VGND VGND VPWR VPWR io_oeb[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput387 _129_/LO VGND VGND VPWR VPWR io_oeb[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput398 _138_/LO VGND VGND VPWR VPWR io_oeb[37] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ VGND VGND VPWR VPWR _140_/HI _140_/LO sky130_fd_sc_hd__conb_1
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__buf_4
XANTENNA_input188_A la_oenb[119] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input355_A wbs_dat_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input49_A la_data_in[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ _350_/CLK _338_/D VGND VGND VPWR VPWR _338_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output574_A _297_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_269_ VGND VGND VPWR VPWR _269_/HI _269_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input103_A la_data_in[42] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_123_ VGND VGND VPWR VPWR _123_/HI _123_/LO sky130_fd_sc_hd__conb_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_054_ _350_/Q _052_/X _349_/Q _053_/X VGND VGND VPWR VPWR _349_/D sky130_fd_sc_hd__a22o_4
XFILLER_109_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput20 io_in[27] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_1
Xinput31 io_in[37] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__buf_1
Xinput42 la_data_in[102] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__buf_1
Xinput53 la_data_in[112] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_1
Xinput64 la_data_in[122] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_1
XFILLER_116_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput75 la_data_in[17] VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_1
Xinput86 la_data_in[27] VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_1
Xinput97 la_data_in[37] VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_1
XANTENNA__340__D _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input318_A wbs_adr_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input220_A la_oenb[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ VGND VGND VPWR VPWR _106_/HI _106_/LO sky130_fd_sc_hd__conb_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output537_A _236_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__335__D _335_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__095__A _344_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__346__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input170_A la_oenb[102] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input268_A la_oenb[76] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput210 la_oenb[23] VGND VGND VPWR VPWR input210/X sky130_fd_sc_hd__buf_1
XFILLER_68_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input31_A io_in[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput254 la_oenb[63] VGND VGND VPWR VPWR input254/X sky130_fd_sc_hd__buf_1
Xinput243 la_oenb[53] VGND VGND VPWR VPWR input243/X sky130_fd_sc_hd__buf_1
Xinput221 la_oenb[33] VGND VGND VPWR VPWR input221/X sky130_fd_sc_hd__buf_1
Xinput232 la_oenb[43] VGND VGND VPWR VPWR input232/X sky130_fd_sc_hd__buf_1
Xinput265 la_oenb[73] VGND VGND VPWR VPWR input265/X sky130_fd_sc_hd__buf_1
Xinput276 la_oenb[83] VGND VGND VPWR VPWR input276/X sky130_fd_sc_hd__buf_1
Xinput287 la_oenb[93] VGND VGND VPWR VPWR input287/X sky130_fd_sc_hd__buf_1
XFILLER_75_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput298 wbs_adr_i[10] VGND VGND VPWR VPWR input298/X sky130_fd_sc_hd__buf_1
XFILLER_29_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output487_A _190_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input79_A la_data_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output402_A _110_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput503 _205_/LO VGND VGND VPWR VPWR la_data_out[38] sky130_fd_sc_hd__clkbuf_2
Xoutput536 _235_/LO VGND VGND VPWR VPWR la_data_out[68] sky130_fd_sc_hd__clkbuf_2
Xoutput525 _225_/LO VGND VGND VPWR VPWR la_data_out[58] sky130_fd_sc_hd__clkbuf_2
Xoutput514 _215_/LO VGND VGND VPWR VPWR la_data_out[48] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput547 _245_/LO VGND VGND VPWR VPWR la_data_out[78] sky130_fd_sc_hd__clkbuf_2
Xoutput558 _255_/LO VGND VGND VPWR VPWR la_data_out[88] sky130_fd_sc_hd__clkbuf_2
Xoutput569 _265_/LO VGND VGND VPWR VPWR la_data_out[98] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__067__A2 _063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__058__A2 _052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input133_A la_data_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input300_A wbs_adr_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_285_ VGND VGND VPWR VPWR _285_/HI _285_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 io_in[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_1
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__343__D _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput377 _120_/LO VGND VGND VPWR VPWR io_oeb[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput399 _107_/LO VGND VGND VPWR VPWR io_oeb[3] sky130_fd_sc_hd__clkbuf_2
Xoutput388 _103_/HI VGND VGND VPWR VPWR io_oeb[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_070_ _331_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__buf_4
XFILLER_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input348_A wbs_dat_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input250_A la_oenb[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ _349_/CLK _337_/D VGND VGND VPWR VPWR _337_/Q sky130_fd_sc_hd__dfxtp_4
X_268_ VGND VGND VPWR VPWR _268_/HI _268_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_199_ VGND VGND VPWR VPWR _199_/HI _199_/LO sky130_fd_sc_hd__conb_1
XFILLER_115_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__338__D _338_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input298_A wbs_adr_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_122_ VGND VGND VPWR VPWR _122_/HI _122_/LO sky130_fd_sc_hd__conb_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_053_ _334_/Q VGND VGND VPWR VPWR _053_/X sky130_fd_sc_hd__buf_6
XFILLER_109_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input61_A la_data_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput10 io_in[18] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__buf_1
Xinput21 io_in[28] VGND VGND VPWR VPWR _098_/B1 sky130_fd_sc_hd__clkbuf_2
Xinput43 la_data_in[103] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__buf_1
Xinput54 la_data_in[113] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_1
Xinput32 io_in[3] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__buf_1
Xinput76 la_data_in[18] VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__buf_1
Xinput98 la_data_in[38] VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__buf_1
Xinput87 la_data_in[28] VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__buf_1
Xinput65 la_data_in[123] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__buf_1
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input213_A la_oenb[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_105_ VGND VGND VPWR VPWR _105_/HI _105_/LO sky130_fd_sc_hd__conb_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output432_A _338_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__095__B _095_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input163_A la_data_in[97] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput211 la_oenb[24] VGND VGND VPWR VPWR input211/X sky130_fd_sc_hd__buf_1
Xinput200 la_oenb[14] VGND VGND VPWR VPWR input200/X sky130_fd_sc_hd__buf_1
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input330_A wbs_dat_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput222 la_oenb[34] VGND VGND VPWR VPWR input222/X sky130_fd_sc_hd__buf_1
Xinput244 la_oenb[54] VGND VGND VPWR VPWR input244/X sky130_fd_sc_hd__buf_1
Xinput233 la_oenb[44] VGND VGND VPWR VPWR input233/X sky130_fd_sc_hd__buf_1
XFILLER_68_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput266 la_oenb[74] VGND VGND VPWR VPWR input266/X sky130_fd_sc_hd__buf_1
Xinput255 la_oenb[64] VGND VGND VPWR VPWR input255/X sky130_fd_sc_hd__buf_1
Xinput277 la_oenb[84] VGND VGND VPWR VPWR input277/X sky130_fd_sc_hd__buf_1
Xinput288 la_oenb[94] VGND VGND VPWR VPWR input288/X sky130_fd_sc_hd__buf_1
XANTENNA_input24_A io_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput299 wbs_adr_i[11] VGND VGND VPWR VPWR input299/X sky130_fd_sc_hd__buf_1
XFILLER_84_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output382_A _124_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__346__D _346_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input280_A la_oenb[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output597_A _328_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput504 _206_/LO VGND VGND VPWR VPWR la_data_out[39] sky130_fd_sc_hd__clkbuf_2
Xoutput526 _226_/LO VGND VGND VPWR VPWR la_data_out[59] sky130_fd_sc_hd__clkbuf_2
Xoutput515 _216_/LO VGND VGND VPWR VPWR la_data_out[49] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput548 _246_/LO VGND VGND VPWR VPWR la_data_out[79] sky130_fd_sc_hd__clkbuf_2
Xoutput537 _236_/LO VGND VGND VPWR VPWR la_data_out[69] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput559 _256_/LO VGND VGND VPWR VPWR la_data_out[89] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__336__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input126_A la_data_in[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_284_ VGND VGND VPWR VPWR _284_/HI _284_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input91_A la_data_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 io_in[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__buf_1
XANTENNA_output512_A _213_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput378 _121_/LO VGND VGND VPWR VPWR io_oeb[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput389 _130_/LO VGND VGND VPWR VPWR io_oeb[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input243_A la_oenb[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_336_ _349_/CLK _336_/D VGND VGND VPWR VPWR _336_/Q sky130_fd_sc_hd__dfxtp_2
X_267_ VGND VGND VPWR VPWR _267_/HI _267_/LO sky130_fd_sc_hd__conb_1
X_198_ VGND VGND VPWR VPWR _198_/HI _198_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output462_A _283_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ VGND VGND VPWR VPWR _121_/HI _121_/LO sky130_fd_sc_hd__conb_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input193_A la_oenb[123] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_052_ _052_/A VGND VGND VPWR VPWR _052_/X sky130_fd_sc_hd__buf_6
XFILLER_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input360_A wbs_dat_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input54_A la_data_in[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput11 io_in[19] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_1
X_319_ VGND VGND VPWR VPWR _319_/HI _319_/LO sky130_fd_sc_hd__conb_1
Xinput22 io_in[29] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_1
Xinput44 la_data_in[104] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_1
Xinput55 la_data_in[114] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_1
Xinput33 io_in[4] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__buf_1
XFILLER_115_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput88 la_data_in[29] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__buf_1
Xinput77 la_data_in[19] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__buf_1
Xinput66 la_data_in[124] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__buf_1
Xinput99 la_data_in[39] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__buf_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__349__D _349_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input206_A la_oenb[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_104_ VGND VGND VPWR VPWR _104_/HI _104_/LO sky130_fd_sc_hd__conb_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output425_A _331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput201 la_oenb[15] VGND VGND VPWR VPWR input201/X sky130_fd_sc_hd__buf_1
XANTENNA_input156_A la_data_in[90] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput212 la_oenb[25] VGND VGND VPWR VPWR input212/X sky130_fd_sc_hd__buf_1
Xinput245 la_oenb[55] VGND VGND VPWR VPWR input245/X sky130_fd_sc_hd__buf_1
Xinput223 la_oenb[35] VGND VGND VPWR VPWR input223/X sky130_fd_sc_hd__buf_1
Xinput234 la_oenb[45] VGND VGND VPWR VPWR input234/X sky130_fd_sc_hd__buf_1
XFILLER_48_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input323_A wbs_adr_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput267 la_oenb[75] VGND VGND VPWR VPWR input267/X sky130_fd_sc_hd__buf_1
Xinput256 la_oenb[65] VGND VGND VPWR VPWR input256/X sky130_fd_sc_hd__buf_1
Xinput278 la_oenb[85] VGND VGND VPWR VPWR input278/X sky130_fd_sc_hd__buf_1
XANTENNA_input17_A io_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput289 la_oenb[95] VGND VGND VPWR VPWR input289/X sky130_fd_sc_hd__buf_1
XFILLER_17_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output375_A _118_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output542_A _240_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input9_A io_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input273_A la_oenb[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output492_A _195_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput516 _171_/LO VGND VGND VPWR VPWR la_data_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput505 _170_/LO VGND VGND VPWR VPWR la_data_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput527 _172_/LO VGND VGND VPWR VPWR la_data_out[5] sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_1_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput538 _173_/LO VGND VGND VPWR VPWR la_data_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput549 _174_/LO VGND VGND VPWR VPWR la_data_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input119_A la_data_in[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_283_ VGND VGND VPWR VPWR _283_/HI _283_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input84_A la_data_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 io_in[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_1
XANTENNA_output505_A _170_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput368 _104_/LO VGND VGND VPWR VPWR io_oeb[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput379 _105_/LO VGND VGND VPWR VPWR io_oeb[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input236_A la_oenb[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_335_ _349_/CLK _335_/D VGND VGND VPWR VPWR _335_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_266_ VGND VGND VPWR VPWR _266_/HI _266_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_197_ VGND VGND VPWR VPWR _197_/HI _197_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output455_A _177_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__349__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_120_ VGND VGND VPWR VPWR _120_/HI _120_/LO sky130_fd_sc_hd__conb_1
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_051_ _062_/A VGND VGND VPWR VPWR _052_/A sky130_fd_sc_hd__clkinv_8
XFILLER_3_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input186_A la_oenb[117] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input353_A wbs_dat_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input47_A la_data_in[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput12 io_in[1] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_1
X_318_ VGND VGND VPWR VPWR _318_/HI _318_/LO sky130_fd_sc_hd__conb_1
X_249_ VGND VGND VPWR VPWR _249_/HI _249_/LO sky130_fd_sc_hd__conb_1
Xinput45 la_data_in[105] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_1
Xinput23 io_in[2] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__buf_1
Xinput34 io_in[5] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__buf_1
XFILLER_116_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput89 la_data_in[2] VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__buf_1
Xinput78 la_data_in[1] VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_1
Xinput56 la_data_in[115] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_1
Xinput67 la_data_in[125] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__buf_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input101_A la_data_in[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_103_ VGND VGND VPWR VPWR _103_/HI _103_/LO sky130_fd_sc_hd__conb_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output418_A _159_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput202 la_oenb[16] VGND VGND VPWR VPWR input202/X sky130_fd_sc_hd__buf_1
Xinput213 la_oenb[26] VGND VGND VPWR VPWR input213/X sky130_fd_sc_hd__buf_1
Xinput224 la_oenb[36] VGND VGND VPWR VPWR input224/X sky130_fd_sc_hd__buf_1
Xinput235 la_oenb[46] VGND VGND VPWR VPWR input235/X sky130_fd_sc_hd__buf_1
XANTENNA_input149_A la_data_in[84] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput268 la_oenb[76] VGND VGND VPWR VPWR input268/X sky130_fd_sc_hd__buf_1
Xinput257 la_oenb[66] VGND VGND VPWR VPWR input257/X sky130_fd_sc_hd__buf_1
Xinput246 la_oenb[56] VGND VGND VPWR VPWR input246/X sky130_fd_sc_hd__buf_1
Xinput279 la_oenb[86] VGND VGND VPWR VPWR input279/X sky130_fd_sc_hd__buf_1
XFILLER_48_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input316_A wbs_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output368_A _104_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output535_A _234_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input266_A la_oenb[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output485_A _188_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput506 _207_/LO VGND VGND VPWR VPWR la_data_out[40] sky130_fd_sc_hd__clkbuf_2
Xoutput517 _217_/LO VGND VGND VPWR VPWR la_data_out[50] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput539 _237_/LO VGND VGND VPWR VPWR la_data_out[70] sky130_fd_sc_hd__clkbuf_2
Xoutput528 _227_/LO VGND VGND VPWR VPWR la_data_out[60] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_282_ VGND VGND VPWR VPWR _282_/HI _282_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input77_A la_data_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output400_A _108_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput369 _112_/LO VGND VGND VPWR VPWR io_oeb[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input131_A la_data_in[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input229_A la_oenb[40] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _350_/CLK _334_/D hold1/X VGND VGND VPWR VPWR _334_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_265_ VGND VGND VPWR VPWR _265_/HI _265_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_196_ VGND VGND VPWR VPWR _196_/HI _196_/LO sky130_fd_sc_hd__conb_1
XFILLER_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output448_A _270_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__060__B1 _343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_050_ _072_/A _333_/Q VGND VGND VPWR VPWR _062_/A sky130_fd_sc_hd__nand2_8
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input179_A la_oenb[110] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input346_A wbs_dat_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output398_A _138_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_317_ VGND VGND VPWR VPWR _317_/HI _317_/LO sky130_fd_sc_hd__conb_1
Xinput13 io_in[20] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_1
XFILLER_30_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_248_ VGND VGND VPWR VPWR _248_/HI _248_/LO sky130_fd_sc_hd__conb_1
Xinput46 la_data_in[106] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_1
Xinput35 io_in[6] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__buf_1
Xinput24 io_in[30] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_1
X_179_ VGND VGND VPWR VPWR _179_/HI _179_/LO sky130_fd_sc_hd__conb_1
Xinput79 la_data_in[20] VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__buf_1
XANTENNA_output565_A _261_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput57 la_data_in[116] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_1
Xinput68 la_data_in[126] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__buf_1
XFILLER_115_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input296_A wb_rst_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_102_ VGND VGND VPWR VPWR _102_/HI _102_/LO sky130_fd_sc_hd__conb_1
XFILLER_113_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__339__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput203 la_oenb[17] VGND VGND VPWR VPWR input203/X sky130_fd_sc_hd__buf_1
Xinput214 la_oenb[27] VGND VGND VPWR VPWR input214/X sky130_fd_sc_hd__buf_1
Xinput236 la_oenb[47] VGND VGND VPWR VPWR input236/X sky130_fd_sc_hd__buf_1
Xinput225 la_oenb[37] VGND VGND VPWR VPWR input225/X sky130_fd_sc_hd__buf_1
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput269 la_oenb[77] VGND VGND VPWR VPWR input269/X sky130_fd_sc_hd__buf_1
Xinput258 la_oenb[67] VGND VGND VPWR VPWR input258/X sky130_fd_sc_hd__buf_1
Xinput247 la_oenb[57] VGND VGND VPWR VPWR input247/X sky130_fd_sc_hd__buf_1
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input211_A la_oenb[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input309_A wbs_adr_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output528_A _227_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output430_A _336_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input259_A la_oenb[68] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input161_A la_data_in[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input22_A io_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output478_A _182_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput507 _208_/LO VGND VGND VPWR VPWR la_data_out[41] sky130_fd_sc_hd__clkbuf_2
Xoutput518 _218_/LO VGND VGND VPWR VPWR la_data_out[51] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput529 _228_/LO VGND VGND VPWR VPWR la_data_out[61] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ _350_/CLK _350_/D VGND VGND VPWR VPWR _350_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_281_ VGND VGND VPWR VPWR _281_/HI _281_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output595_A _326_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input124_A la_data_in[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ _349_/CLK _333_/D hold1/X VGND VGND VPWR VPWR _333_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ VGND VGND VPWR VPWR _264_/HI _264_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_195_ VGND VGND VPWR VPWR _195_/HI _195_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output510_A _211_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__060__B2 _334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__060__A1 _344_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input339_A wbs_dat_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input241_A la_oenb[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_316_ VGND VGND VPWR VPWR _316_/HI _316_/LO sky130_fd_sc_hd__conb_1
XFILLER_30_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput14 io_in[21] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__buf_1
X_247_ VGND VGND VPWR VPWR _247_/HI _247_/LO sky130_fd_sc_hd__conb_1
Xinput36 io_in[7] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__buf_1
Xinput25 io_in[31] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__buf_1
XFILLER_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_178_ VGND VGND VPWR VPWR _178_/HI _178_/LO sky130_fd_sc_hd__conb_1
Xinput47 la_data_in[107] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_1
Xinput58 la_data_in[117] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_1
Xinput69 la_data_in[127] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_1
XANTENNA_output460_A _281_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output558_A _255_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_101_ VGND VGND VPWR VPWR _101_/HI _101_/LO sky130_fd_sc_hd__conb_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input191_A la_oenb[121] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input289_A la_oenb[95] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input52_A la_data_in[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput226 la_oenb[38] VGND VGND VPWR VPWR input226/X sky130_fd_sc_hd__buf_1
Xinput204 la_oenb[18] VGND VGND VPWR VPWR input204/X sky130_fd_sc_hd__buf_1
Xinput215 la_oenb[28] VGND VGND VPWR VPWR input215/X sky130_fd_sc_hd__buf_1
XFILLER_88_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput248 la_oenb[58] VGND VGND VPWR VPWR input248/X sky130_fd_sc_hd__buf_1
Xinput259 la_oenb[68] VGND VGND VPWR VPWR input259/X sky130_fd_sc_hd__buf_1
Xinput237 la_oenb[48] VGND VGND VPWR VPWR input237/X sky130_fd_sc_hd__buf_1
XFILLER_75_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input204_A la_oenb[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output423_A _164_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input154_A la_data_in[89] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input321_A wbs_adr_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input15_A io_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output373_A _116_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput508 _209_/LO VGND VGND VPWR VPWR la_data_out[42] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput519 _219_/LO VGND VGND VPWR VPWR la_data_out[52] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output540_A _238_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input7_A io_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__081__C1 _080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_280_ VGND VGND VPWR VPWR _280_/HI _280_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input271_A la_oenb[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output490_A _193_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output588_A _319_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input117_A la_data_in[55] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _332_/A VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__clkbuf_4
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ VGND VGND VPWR VPWR _263_/HI _263_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input82_A la_data_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_194_ VGND VGND VPWR VPWR _194_/HI _194_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output503_A _205_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__060__A2 _052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input234_A la_oenb[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_315_ VGND VGND VPWR VPWR _315_/HI _315_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput15 io_in[22] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_1
Xinput37 io_in[8] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_1
Xinput26 io_in[32] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__buf_1
X_246_ VGND VGND VPWR VPWR _246_/HI _246_/LO sky130_fd_sc_hd__conb_1
X_177_ VGND VGND VPWR VPWR _177_/HI _177_/LO sky130_fd_sc_hd__conb_1
Xinput48 la_data_in[108] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__buf_1
Xinput59 la_data_in[118] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_1
XFILLER_115_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output453_A _275_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_100_ _063_/A _052_/X _071_/X VGND VGND VPWR VPWR _350_/D sky130_fd_sc_hd__o21ai_4
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input184_A la_oenb[115] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input351_A wbs_dat_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input45_A la_data_in[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output570_A _266_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_229_ VGND VGND VPWR VPWR _229_/HI _229_/LO sky130_fd_sc_hd__conb_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput216 la_oenb[29] VGND VGND VPWR VPWR input216/X sky130_fd_sc_hd__buf_1
Xinput205 la_oenb[19] VGND VGND VPWR VPWR input205/X sky130_fd_sc_hd__buf_1
Xinput227 la_oenb[39] VGND VGND VPWR VPWR input227/X sky130_fd_sc_hd__buf_1
Xinput238 la_oenb[49] VGND VGND VPWR VPWR input238/X sky130_fd_sc_hd__buf_1
Xinput249 la_oenb[59] VGND VGND VPWR VPWR input249/X sky130_fd_sc_hd__buf_1
XFILLER_75_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output416_A _158_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input147_A la_data_in[82] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input314_A wbs_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput509 _210_/LO VGND VGND VPWR VPWR la_data_out[43] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output533_A _232_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__090__B1 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__081__B1 _071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input264_A la_oenb[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output483_A _168_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__054__B1 _349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_331_ _331_/A VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__buf_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ VGND VGND VPWR VPWR _262_/HI _262_/LO sky130_fd_sc_hd__conb_1
X_193_ VGND VGND VPWR VPWR _193_/HI _193_/LO sky130_fd_sc_hd__conb_1
XFILLER_108_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input75_A la_data_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input227_A la_oenb[39] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_314_ VGND VGND VPWR VPWR _314_/HI _314_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_245_ VGND VGND VPWR VPWR _245_/HI _245_/LO sky130_fd_sc_hd__conb_1
XFILLER_52_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput16 io_in[23] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_1
Xinput27 io_in[33] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__buf_1
Xinput38 io_in[9] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_1
X_176_ VGND VGND VPWR VPWR _176_/HI _176_/LO sky130_fd_sc_hd__conb_1
Xinput49 la_data_in[109] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_1
XFILLER_108_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output446_A _268_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input177_A la_oenb[109] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input344_A wbs_dat_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input38_A io_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_228_ VGND VGND VPWR VPWR _228_/HI _228_/LO sky130_fd_sc_hd__conb_1
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output563_A _259_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_159_ VGND VGND VPWR VPWR _159_/HI _159_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_26_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput217 la_oenb[2] VGND VGND VPWR VPWR input217/X sky130_fd_sc_hd__buf_1
Xinput206 la_oenb[1] VGND VGND VPWR VPWR input206/X sky130_fd_sc_hd__buf_1
Xinput239 la_oenb[4] VGND VGND VPWR VPWR input239/X sky130_fd_sc_hd__buf_1
Xinput228 la_oenb[3] VGND VGND VPWR VPWR input228/X sky130_fd_sc_hd__buf_1
XFILLER_29_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input294_A la_oenb[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output409_A _151_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input307_A wbs_adr_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output526_A _226_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__090__A1 _088_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__081__A1 _079_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input257_A la_oenb[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input20_A io_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output476_A _180_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__052__A _052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__054__B2 _053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__054__A1 _350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ VGND VGND VPWR VPWR _330_/HI _330_/LO sky130_fd_sc_hd__conb_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ VGND VGND VPWR VPWR _261_/HI _261_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_192_ VGND VGND VPWR VPWR _192_/HI _192_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input68_A la_data_in[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output593_A _324_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input122_A la_data_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_313_ VGND VGND VPWR VPWR _313_/HI _313_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_244_ VGND VGND VPWR VPWR _244_/HI _244_/LO sky130_fd_sc_hd__conb_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 io_in[24] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_1
Xinput28 io_in[34] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__buf_1
Xinput39 la_data_in[0] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__buf_1
X_175_ VGND VGND VPWR VPWR _175_/HI _175_/LO sky130_fd_sc_hd__conb_1
XFILLER_108_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output439_A _144_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output606_A _307_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput490 _193_/LO VGND VGND VPWR VPWR la_data_out[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input337_A wbs_dat_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_227_ VGND VGND VPWR VPWR _227_/HI _227_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output389_A _130_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_158_ VGND VGND VPWR VPWR _158_/HI _158_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output556_A _253_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_089_ _072_/A _073_/A _345_/Q _336_/Q VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__a31o_1
XFILLER_97_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput218 la_oenb[30] VGND VGND VPWR VPWR input218/X sky130_fd_sc_hd__buf_1
Xinput207 la_oenb[20] VGND VGND VPWR VPWR input207/X sky130_fd_sc_hd__buf_1
Xinput229 la_oenb[40] VGND VGND VPWR VPWR input229/X sky130_fd_sc_hd__buf_1
XFILLER_29_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input287_A la_oenb[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input50_A la_data_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__093__C1 _092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__084__C1 _083_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input202_A la_oenb[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input98_A la_data_in[38] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output421_A _162_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__075__C1 _074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output519_A _219_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__090__A2 _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__081__A2 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input152_A la_data_in[87] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input13_A io_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__342__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output371_A _114_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output469_A _289_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input5_A io_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__054__A2 _052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ VGND VGND VPWR VPWR _260_/HI _260_/LO sky130_fd_sc_hd__conb_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_191_ VGND VGND VPWR VPWR _191_/HI _191_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input367_A wbs_we_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output586_A _318_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__063__A _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input115_A la_data_in[53] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_312_ VGND VGND VPWR VPWR _312_/HI _312_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_243_ VGND VGND VPWR VPWR _243_/HI _243_/LO sky130_fd_sc_hd__conb_1
Xinput18 io_in[25] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__buf_1
XANTENNA_input80_A la_data_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput29 io_in[35] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_1
X_174_ VGND VGND VPWR VPWR _174_/HI _174_/LO sky130_fd_sc_hd__conb_1
XFILLER_97_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output501_A _203_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput480 _184_/LO VGND VGND VPWR VPWR la_data_out[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput491 _194_/LO VGND VGND VPWR VPWR la_data_out[27] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input232_A la_oenb[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_226_ VGND VGND VPWR VPWR _226_/HI _226_/LO sky130_fd_sc_hd__conb_1
X_157_ VGND VGND VPWR VPWR _157_/HI _157_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_088_ _344_/Q VGND VGND VPWR VPWR _088_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output549_A _174_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output451_A _273_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput208 la_oenb[21] VGND VGND VPWR VPWR input208/X sky130_fd_sc_hd__buf_1
Xinput219 la_oenb[31] VGND VGND VPWR VPWR input219/X sky130_fd_sc_hd__buf_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input182_A la_oenb[113] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input43_A la_data_in[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output499_A _201_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ VGND VGND VPWR VPWR _209_/HI _209_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__093__B1 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_adc.COMP_clk _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__071__A _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__084__B1 _071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__075__B1 _071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output414_A _156_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__090__A3 _331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__081__A3 _070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__066__A _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input145_A la_data_in[80] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__057__B1 _346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input312_A wbs_adr_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output531_A _230_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_190_ VGND VGND VPWR VPWR _190_/HI _190_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input262_A la_oenb[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output481_A _185_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output579_A _311_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__063__B _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input108_A la_data_in[47] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_311_ VGND VGND VPWR VPWR _311_/HI _311_/LO sky130_fd_sc_hd__conb_1
X_242_ VGND VGND VPWR VPWR _242_/HI _242_/LO sky130_fd_sc_hd__conb_1
Xinput19 io_in[26] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__buf_1
X_173_ VGND VGND VPWR VPWR _173_/HI _173_/LO sky130_fd_sc_hd__conb_1
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input73_A la_data_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput470 _290_/LO VGND VGND VPWR VPWR la_data_out[123] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput492 _195_/LO VGND VGND VPWR VPWR la_data_out[28] sky130_fd_sc_hd__clkbuf_2
Xoutput481 _185_/LO VGND VGND VPWR VPWR la_data_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input225_A la_oenb[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_225_ VGND VGND VPWR VPWR _225_/HI _225_/LO sky130_fd_sc_hd__conb_1
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_156_ VGND VGND VPWR VPWR _156_/HI _156_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ _085_/Y _069_/A _070_/X _071_/A _086_/X VGND VGND VPWR VPWR _337_/D sky130_fd_sc_hd__o311a_2
XFILLER_6_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output444_A _167_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput209 la_oenb[22] VGND VGND VPWR VPWR input209/X sky130_fd_sc_hd__buf_1
XFILLER_102_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__069__A _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input175_A la_oenb[107] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input342_A wbs_dat_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input36_A io_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output394_A _134_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ VGND VGND VPWR VPWR _208_/HI _208_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output561_A _257_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_139_ VGND VGND VPWR VPWR _139_/HI _139_/LO sky130_fd_sc_hd__conb_1
XFILLER_99_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__093__A1 _095_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__084__A1 _082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input292_A la_oenb[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__075__A1 _068_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output407_A _149_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__082__A _346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__057__A1 _347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__057__B2 _053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input138_A la_data_in[74] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input305_A wbs_adr_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output524_A _224_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input255_A la_oenb[64] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output474_A _294_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__063__C _331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_310_ VGND VGND VPWR VPWR _310_/HI _310_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_241_ VGND VGND VPWR VPWR _241_/HI _241_/LO sky130_fd_sc_hd__conb_1
X_172_ VGND VGND VPWR VPWR _172_/HI _172_/LO sky130_fd_sc_hd__conb_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input66_A la_data_in[124] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output591_A _322_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput460 _281_/LO VGND VGND VPWR VPWR la_data_out[114] sky130_fd_sc_hd__clkbuf_2
Xoutput471 _291_/LO VGND VGND VPWR VPWR la_data_out[124] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput493 _196_/LO VGND VGND VPWR VPWR la_data_out[29] sky130_fd_sc_hd__clkbuf_2
Xoutput482 _186_/LO VGND VGND VPWR VPWR la_data_out[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input218_A la_oenb[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input120_A la_data_in[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_224_ VGND VGND VPWR VPWR _224_/HI _224_/LO sky130_fd_sc_hd__conb_1
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_155_ VGND VGND VPWR VPWR _155_/HI _155_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_086_ _072_/A _073_/A _346_/Q _337_/Q VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__a31o_1
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output437_A _142_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output604_A _305_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__085__A _345_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input168_A la_oenb[100] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__087__C1 _086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input335_A wbs_dat_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input29_A io_in[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__345__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output387_A _129_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_207_ VGND VGND VPWR VPWR _207_/HI _207_/LO sky130_fd_sc_hd__conb_1
X_138_ VGND VGND VPWR VPWR _138_/HI _138_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output554_A _251_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_069_ _069_/A VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_99_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__078__C1 _077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__093__A2 _331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__084__A2 _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input285_A la_oenb[91] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__075__A2 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__057__A2 _052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input200_A la_oenb[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input96_A la_data_in[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput360 wbs_dat_i[8] VGND VGND VPWR VPWR input360/X sky130_fd_sc_hd__buf_1
XFILLER_48_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__333__D _333_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input150_A la_data_in[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input248_A la_oenb[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input11_A io_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output467_A _287_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput190 la_oenb[120] VGND VGND VPWR VPWR input190/X sky130_fd_sc_hd__buf_1
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input3_A io_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__088__A _344_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_240_ VGND VGND VPWR VPWR _240_/HI _240_/LO sky130_fd_sc_hd__conb_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_171_ VGND VGND VPWR VPWR _171_/HI _171_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input198_A la_oenb[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input365_A wbs_sel_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input59_A la_data_in[118] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output584_A _316_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput450 _272_/LO VGND VGND VPWR VPWR la_data_out[105] sky130_fd_sc_hd__clkbuf_2
Xoutput461 _282_/LO VGND VGND VPWR VPWR la_data_out[115] sky130_fd_sc_hd__clkbuf_2
Xoutput494 _169_/LO VGND VGND VPWR VPWR la_data_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput483 _168_/LO VGND VGND VPWR VPWR la_data_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput472 _292_/LO VGND VGND VPWR VPWR la_data_out[125] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input113_A la_data_in[51] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ VGND VGND VPWR VPWR _223_/HI _223_/LO sky130_fd_sc_hd__conb_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_154_ VGND VGND VPWR VPWR _154_/HI _154_/LO sky130_fd_sc_hd__conb_1
X_085_ _345_/Q VGND VGND VPWR VPWR _085_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__341__D _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__087__B1 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input230_A la_oenb[41] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input328_A wbs_adr_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_206_ VGND VGND VPWR VPWR _206_/HI _206_/LO sky130_fd_sc_hd__conb_1
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_137_ VGND VGND VPWR VPWR _137_/HI _137_/LO sky130_fd_sc_hd__conb_1
X_068_ _349_/Q VGND VGND VPWR VPWR _068_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_98_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__078__B1 _071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__093__A3 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__336__D _336_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__084__A3 _070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__096__A _350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input180_A la_oenb[111] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_oenb[85] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input41_A la_data_in[101] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__075__A3 _070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output497_A _199_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__335__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input89_A la_data_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput350 wbs_dat_i[28] VGND VGND VPWR VPWR input350/X sky130_fd_sc_hd__buf_1
Xinput361 wbs_dat_i[9] VGND VGND VPWR VPWR input361/X sky130_fd_sc_hd__buf_1
XFILLER_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output412_A _154_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input143_A la_data_in[79] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input310_A wbs_adr_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput180 la_oenb[111] VGND VGND VPWR VPWR input180/X sky130_fd_sc_hd__buf_1
XFILLER_64_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput191 la_oenb[121] VGND VGND VPWR VPWR input191/X sky130_fd_sc_hd__buf_1
XFILLER_48_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ VGND VGND VPWR VPWR _170_/HI _170_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input260_A la_oenb[69] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input358_A wbs_dat_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output577_A _309_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_299_ VGND VGND VPWR VPWR _299_/HI _299_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__339__D _339_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput451 _273_/LO VGND VGND VPWR VPWR la_data_out[106] sky130_fd_sc_hd__clkbuf_2
Xoutput462 _283_/LO VGND VGND VPWR VPWR la_data_out[116] sky130_fd_sc_hd__clkbuf_2
Xoutput440 _145_/LO VGND VGND VPWR VPWR io_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput495 _197_/LO VGND VGND VPWR VPWR la_data_out[30] sky130_fd_sc_hd__clkbuf_2
Xoutput484 _187_/LO VGND VGND VPWR VPWR la_data_out[20] sky130_fd_sc_hd__clkbuf_2
Xoutput473 _293_/LO VGND VGND VPWR VPWR la_data_out[126] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A la_data_in[45] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_222_ VGND VGND VPWR VPWR _222_/HI _222_/LO sky130_fd_sc_hd__conb_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_153_ VGND VGND VPWR VPWR _153_/HI _153_/LO sky130_fd_sc_hd__conb_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_084_ _082_/Y _069_/A _070_/X _071_/X _083_/X VGND VGND VPWR VPWR _338_/D sky130_fd_sc_hd__o311a_2
XANTENNA_input71_A la_data_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input223_A la_oenb[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_205_ VGND VGND VPWR VPWR _205_/HI _205_/LO sky130_fd_sc_hd__conb_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_136_ VGND VGND VPWR VPWR _136_/HI _136_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_067_ _342_/Q _063_/X _066_/Y VGND VGND VPWR VPWR _342_/D sky130_fd_sc_hd__a21o_2
XANTENNA_output442_A _147_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__078__A1 _076_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__096__B _349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input173_A la_oenb[105] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input340_A wbs_dat_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input34_A io_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output392_A _132_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_119_ VGND VGND VPWR VPWR _119_/HI _119_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__347__D _347_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input290_A la_oenb[96] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput351 wbs_dat_i[29] VGND VGND VPWR VPWR input351/X sky130_fd_sc_hd__buf_1
Xinput362 wbs_sel_i[0] VGND VGND VPWR VPWR input362/X sky130_fd_sc_hd__buf_1
Xinput340 wbs_dat_i[19] VGND VGND VPWR VPWR input340/X sky130_fd_sc_hd__buf_1
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input136_A la_data_in[72] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input303_A wbs_adr_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output522_A _222_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput170 la_oenb[102] VGND VGND VPWR VPWR input170/X sky130_fd_sc_hd__buf_1
Xinput181 la_oenb[112] VGND VGND VPWR VPWR input181/X sky130_fd_sc_hd__buf_1
Xinput192 la_oenb[122] VGND VGND VPWR VPWR input192/X sky130_fd_sc_hd__buf_1
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput600 _330_/LO VGND VGND VPWR VPWR wbs_dat_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input253_A la_oenb[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__348__CLK _349_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_298_ VGND VGND VPWR VPWR _298_/HI _298_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output472_A _292_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput452 _274_/LO VGND VGND VPWR VPWR la_data_out[107] sky130_fd_sc_hd__clkbuf_2
Xoutput430 _336_/Q VGND VGND VPWR VPWR io_out[31] sky130_fd_sc_hd__clkbuf_2
Xoutput441 _146_/LO VGND VGND VPWR VPWR io_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput496 _198_/LO VGND VGND VPWR VPWR la_data_out[31] sky130_fd_sc_hd__clkbuf_2
Xoutput485 _188_/LO VGND VGND VPWR VPWR la_data_out[21] sky130_fd_sc_hd__clkbuf_2
Xoutput463 _284_/LO VGND VGND VPWR VPWR la_data_out[117] sky130_fd_sc_hd__clkbuf_2
Xoutput474 _294_/LO VGND VGND VPWR VPWR la_data_out[127] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__099__B _099_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_221_ VGND VGND VPWR VPWR _221_/HI _221_/LO sky130_fd_sc_hd__conb_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_152_ VGND VGND VPWR VPWR _152_/HI _152_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_083_ _094_/A _094_/B _347_/Q _338_/Q VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__a31o_2
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input64_A la_data_in[122] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__087__A2 _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input216_A la_oenb[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_204_ VGND VGND VPWR VPWR _204_/HI _204_/LO sky130_fd_sc_hd__conb_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_135_ VGND VGND VPWR VPWR _135_/HI _135_/LO sky130_fd_sc_hd__conb_1
X_066_ _071_/A VGND VGND VPWR VPWR _066_/Y sky130_fd_sc_hd__inv_4
XFILLER_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__078__A2 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output435_A _341_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__096__C _348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input166_A la_data_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input333_A wbs_dat_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input27_A io_in[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output385_A _127_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_118_ VGND VGND VPWR VPWR _118_/HI _118_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output552_A _249_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_049_ _334_/Q VGND VGND VPWR VPWR _072_/A sky130_fd_sc_hd__clkinv_8
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input283_A la_oenb[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput330 wbs_dat_i[0] VGND VGND VPWR VPWR input330/X sky130_fd_sc_hd__buf_1
XFILLER_88_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput352 wbs_dat_i[2] VGND VGND VPWR VPWR input352/X sky130_fd_sc_hd__buf_1
Xinput341 wbs_dat_i[1] VGND VGND VPWR VPWR input341/X sky130_fd_sc_hd__buf_1
Xinput363 wbs_sel_i[1] VGND VGND VPWR VPWR input363/X sky130_fd_sc_hd__buf_1
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input129_A la_data_in[66] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input94_A la_data_in[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output515_A _216_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput160 la_data_in[94] VGND VGND VPWR VPWR input160/X sky130_fd_sc_hd__buf_1
Xinput171 la_oenb[103] VGND VGND VPWR VPWR input171/X sky130_fd_sc_hd__buf_1
Xinput182 la_oenb[113] VGND VGND VPWR VPWR input182/X sky130_fd_sc_hd__buf_1
Xinput193 la_oenb[123] VGND VGND VPWR VPWR input193/X sky130_fd_sc_hd__buf_1
XFILLER_17_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput601 _302_/LO VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input246_A la_oenb[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_297_ VGND VGND VPWR VPWR _297_/HI _297_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput420 _161_/LO VGND VGND VPWR VPWR io_out[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput442 _147_/LO VGND VGND VPWR VPWR io_out[8] sky130_fd_sc_hd__clkbuf_2
Xoutput453 _275_/LO VGND VGND VPWR VPWR la_data_out[108] sky130_fd_sc_hd__clkbuf_2
Xoutput431 _337_/Q VGND VGND VPWR VPWR io_out[32] sky130_fd_sc_hd__clkbuf_2
Xoutput486 _189_/LO VGND VGND VPWR VPWR la_data_out[22] sky130_fd_sc_hd__clkbuf_2
Xoutput475 _179_/LO VGND VGND VPWR VPWR la_data_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput464 _285_/LO VGND VGND VPWR VPWR la_data_out[118] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput497 _199_/LO VGND VGND VPWR VPWR la_data_out[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input1_A io_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_220_ VGND VGND VPWR VPWR _220_/HI _220_/LO sky130_fd_sc_hd__conb_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_151_ VGND VGND VPWR VPWR _151_/HI _151_/LO sky130_fd_sc_hd__conb_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input196_A la_oenb[126] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ _346_/Q VGND VGND VPWR VPWR _082_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input363_A wbs_sel_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input57_A la_data_in[116] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output582_A _314_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_349_ _349_/CLK _349_/D VGND VGND VPWR VPWR _349_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_115_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__338__CLK _350_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__087__A3 _070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xadc.COMP analog_io[1] analog_io[0] _331_/A adc.COMP/VDD adc.COMP/VSS _349_/CLK VPWR
+ VGND ACMP
XANTENNA_input111_A la_data_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input209_A la_oenb[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_203_ VGND VGND VPWR VPWR _203_/HI _203_/LO sky130_fd_sc_hd__conb_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_134_ VGND VGND VPWR VPWR _134_/HI _134_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_065_ _334_/Q _073_/A VGND VGND VPWR VPWR _071_/A sky130_fd_sc_hd__or2_4
XFILLER_3_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__078__A3 _070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output428_A _141_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__096__D _347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input159_A la_data_in[93] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input326_A wbs_adr_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output378_A _121_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_117_ VGND VGND VPWR VPWR _117_/HI _117_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input276_A la_oenb[83] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput320 wbs_adr_i[30] VGND VGND VPWR VPWR input320/X sky130_fd_sc_hd__buf_1
XFILLER_96_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput353 wbs_dat_i[30] VGND VGND VPWR VPWR input353/X sky130_fd_sc_hd__buf_1
Xinput331 wbs_dat_i[10] VGND VGND VPWR VPWR input331/X sky130_fd_sc_hd__buf_1
Xinput342 wbs_dat_i[20] VGND VGND VPWR VPWR input342/X sky130_fd_sc_hd__buf_1
XFILLER_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput364 wbs_sel_i[2] VGND VGND VPWR VPWR input364/X sky130_fd_sc_hd__buf_1
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output495_A _197_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_adc.COMP_INN analog_io[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input87_A la_data_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput150 la_data_in[85] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__buf_1
Xinput161 la_data_in[95] VGND VGND VPWR VPWR input161/X sky130_fd_sc_hd__buf_1
Xinput172 la_oenb[104] VGND VGND VPWR VPWR input172/X sky130_fd_sc_hd__buf_1
XANTENNA_output410_A _152_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output508_A _209_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput183 la_oenb[114] VGND VGND VPWR VPWR input183/X sky130_fd_sc_hd__buf_1
Xinput194 la_oenb[124] VGND VGND VPWR VPWR input194/X sky130_fd_sc_hd__buf_1
XFILLER_36_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput602 _303_/LO VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_98_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input239_A la_oenb[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input141_A la_data_in[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_296_ VGND VGND VPWR VPWR _296_/HI _296_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output458_A _279_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput410 _152_/LO VGND VGND VPWR VPWR io_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput421 _162_/LO VGND VGND VPWR VPWR io_out[23] sky130_fd_sc_hd__clkbuf_2
Xoutput443 _148_/LO VGND VGND VPWR VPWR io_out[9] sky130_fd_sc_hd__clkbuf_2
Xoutput432 _338_/Q VGND VGND VPWR VPWR io_out[33] sky130_fd_sc_hd__clkbuf_2
Xoutput487 _190_/LO VGND VGND VPWR VPWR la_data_out[23] sky130_fd_sc_hd__clkbuf_2
Xoutput476 _180_/LO VGND VGND VPWR VPWR la_data_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput454 _276_/LO VGND VGND VPWR VPWR la_data_out[109] sky130_fd_sc_hd__clkbuf_2
Xoutput465 _286_/LO VGND VGND VPWR VPWR la_data_out[119] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput498 _200_/LO VGND VGND VPWR VPWR la_data_out[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_150_ VGND VGND VPWR VPWR _150_/HI _150_/LO sky130_fd_sc_hd__conb_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input189_A la_oenb[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_081_ _079_/Y _099_/A _070_/X _071_/X _080_/X VGND VGND VPWR VPWR _339_/D sky130_fd_sc_hd__o311a_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input356_A wbs_dat_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_348_ _349_/CLK _348_/D VGND VGND VPWR VPWR _348_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_output575_A _298_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_279_ VGND VGND VPWR VPWR _279_/HI _279_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input104_A la_data_in[43] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_202_ VGND VGND VPWR VPWR _202_/HI _202_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_133_ VGND VGND VPWR VPWR _133_/HI _133_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_064_ _333_/Q VGND VGND VPWR VPWR _073_/A sky130_fd_sc_hd__buf_6
XFILLER_3_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input319_A wbs_adr_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input221_A la_oenb[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_116_ VGND VGND VPWR VPWR _116_/HI _116_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output440_A _145_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output538_A _173_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input171_A la_oenb[103] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input269_A la_oenb[77] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput321 wbs_adr_i[31] VGND VGND VPWR VPWR input321/X sky130_fd_sc_hd__buf_1
Xinput310 wbs_adr_i[21] VGND VGND VPWR VPWR input310/X sky130_fd_sc_hd__buf_1
Xinput354 wbs_dat_i[31] VGND VGND VPWR VPWR input354/X sky130_fd_sc_hd__buf_1
Xinput343 wbs_dat_i[21] VGND VGND VPWR VPWR input343/X sky130_fd_sc_hd__buf_1
Xinput332 wbs_dat_i[11] VGND VGND VPWR VPWR input332/X sky130_fd_sc_hd__buf_1
XANTENNA_input32_A io_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput365 wbs_sel_i[3] VGND VGND VPWR VPWR input365/X sky130_fd_sc_hd__buf_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output488_A _191_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output390_A _106_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput140 la_data_in[76] VGND VGND VPWR VPWR input140/X sky130_fd_sc_hd__buf_1
Xinput151 la_data_in[86] VGND VGND VPWR VPWR input151/X sky130_fd_sc_hd__buf_1
Xinput162 la_data_in[96] VGND VGND VPWR VPWR input162/X sky130_fd_sc_hd__buf_1
XFILLER_64_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput173 la_oenb[105] VGND VGND VPWR VPWR input173/X sky130_fd_sc_hd__buf_1
Xinput184 la_oenb[115] VGND VGND VPWR VPWR input184/X sky130_fd_sc_hd__buf_1
Xinput195 la_oenb[125] VGND VGND VPWR VPWR input195/X sky130_fd_sc_hd__buf_1
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput603 _304_/LO VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input134_A la_data_in[70] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input301_A wbs_adr_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_295_ VGND VGND VPWR VPWR _295_/HI _295_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output520_A _220_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput411 _153_/LO VGND VGND VPWR VPWR io_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput400 _108_/LO VGND VGND VPWR VPWR io_oeb[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput422 _163_/LO VGND VGND VPWR VPWR io_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput444 _167_/LO VGND VGND VPWR VPWR la_data_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput433 _339_/Q VGND VGND VPWR VPWR io_out[34] sky130_fd_sc_hd__clkbuf_2
Xoutput455 _177_/LO VGND VGND VPWR VPWR la_data_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput466 _178_/LO VGND VGND VPWR VPWR la_data_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput477 _181_/LO VGND VGND VPWR VPWR la_data_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput499 _201_/LO VGND VGND VPWR VPWR la_data_out[34] sky130_fd_sc_hd__clkbuf_2
Xoutput488 _191_/LO VGND VGND VPWR VPWR la_data_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_080_ _094_/A _094_/B _348_/Q _339_/Q VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__a31o_4
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input349_A wbs_dat_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input251_A la_oenb[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_347_ _349_/CLK _347_/D VGND VGND VPWR VPWR _347_/Q sky130_fd_sc_hd__dfxtp_4
X_278_ VGND VGND VPWR VPWR _278_/HI _278_/LO sky130_fd_sc_hd__conb_1
XANTENNA_output568_A _264_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output470_A _290_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_201_ VGND VGND VPWR VPWR _201_/HI _201_/LO sky130_fd_sc_hd__conb_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_132_ VGND VGND VPWR VPWR _132_/HI _132_/LO sky130_fd_sc_hd__conb_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input299_A wbs_adr_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_063_ _063_/A _069_/A _331_/A VGND VGND VPWR VPWR _063_/X sky130_fd_sc_hd__or3_4
XFILLER_109_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input62_A la_data_in[120] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input214_A la_oenb[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_115_ VGND VGND VPWR VPWR _115_/HI _115_/LO sky130_fd_sc_hd__conb_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output433_A _339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__080__B1 _339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input164_A la_data_in[98] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput300 wbs_adr_i[12] VGND VGND VPWR VPWR input300/X sky130_fd_sc_hd__buf_1
Xinput311 wbs_adr_i[22] VGND VGND VPWR VPWR input311/X sky130_fd_sc_hd__buf_1
XFILLER_102_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput344 wbs_dat_i[22] VGND VGND VPWR VPWR input344/X sky130_fd_sc_hd__buf_1
XANTENNA_input331_A wbs_dat_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput322 wbs_adr_i[3] VGND VGND VPWR VPWR input322/X sky130_fd_sc_hd__buf_1
Xinput333 wbs_dat_i[12] VGND VGND VPWR VPWR input333/X sky130_fd_sc_hd__buf_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput355 wbs_dat_i[3] VGND VGND VPWR VPWR input355/X sky130_fd_sc_hd__buf_1
Xinput366 wbs_stb_i VGND VGND VPWR VPWR input366/X sky130_fd_sc_hd__buf_1
XANTENNA_input25_A io_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output383_A _125_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_adc.COMP_INP analog_io[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output550_A _247_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input281_A la_oenb[88] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput141 la_data_in[77] VGND VGND VPWR VPWR input141/X sky130_fd_sc_hd__buf_1
Xinput130 la_data_in[67] VGND VGND VPWR VPWR input130/X sky130_fd_sc_hd__buf_1
Xinput152 la_data_in[87] VGND VGND VPWR VPWR input152/X sky130_fd_sc_hd__buf_1
Xinput163 la_data_in[97] VGND VGND VPWR VPWR input163/X sky130_fd_sc_hd__buf_1
XFILLER_64_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput174 la_oenb[106] VGND VGND VPWR VPWR input174/X sky130_fd_sc_hd__buf_1
Xinput185 la_oenb[116] VGND VGND VPWR VPWR input185/X sky130_fd_sc_hd__buf_1
Xinput196 la_oenb[126] VGND VGND VPWR VPWR input196/X sky130_fd_sc_hd__buf_1
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output598_A _301_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput604 _305_/LO VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

