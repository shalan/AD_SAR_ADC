magic
tech sky130A
magscale 1 2
timestamp 1626122236
<< locali >>
rect 58081 44183 58115 44489
rect 68937 34935 68971 35581
rect 27629 15895 27663 16541
rect 21373 13379 21407 13481
rect 37381 12903 37415 13277
rect 24501 4879 24535 5525
rect 2513 2907 2547 3145
rect 19073 3111 19107 4097
rect 19165 3179 19199 4029
rect 19165 1819 19199 2601
rect 19257 2567 19291 4437
rect 20729 3179 20763 3485
rect 21741 2907 21775 3213
rect 22109 1955 22143 3213
rect 22477 1479 22511 3077
rect 22569 2703 22603 3553
rect 22937 2159 22971 3689
rect 23397 2703 23431 2805
rect 25237 1819 25271 5525
rect 25329 1887 25363 2941
rect 25605 1887 25639 2805
rect 25789 1887 25823 3281
rect 25881 1887 25915 3417
rect 26065 1887 26099 3077
rect 26341 1955 26375 3145
rect 26525 1955 26559 3757
rect 26617 1955 26651 3009
rect 26801 1887 26835 2873
rect 26893 1955 26927 4029
rect 27169 1955 27203 3621
rect 27353 1887 27387 3621
rect 27445 1955 27479 3281
rect 27629 1955 27663 2805
rect 27905 1955 27939 3893
rect 28641 1751 28675 4505
rect 28733 1955 28767 3689
rect 29009 1955 29043 3961
rect 29193 1955 29227 3349
rect 29469 1547 29503 3145
rect 29561 1751 29595 3077
rect 30297 1547 30331 3825
rect 30481 1343 30515 3417
rect 30573 1547 30607 4097
rect 30757 1343 30791 3485
rect 30849 1547 30883 3553
rect 30941 1683 30975 1989
rect 31125 1683 31159 3757
rect 31309 1683 31343 2873
rect 31493 1547 31527 9401
rect 31585 3655 31619 6205
rect 31769 4879 31803 5525
rect 31953 4675 31987 5593
rect 32045 4879 32079 5525
rect 32321 4879 32355 5525
rect 32505 4879 32539 5525
rect 32689 3519 32723 4165
rect 31585 1683 31619 3213
rect 32965 2839 32999 5185
rect 32171 2805 32321 2839
rect 33333 2703 33367 3757
rect 33425 2567 33459 5049
rect 33609 2363 33643 8517
rect 33885 3111 33919 3689
rect 33977 2567 34011 3213
rect 34069 1003 34103 9537
rect 34161 1955 34195 3689
rect 34345 1275 34379 4437
rect 34437 1955 34471 8585
rect 37381 6239 37415 6817
rect 34989 4539 35023 5185
rect 34897 3179 34931 3485
rect 34989 3383 35023 3485
rect 35725 3179 35759 3893
rect 35817 3655 35851 4029
rect 37289 3519 37323 3961
rect 37473 3655 37507 7837
rect 37381 3315 37415 3485
rect 35633 3111 35667 3145
rect 35633 3077 35759 3111
rect 35725 2907 35759 3077
rect 35449 1819 35483 2397
rect 36001 1343 36035 2805
rect 37289 2023 37323 2329
rect 36461 1479 36495 1921
rect 36553 1615 36587 1853
rect 39773 1071 39807 2057
<< viali >>
rect 16497 67337 16531 67371
rect 1777 67269 1811 67303
rect 2881 67269 2915 67303
rect 8677 67269 8711 67303
rect 10609 67269 10643 67303
rect 18429 67269 18463 67303
rect 24225 67269 24259 67303
rect 26157 67269 26191 67303
rect 32045 67269 32079 67303
rect 33977 67269 34011 67303
rect 39773 67269 39807 67303
rect 41705 67269 41739 67303
rect 47593 67269 47627 67303
rect 49617 67269 49651 67303
rect 55321 67269 55355 67303
rect 57621 67269 57655 67303
rect 63141 67269 63175 67303
rect 65625 67269 65659 67303
rect 67373 67269 67407 67303
rect 4997 67133 5031 67167
rect 5457 67133 5491 67167
rect 12725 67133 12759 67167
rect 13185 67133 13219 67167
rect 20545 67133 20579 67167
rect 21005 67133 21039 67167
rect 24409 67133 24443 67167
rect 28457 67133 28491 67167
rect 28917 67133 28951 67167
rect 36461 67133 36495 67167
rect 36921 67133 36955 67167
rect 44465 67133 44499 67167
rect 44925 67133 44959 67167
rect 52469 67133 52503 67167
rect 52929 67133 52963 67167
rect 59369 67133 59403 67167
rect 59921 67133 59955 67167
rect 66637 67133 66671 67167
rect 1961 67065 1995 67099
rect 3065 67065 3099 67099
rect 8493 67065 8527 67099
rect 10793 67065 10827 67099
rect 16589 67065 16623 67099
rect 17233 67065 17267 67099
rect 18613 67065 18647 67099
rect 26341 67065 26375 67099
rect 32229 67065 32263 67099
rect 34161 67065 34195 67099
rect 39957 67065 39991 67099
rect 41889 67065 41923 67099
rect 47777 67065 47811 67099
rect 49801 67065 49835 67099
rect 55505 67065 55539 67099
rect 57805 67065 57839 67099
rect 63325 67065 63359 67099
rect 65809 67065 65843 67099
rect 67189 67065 67223 67099
rect 67925 67065 67959 67099
rect 3893 66997 3927 67031
rect 9321 66997 9355 67031
rect 19165 66997 19199 67031
rect 25605 66997 25639 67031
rect 33241 66997 33275 67031
rect 39221 66997 39255 67031
rect 50445 66997 50479 67031
rect 54769 66997 54803 67031
rect 62589 66997 62623 67031
rect 64705 66997 64739 67031
rect 33793 66793 33827 66827
rect 66913 66793 66947 66827
rect 68017 66793 68051 66827
rect 1777 66725 1811 66759
rect 1961 66657 1995 66691
rect 2697 66657 2731 66691
rect 3157 66657 3191 66691
rect 57437 66657 57471 66691
rect 66269 66657 66303 66691
rect 67925 66657 67959 66691
rect 3985 66453 4019 66487
rect 11069 66453 11103 66487
rect 30481 66453 30515 66487
rect 41521 66453 41555 66487
rect 65349 66453 65383 66487
rect 2237 66113 2271 66147
rect 66269 66113 66303 66147
rect 1593 66045 1627 66079
rect 14841 66045 14875 66079
rect 36185 66045 36219 66079
rect 36461 66045 36495 66079
rect 65349 66045 65383 66079
rect 65809 66045 65843 66079
rect 65993 66045 66027 66079
rect 66361 66045 66395 66079
rect 68109 66045 68143 66079
rect 64705 65977 64739 66011
rect 34253 65909 34287 65943
rect 34897 65909 34931 65943
rect 36921 65909 36955 65943
rect 66729 65909 66763 65943
rect 65533 65705 65567 65739
rect 68109 65705 68143 65739
rect 1961 65569 1995 65603
rect 44649 65433 44683 65467
rect 1869 65365 1903 65399
rect 2605 65365 2639 65399
rect 23029 65365 23063 65399
rect 48697 65365 48731 65399
rect 66821 65365 66855 65399
rect 17325 64957 17359 64991
rect 41337 64957 41371 64991
rect 66913 64957 66947 64991
rect 67517 64957 67551 64991
rect 67741 64957 67775 64991
rect 66361 64889 66395 64923
rect 67373 64889 67407 64923
rect 67925 64889 67959 64923
rect 67649 64821 67683 64855
rect 2237 64277 2271 64311
rect 52469 64277 52503 64311
rect 67005 64277 67039 64311
rect 15393 64005 15427 64039
rect 14289 63937 14323 63971
rect 68109 63937 68143 63971
rect 14013 63869 14047 63903
rect 14749 63869 14783 63903
rect 67925 63801 67959 63835
rect 12909 63733 12943 63767
rect 67281 63733 67315 63767
rect 11345 63393 11379 63427
rect 11989 63393 12023 63427
rect 67925 63393 67959 63427
rect 11897 63257 11931 63291
rect 68109 63257 68143 63291
rect 12725 63189 12759 63223
rect 13185 63189 13219 63223
rect 48881 63189 48915 63223
rect 67281 63189 67315 63223
rect 67373 62985 67407 63019
rect 7021 62917 7055 62951
rect 36829 62849 36863 62883
rect 49341 62849 49375 62883
rect 1593 62781 1627 62815
rect 2053 62781 2087 62815
rect 9781 62781 9815 62815
rect 47409 62781 47443 62815
rect 67281 62781 67315 62815
rect 49617 62713 49651 62747
rect 67097 62713 67131 62747
rect 48789 62645 48823 62679
rect 51089 62645 51123 62679
rect 66545 62645 66579 62679
rect 66913 62441 66947 62475
rect 48973 62373 49007 62407
rect 20269 62305 20303 62339
rect 20361 62305 20395 62339
rect 21005 62237 21039 62271
rect 13553 62169 13587 62203
rect 36921 61829 36955 61863
rect 17509 61693 17543 61727
rect 1961 61625 1995 61659
rect 1869 61557 1903 61591
rect 2513 61557 2547 61591
rect 67465 61217 67499 61251
rect 68109 61217 68143 61251
rect 51457 60673 51491 60707
rect 1777 60129 1811 60163
rect 1961 60129 1995 60163
rect 2513 60129 2547 60163
rect 52233 60129 52267 60163
rect 52377 60129 52411 60163
rect 52469 60129 52503 60163
rect 52653 60129 52687 60163
rect 57161 60129 57195 60163
rect 15669 60061 15703 60095
rect 44373 59925 44407 59959
rect 47409 59925 47443 59959
rect 51457 59925 51491 59959
rect 52101 59925 52135 59959
rect 53205 59925 53239 59959
rect 16129 59517 16163 59551
rect 16405 59517 16439 59551
rect 67097 59517 67131 59551
rect 17049 59449 17083 59483
rect 14841 59381 14875 59415
rect 17509 59381 17543 59415
rect 51641 59381 51675 59415
rect 52837 59381 52871 59415
rect 10517 58973 10551 59007
rect 43269 58905 43303 58939
rect 13461 58837 13495 58871
rect 64337 58837 64371 58871
rect 48789 58565 48823 58599
rect 68109 58565 68143 58599
rect 23213 58497 23247 58531
rect 44005 58497 44039 58531
rect 44097 58497 44131 58531
rect 44281 58497 44315 58531
rect 22753 58429 22787 58463
rect 27997 58429 28031 58463
rect 34529 58429 34563 58463
rect 44189 58429 44223 58463
rect 67925 58361 67959 58395
rect 42533 58293 42567 58327
rect 43269 58293 43303 58327
rect 43821 58293 43855 58327
rect 67281 58293 67315 58327
rect 6837 58089 6871 58123
rect 6009 58021 6043 58055
rect 65533 58021 65567 58055
rect 5641 57953 5675 57987
rect 6101 57953 6135 57987
rect 65073 57953 65107 57987
rect 6377 57885 6411 57919
rect 7481 57885 7515 57919
rect 5457 57817 5491 57851
rect 28089 57817 28123 57851
rect 4721 57749 4755 57783
rect 8217 57749 8251 57783
rect 36185 57749 36219 57783
rect 43453 57749 43487 57783
rect 45293 57749 45327 57783
rect 55137 57749 55171 57783
rect 64429 57749 64463 57783
rect 67281 57545 67315 57579
rect 17325 57477 17359 57511
rect 35633 57409 35667 57443
rect 1593 57341 1627 57375
rect 2053 57341 2087 57375
rect 25513 57341 25547 57375
rect 67925 57341 67959 57375
rect 68109 57273 68143 57307
rect 6929 57205 6963 57239
rect 10793 56661 10827 56695
rect 1777 56321 1811 56355
rect 18245 56253 18279 56287
rect 30297 56253 30331 56287
rect 67465 56253 67499 56287
rect 68109 56253 68143 56287
rect 1961 56185 1995 56219
rect 2513 56117 2547 56151
rect 9965 55777 9999 55811
rect 10057 55709 10091 55743
rect 11069 55573 11103 55607
rect 13093 55573 13127 55607
rect 38025 55573 38059 55607
rect 10241 55301 10275 55335
rect 37381 55301 37415 55335
rect 38761 55301 38795 55335
rect 61117 55301 61151 55335
rect 2605 55233 2639 55267
rect 41981 55233 42015 55267
rect 67189 55233 67223 55267
rect 1961 55165 1995 55199
rect 38577 55165 38611 55199
rect 38669 55165 38703 55199
rect 38853 55165 38887 55199
rect 39037 55165 39071 55199
rect 39589 55097 39623 55131
rect 1869 55029 1903 55063
rect 38393 55029 38427 55063
rect 38117 54485 38151 54519
rect 44833 54485 44867 54519
rect 62129 54485 62163 54519
rect 5641 54077 5675 54111
rect 48789 54077 48823 54111
rect 33333 53737 33367 53771
rect 32321 53669 32355 53703
rect 28089 53601 28123 53635
rect 28733 53601 28767 53635
rect 33057 53601 33091 53635
rect 67925 53601 67959 53635
rect 29377 53533 29411 53567
rect 32873 53533 32907 53567
rect 32965 53533 32999 53567
rect 33149 53533 33183 53567
rect 31769 53465 31803 53499
rect 68109 53465 68143 53499
rect 7757 53397 7791 53431
rect 53941 53397 53975 53431
rect 55505 53397 55539 53431
rect 67281 53397 67315 53431
rect 55781 53193 55815 53227
rect 54677 53125 54711 53159
rect 40693 53057 40727 53091
rect 41337 52989 41371 53023
rect 51089 52989 51123 53023
rect 54401 52989 54435 53023
rect 54585 52989 54619 53023
rect 54769 52989 54803 53023
rect 54861 52989 54895 53023
rect 55597 52989 55631 53023
rect 62865 52989 62899 53023
rect 65257 52989 65291 53023
rect 32137 52921 32171 52955
rect 55045 52921 55079 52955
rect 62773 52921 62807 52955
rect 32781 52853 32815 52887
rect 53021 52853 53055 52887
rect 53849 52853 53883 52887
rect 63233 52649 63267 52683
rect 1593 52513 1627 52547
rect 2053 52513 2087 52547
rect 54033 52445 54067 52479
rect 55321 52445 55355 52479
rect 27077 52309 27111 52343
rect 67281 52105 67315 52139
rect 68109 51969 68143 52003
rect 15853 51901 15887 51935
rect 67925 51901 67959 51935
rect 15301 51425 15335 51459
rect 15853 51425 15887 51459
rect 15117 51357 15151 51391
rect 31493 51357 31527 51391
rect 46213 51357 46247 51391
rect 67373 51221 67407 51255
rect 1869 51017 1903 51051
rect 2605 51017 2639 51051
rect 34437 50881 34471 50915
rect 1961 50813 1995 50847
rect 17969 50813 18003 50847
rect 54217 50813 54251 50847
rect 67465 50813 67499 50847
rect 68109 50813 68143 50847
rect 17601 50745 17635 50779
rect 18613 50677 18647 50711
rect 34437 50201 34471 50235
rect 3157 50133 3191 50167
rect 23305 50133 23339 50167
rect 34897 49861 34931 49895
rect 1777 49793 1811 49827
rect 2605 49793 2639 49827
rect 20085 49793 20119 49827
rect 21373 49793 21407 49827
rect 35449 49793 35483 49827
rect 1961 49725 1995 49759
rect 20821 49725 20855 49759
rect 34345 49725 34379 49759
rect 34529 49725 34563 49759
rect 34718 49725 34752 49759
rect 36001 49725 36035 49759
rect 34621 49657 34655 49691
rect 33793 49589 33827 49623
rect 33977 49045 34011 49079
rect 67925 48161 67959 48195
rect 68109 48025 68143 48059
rect 45017 47957 45051 47991
rect 31769 47209 31803 47243
rect 1869 47141 1903 47175
rect 25421 47073 25455 47107
rect 32413 47073 32447 47107
rect 67925 47073 67959 47107
rect 26065 47005 26099 47039
rect 2053 46937 2087 46971
rect 32597 46937 32631 46971
rect 39681 46937 39715 46971
rect 49617 46937 49651 46971
rect 67281 46937 67315 46971
rect 68109 46937 68143 46971
rect 1685 46665 1719 46699
rect 7573 46529 7607 46563
rect 21281 46461 21315 46495
rect 2513 46121 2547 46155
rect 1961 46053 1995 46087
rect 1777 45917 1811 45951
rect 39313 45781 39347 45815
rect 39957 45509 39991 45543
rect 58081 45509 58115 45543
rect 13001 45373 13035 45407
rect 39405 45373 39439 45407
rect 40089 45373 40123 45407
rect 40325 45373 40359 45407
rect 40509 45373 40543 45407
rect 67465 45373 67499 45407
rect 68109 45373 68143 45407
rect 40233 45305 40267 45339
rect 40969 45237 41003 45271
rect 1961 44965 1995 44999
rect 2513 44965 2547 44999
rect 58725 44965 58759 44999
rect 59553 44965 59587 44999
rect 17058 44897 17092 44931
rect 58541 44897 58575 44931
rect 58817 44897 58851 44931
rect 58909 44897 58943 44931
rect 17325 44829 17359 44863
rect 15945 44761 15979 44795
rect 59093 44761 59127 44795
rect 1869 44693 1903 44727
rect 15301 44693 15335 44727
rect 17877 44693 17911 44727
rect 39589 44693 39623 44727
rect 58081 44693 58115 44727
rect 58081 44489 58115 44523
rect 58265 44489 58299 44523
rect 10701 44285 10735 44319
rect 58081 44149 58115 44183
rect 30481 43809 30515 43843
rect 31125 43809 31159 43843
rect 62405 43809 62439 43843
rect 62865 43809 62899 43843
rect 62129 43741 62163 43775
rect 30665 43605 30699 43639
rect 35725 43605 35759 43639
rect 65441 43605 65475 43639
rect 2973 43265 3007 43299
rect 3249 43197 3283 43231
rect 4353 43197 4387 43231
rect 13001 43197 13035 43231
rect 13645 43197 13679 43231
rect 50077 43197 50111 43231
rect 1869 43061 1903 43095
rect 3709 43061 3743 43095
rect 13093 43061 13127 43095
rect 49433 42721 49467 42755
rect 67925 42721 67959 42755
rect 68109 42721 68143 42755
rect 48881 42653 48915 42687
rect 50261 42653 50295 42687
rect 11713 42517 11747 42551
rect 12817 42517 12851 42551
rect 20177 42517 20211 42551
rect 18705 42245 18739 42279
rect 1593 42109 1627 42143
rect 2053 42109 2087 42143
rect 26617 42109 26651 42143
rect 51365 42109 51399 42143
rect 17685 41769 17719 41803
rect 67281 41769 67315 41803
rect 30757 41701 30791 41735
rect 31309 41701 31343 41735
rect 67925 41701 67959 41735
rect 16037 41633 16071 41667
rect 17872 41633 17906 41667
rect 17969 41633 18003 41667
rect 18107 41633 18141 41667
rect 18245 41633 18279 41667
rect 32689 41633 32723 41667
rect 33517 41633 33551 41667
rect 32965 41565 32999 41599
rect 18797 41497 18831 41531
rect 35909 41497 35943 41531
rect 68109 41497 68143 41531
rect 16681 41429 16715 41463
rect 57713 41429 57747 41463
rect 43545 41021 43579 41055
rect 47041 41021 47075 41055
rect 66177 41021 66211 41055
rect 17509 40885 17543 40919
rect 18613 40885 18647 40919
rect 1869 40681 1903 40715
rect 1961 40545 1995 40579
rect 22937 40545 22971 40579
rect 23581 40545 23615 40579
rect 2513 40341 2547 40375
rect 23029 40341 23063 40375
rect 67465 39933 67499 39967
rect 68109 39933 68143 39967
rect 2605 39593 2639 39627
rect 1961 39525 1995 39559
rect 1777 39457 1811 39491
rect 29377 39253 29411 39287
rect 33517 39253 33551 39287
rect 34253 38981 34287 39015
rect 34345 38913 34379 38947
rect 34124 38845 34158 38879
rect 48973 38845 49007 38879
rect 33977 38777 34011 38811
rect 34713 38777 34747 38811
rect 33425 38709 33459 38743
rect 35265 38709 35299 38743
rect 33609 38165 33643 38199
rect 40969 38165 41003 38199
rect 46121 37893 46155 37927
rect 35725 37757 35759 37791
rect 40693 37757 40727 37791
rect 67925 37689 67959 37723
rect 68109 37689 68143 37723
rect 1593 36669 1627 36703
rect 2053 36669 2087 36703
rect 5549 36193 5583 36227
rect 67373 36193 67407 36227
rect 67925 36193 67959 36227
rect 68109 36193 68143 36227
rect 41797 36125 41831 36159
rect 42073 36125 42107 36159
rect 2881 35989 2915 36023
rect 41245 35989 41279 36023
rect 43177 35989 43211 36023
rect 51457 35989 51491 36023
rect 1777 35581 1811 35615
rect 7205 35581 7239 35615
rect 44465 35581 44499 35615
rect 55873 35581 55907 35615
rect 61301 35581 61335 35615
rect 61577 35581 61611 35615
rect 67465 35581 67499 35615
rect 68109 35581 68143 35615
rect 68937 35581 68971 35615
rect 1961 35513 1995 35547
rect 2605 35445 2639 35479
rect 41521 35445 41555 35479
rect 60749 35445 60783 35479
rect 62681 35445 62715 35479
rect 30941 35105 30975 35139
rect 31493 35105 31527 35139
rect 67925 35105 67959 35139
rect 32781 34901 32815 34935
rect 60841 34901 60875 34935
rect 68937 34901 68971 34935
rect 8401 34697 8435 34731
rect 9045 34697 9079 34731
rect 64705 34697 64739 34731
rect 32045 34629 32079 34663
rect 33425 34629 33459 34663
rect 34897 34629 34931 34663
rect 7113 34561 7147 34595
rect 33149 34561 33183 34595
rect 45109 34561 45143 34595
rect 6837 34493 6871 34527
rect 9597 34493 9631 34527
rect 30297 34493 30331 34527
rect 33344 34493 33378 34527
rect 33517 34493 33551 34527
rect 33609 34493 33643 34527
rect 33793 34493 33827 34527
rect 44465 34493 44499 34527
rect 34253 34357 34287 34391
rect 1869 34153 1903 34187
rect 32413 34153 32447 34187
rect 32965 34085 32999 34119
rect 1961 34017 1995 34051
rect 10149 34017 10183 34051
rect 2513 33813 2547 33847
rect 55321 33813 55355 33847
rect 36921 33541 36955 33575
rect 25145 33405 25179 33439
rect 39313 33405 39347 33439
rect 62957 33405 62991 33439
rect 64889 32725 64923 32759
rect 7021 32317 7055 32351
rect 67925 32249 67959 32283
rect 68109 32249 68143 32283
rect 36645 31909 36679 31943
rect 55413 31909 55447 31943
rect 55781 31909 55815 31943
rect 56425 31909 56459 31943
rect 1593 31841 1627 31875
rect 2053 31841 2087 31875
rect 26893 31841 26927 31875
rect 27537 31841 27571 31875
rect 37197 31841 37231 31875
rect 37473 31841 37507 31875
rect 37749 31841 37783 31875
rect 37933 31841 37967 31875
rect 39037 31841 39071 31875
rect 54861 31841 54895 31875
rect 55597 31841 55631 31875
rect 37565 31773 37599 31807
rect 38485 31773 38519 31807
rect 37657 31705 37691 31739
rect 42441 31705 42475 31739
rect 36829 31433 36863 31467
rect 25973 30889 26007 30923
rect 37841 30821 37875 30855
rect 67925 30821 67959 30855
rect 68109 30821 68143 30855
rect 8125 30753 8159 30787
rect 25421 30753 25455 30787
rect 37697 30753 37731 30787
rect 37933 30753 37967 30787
rect 38117 30753 38151 30787
rect 39129 30753 39163 30787
rect 4445 30617 4479 30651
rect 25237 30549 25271 30583
rect 36921 30549 36955 30583
rect 37565 30549 37599 30583
rect 38577 30549 38611 30583
rect 1777 30277 1811 30311
rect 2697 30277 2731 30311
rect 37105 30277 37139 30311
rect 49065 30209 49099 30243
rect 12081 30141 12115 30175
rect 27813 30141 27847 30175
rect 38945 30141 38979 30175
rect 48605 30141 48639 30175
rect 49157 30141 49191 30175
rect 1961 30073 1995 30107
rect 27077 29801 27111 29835
rect 27169 29801 27203 29835
rect 28457 29801 28491 29835
rect 27997 29733 28031 29767
rect 26893 29665 26927 29699
rect 27261 29665 27295 29699
rect 35909 29665 35943 29699
rect 67465 29665 67499 29699
rect 68109 29665 68143 29699
rect 27445 29529 27479 29563
rect 2237 29461 2271 29495
rect 7021 29461 7055 29495
rect 21005 29461 21039 29495
rect 26341 29461 26375 29495
rect 27905 29189 27939 29223
rect 1777 29053 1811 29087
rect 1961 29053 1995 29087
rect 2513 29053 2547 29087
rect 29101 29053 29135 29087
rect 59277 29053 59311 29087
rect 30941 28713 30975 28747
rect 54953 28509 54987 28543
rect 13461 28169 13495 28203
rect 31493 28169 31527 28203
rect 32781 28169 32815 28203
rect 18705 28101 18739 28135
rect 17693 28033 17727 28067
rect 31033 28033 31067 28067
rect 31769 28033 31803 28067
rect 31677 27965 31711 27999
rect 31861 27965 31895 27999
rect 31953 27965 31987 27999
rect 32137 27965 32171 27999
rect 35817 27965 35851 27999
rect 60473 27965 60507 27999
rect 33241 27829 33275 27863
rect 17805 27489 17839 27523
rect 18061 27421 18095 27455
rect 16681 27353 16715 27387
rect 7665 27285 7699 27319
rect 18521 27285 18555 27319
rect 31125 27285 31159 27319
rect 64981 27285 65015 27319
rect 18797 27081 18831 27115
rect 67281 27081 67315 27115
rect 68109 26945 68143 26979
rect 1593 26877 1627 26911
rect 2053 26877 2087 26911
rect 31401 26877 31435 26911
rect 67925 26877 67959 26911
rect 18245 26741 18279 26775
rect 43085 26537 43119 26571
rect 47409 26537 47443 26571
rect 50353 26537 50387 26571
rect 27905 26469 27939 26503
rect 29561 26469 29595 26503
rect 47869 26469 47903 26503
rect 24225 26401 24259 26435
rect 28181 26401 28215 26435
rect 28457 26401 28491 26435
rect 29009 26401 29043 26435
rect 30205 26401 30239 26435
rect 38025 26401 38059 26435
rect 42533 26401 42567 26435
rect 42625 26401 42659 26435
rect 48881 26401 48915 26435
rect 49249 26401 49283 26435
rect 49433 26401 49467 26435
rect 49617 26401 49651 26435
rect 49801 26401 49835 26435
rect 48513 26333 48547 26367
rect 1777 26265 1811 26299
rect 27353 26265 27387 26299
rect 62681 26265 62715 26299
rect 27813 25993 27847 26027
rect 67373 25993 67407 26027
rect 55505 25925 55539 25959
rect 67925 25789 67959 25823
rect 55781 25721 55815 25755
rect 68109 25721 68143 25755
rect 47685 25653 47719 25687
rect 48421 25653 48455 25687
rect 11989 25449 12023 25483
rect 66177 25449 66211 25483
rect 1961 25313 1995 25347
rect 11345 25313 11379 25347
rect 10977 25245 11011 25279
rect 1777 25177 1811 25211
rect 2605 25109 2639 25143
rect 7941 25109 7975 25143
rect 36921 24701 36955 24735
rect 64521 24701 64555 24735
rect 67465 24701 67499 24735
rect 68109 24701 68143 24735
rect 23489 24361 23523 24395
rect 21925 24225 21959 24259
rect 22845 24225 22879 24259
rect 33701 24225 33735 24259
rect 67925 24157 67959 24191
rect 12357 24021 12391 24055
rect 29101 24021 29135 24055
rect 54125 24021 54159 24055
rect 1869 23817 1903 23851
rect 2605 23817 2639 23851
rect 57345 23681 57379 23715
rect 1961 23613 1995 23647
rect 53021 23613 53055 23647
rect 54309 23613 54343 23647
rect 54401 23613 54435 23647
rect 54585 23613 54619 23647
rect 53849 23545 53883 23579
rect 54769 23477 54803 23511
rect 56425 23477 56459 23511
rect 58449 23273 58483 23307
rect 67373 23273 67407 23307
rect 53941 23205 53975 23239
rect 55781 23205 55815 23239
rect 67925 23205 67959 23239
rect 56701 23069 56735 23103
rect 56977 23069 57011 23103
rect 68109 23001 68143 23035
rect 11713 22933 11747 22967
rect 37933 22933 37967 22967
rect 30481 22729 30515 22763
rect 39681 22729 39715 22763
rect 62037 22729 62071 22763
rect 9229 22661 9263 22695
rect 13185 22661 13219 22695
rect 29929 22661 29963 22695
rect 7297 22593 7331 22627
rect 7021 22525 7055 22559
rect 30660 22525 30694 22559
rect 31033 22525 31067 22559
rect 32045 22525 32079 22559
rect 38301 22525 38335 22559
rect 38577 22525 38611 22559
rect 46397 22525 46431 22559
rect 30757 22457 30791 22491
rect 30849 22457 30883 22491
rect 31493 22457 31527 22491
rect 8585 22389 8619 22423
rect 9781 22389 9815 22423
rect 56609 22389 56643 22423
rect 30113 22185 30147 22219
rect 38117 22185 38151 22219
rect 15301 21845 15335 21879
rect 67281 21641 67315 21675
rect 68109 21573 68143 21607
rect 1409 21437 1443 21471
rect 2421 21437 2455 21471
rect 13093 21437 13127 21471
rect 31493 21437 31527 21471
rect 33609 21437 33643 21471
rect 36093 21437 36127 21471
rect 67925 21437 67959 21471
rect 1409 21097 1443 21131
rect 33149 20825 33183 20859
rect 37289 20757 37323 20791
rect 27813 20553 27847 20587
rect 28457 20553 28491 20587
rect 29285 20349 29319 20383
rect 30297 20349 30331 20383
rect 67465 20349 67499 20383
rect 68109 20349 68143 20383
rect 1869 20009 1903 20043
rect 27261 20009 27295 20043
rect 30021 20009 30055 20043
rect 1961 19873 1995 19907
rect 2605 19873 2639 19907
rect 29009 19873 29043 19907
rect 29285 19873 29319 19907
rect 29469 19873 29503 19907
rect 30941 19873 30975 19907
rect 31861 19873 31895 19907
rect 31677 19805 31711 19839
rect 28825 19737 28859 19771
rect 29101 19737 29135 19771
rect 29193 19737 29227 19771
rect 28273 19669 28307 19703
rect 33977 19669 34011 19703
rect 50445 19669 50479 19703
rect 53297 19669 53331 19703
rect 49709 19329 49743 19363
rect 67925 19193 67959 19227
rect 68109 19193 68143 19227
rect 67281 19125 67315 19159
rect 2513 18921 2547 18955
rect 1961 18853 1995 18887
rect 51273 18785 51307 18819
rect 1777 18649 1811 18683
rect 9505 18581 9539 18615
rect 18245 18377 18279 18411
rect 61485 18377 61519 18411
rect 17693 18105 17727 18139
rect 17785 17833 17819 17867
rect 67281 17833 67315 17867
rect 67925 17765 67959 17799
rect 17509 17697 17543 17731
rect 17877 17697 17911 17731
rect 68109 17697 68143 17731
rect 47685 17493 47719 17527
rect 10057 17085 10091 17119
rect 18245 17085 18279 17119
rect 55781 17085 55815 17119
rect 61577 17085 61611 17119
rect 56517 16609 56551 16643
rect 56701 16609 56735 16643
rect 57161 16609 57195 16643
rect 67465 16609 67499 16643
rect 68109 16609 68143 16643
rect 27629 16541 27663 16575
rect 18245 16405 18279 16439
rect 18061 16201 18095 16235
rect 1593 15997 1627 16031
rect 2053 15997 2087 16031
rect 7021 15997 7055 16031
rect 56517 16473 56551 16507
rect 56149 16201 56183 16235
rect 27629 15861 27663 15895
rect 11345 15657 11379 15691
rect 67741 15657 67775 15691
rect 5917 15521 5951 15555
rect 10517 15521 10551 15555
rect 11437 15521 11471 15555
rect 17693 15317 17727 15351
rect 18245 15317 18279 15351
rect 9781 15113 9815 15147
rect 68109 14977 68143 15011
rect 66361 14909 66395 14943
rect 67189 14909 67223 14943
rect 67925 14909 67959 14943
rect 1961 14841 1995 14875
rect 17325 14841 17359 14875
rect 1869 14773 1903 14807
rect 2605 14773 2639 14807
rect 18245 14773 18279 14807
rect 15209 14569 15243 14603
rect 17325 14569 17359 14603
rect 16773 14297 16807 14331
rect 16221 14229 16255 14263
rect 17877 14229 17911 14263
rect 38209 14229 38243 14263
rect 67741 14229 67775 14263
rect 18061 14025 18095 14059
rect 67281 14025 67315 14059
rect 14657 13957 14691 13991
rect 38117 13957 38151 13991
rect 39129 13957 39163 13991
rect 14013 13821 14047 13855
rect 15209 13821 15243 13855
rect 15853 13821 15887 13855
rect 16313 13821 16347 13855
rect 17049 13821 17083 13855
rect 17601 13821 17635 13855
rect 38669 13821 38703 13855
rect 39773 13821 39807 13855
rect 67925 13821 67959 13855
rect 68109 13821 68143 13855
rect 1869 13481 1903 13515
rect 12265 13481 12299 13515
rect 21373 13481 21407 13515
rect 1961 13413 1995 13447
rect 21373 13345 21407 13379
rect 14933 13277 14967 13311
rect 37381 13277 37415 13311
rect 38669 13277 38703 13311
rect 40969 13277 41003 13311
rect 2697 13209 2731 13243
rect 15669 13209 15703 13243
rect 18245 13209 18279 13243
rect 13553 13141 13587 13175
rect 16129 13141 16163 13175
rect 16773 13141 16807 13175
rect 17601 13141 17635 13175
rect 2237 12937 2271 12971
rect 14749 12937 14783 12971
rect 17233 12937 17267 12971
rect 37933 13141 37967 13175
rect 39221 13141 39255 13175
rect 39773 13141 39807 13175
rect 40417 13141 40451 13175
rect 41613 13141 41647 13175
rect 39037 12937 39071 12971
rect 40141 12937 40175 12971
rect 53849 12937 53883 12971
rect 15761 12869 15795 12903
rect 37381 12869 37415 12903
rect 16221 12733 16255 12767
rect 41429 12733 41463 12767
rect 14105 12665 14139 12699
rect 15209 12665 15243 12699
rect 15577 12665 15611 12699
rect 38485 12665 38519 12699
rect 41981 12665 42015 12699
rect 12265 12597 12299 12631
rect 12817 12597 12851 12631
rect 13369 12597 13403 12631
rect 15393 12597 15427 12631
rect 15485 12597 15519 12631
rect 17693 12597 17727 12631
rect 37933 12597 37967 12631
rect 39589 12597 39623 12631
rect 40877 12597 40911 12631
rect 12633 12325 12667 12359
rect 16589 12325 16623 12359
rect 18245 12257 18279 12291
rect 67465 12257 67499 12291
rect 68109 12257 68143 12291
rect 13277 12189 13311 12223
rect 16129 12189 16163 12223
rect 17969 12189 18003 12223
rect 41521 12189 41555 12223
rect 42073 12121 42107 12155
rect 11161 12053 11195 12087
rect 12081 12053 12115 12087
rect 13829 12053 13863 12087
rect 14657 12053 14691 12087
rect 15209 12053 15243 12087
rect 38117 12053 38151 12087
rect 38669 12053 38703 12087
rect 39129 12053 39163 12087
rect 39773 12053 39807 12087
rect 40417 12053 40451 12087
rect 40969 12053 41003 12087
rect 42717 12053 42751 12087
rect 43269 12053 43303 12087
rect 48053 12053 48087 12087
rect 38025 11849 38059 11883
rect 41981 11849 42015 11883
rect 38117 11645 38151 11679
rect 39129 11645 39163 11679
rect 10701 11577 10735 11611
rect 43545 11577 43579 11611
rect 44189 11577 44223 11611
rect 10149 11509 10183 11543
rect 12173 11509 12207 11543
rect 12817 11509 12851 11543
rect 13369 11509 13403 11543
rect 14473 11509 14507 11543
rect 14933 11509 14967 11543
rect 15577 11509 15611 11543
rect 16221 11509 16255 11543
rect 16957 11509 16991 11543
rect 17693 11509 17727 11543
rect 18153 11509 18187 11543
rect 38669 11509 38703 11543
rect 39773 11509 39807 11543
rect 40417 11509 40451 11543
rect 41061 11509 41095 11543
rect 42993 11509 43027 11543
rect 44649 11509 44683 11543
rect 66085 11509 66119 11543
rect 66637 11509 66671 11543
rect 67189 11509 67223 11543
rect 67649 11509 67683 11543
rect 67281 11305 67315 11339
rect 67925 11237 67959 11271
rect 1593 11169 1627 11203
rect 2053 11169 2087 11203
rect 9505 11169 9539 11203
rect 11529 11169 11563 11203
rect 37933 11169 37967 11203
rect 48329 11169 48363 11203
rect 10057 11101 10091 11135
rect 44281 11101 44315 11135
rect 65533 11101 65567 11135
rect 10885 11033 10919 11067
rect 11989 11033 12023 11067
rect 12633 11033 12667 11067
rect 13369 11033 13403 11067
rect 14381 11033 14415 11067
rect 15301 11033 15335 11067
rect 15853 11033 15887 11067
rect 16589 11033 16623 11067
rect 17141 11033 17175 11067
rect 17785 11033 17819 11067
rect 38669 11033 38703 11067
rect 39129 11033 39163 11067
rect 39773 11033 39807 11067
rect 40417 11033 40451 11067
rect 40969 11033 41003 11067
rect 41521 11033 41555 11067
rect 42073 11033 42107 11067
rect 42625 11033 42659 11067
rect 43177 11033 43211 11067
rect 43821 11033 43855 11067
rect 44833 11033 44867 11067
rect 45661 11033 45695 11067
rect 66085 11033 66119 11067
rect 66821 11033 66855 11067
rect 68109 11033 68143 11067
rect 17509 10761 17543 10795
rect 18245 10761 18279 10795
rect 10057 10693 10091 10727
rect 4353 10625 4387 10659
rect 4905 10625 4939 10659
rect 45753 10625 45787 10659
rect 10609 10557 10643 10591
rect 37933 10557 37967 10591
rect 45201 10557 45235 10591
rect 67005 10557 67039 10591
rect 9413 10489 9447 10523
rect 12265 10489 12299 10523
rect 39129 10489 39163 10523
rect 46305 10489 46339 10523
rect 66177 10489 66211 10523
rect 8861 10421 8895 10455
rect 11161 10421 11195 10455
rect 11713 10421 11747 10455
rect 13185 10421 13219 10455
rect 13921 10421 13955 10455
rect 14565 10421 14599 10455
rect 15301 10421 15335 10455
rect 16129 10421 16163 10455
rect 38669 10421 38703 10455
rect 39681 10421 39715 10455
rect 40233 10421 40267 10455
rect 40785 10421 40819 10455
rect 41429 10421 41463 10455
rect 41889 10421 41923 10455
rect 42993 10421 43027 10455
rect 43545 10421 43579 10455
rect 44189 10421 44223 10455
rect 44741 10421 44775 10455
rect 46949 10421 46983 10455
rect 47501 10421 47535 10455
rect 64797 10421 64831 10455
rect 65625 10421 65659 10455
rect 67465 10421 67499 10455
rect 68017 10421 68051 10455
rect 2237 10217 2271 10251
rect 9229 10217 9263 10251
rect 45753 10217 45787 10251
rect 13829 10149 13863 10183
rect 14749 10149 14783 10183
rect 67925 10149 67959 10183
rect 15209 10081 15243 10115
rect 18245 10081 18279 10115
rect 37933 10081 37967 10115
rect 38577 10081 38611 10115
rect 44097 10081 44131 10115
rect 8033 10013 8067 10047
rect 13001 9945 13035 9979
rect 17049 9945 17083 9979
rect 47317 9945 47351 9979
rect 66085 9945 66119 9979
rect 68109 9945 68143 9979
rect 2789 9877 2823 9911
rect 3893 9877 3927 9911
rect 4721 9877 4755 9911
rect 5365 9877 5399 9911
rect 6561 9877 6595 9911
rect 7205 9877 7239 9911
rect 8585 9877 8619 9911
rect 9781 9877 9815 9911
rect 10333 9877 10367 9911
rect 10885 9877 10919 9911
rect 11897 9877 11931 9911
rect 12449 9877 12483 9911
rect 15853 9877 15887 9911
rect 16497 9877 16531 9911
rect 17601 9877 17635 9911
rect 39221 9877 39255 9911
rect 39773 9877 39807 9911
rect 40601 9877 40635 9911
rect 41153 9877 41187 9911
rect 41705 9877 41739 9911
rect 42257 9877 42291 9911
rect 42809 9877 42843 9911
rect 43361 9877 43395 9911
rect 44833 9877 44867 9911
rect 46305 9877 46339 9911
rect 46765 9877 46799 9911
rect 47869 9877 47903 9911
rect 63969 9877 64003 9911
rect 64889 9877 64923 9911
rect 65441 9877 65475 9911
rect 67005 9877 67039 9911
rect 1777 9605 1811 9639
rect 2605 9605 2639 9639
rect 4537 9605 4571 9639
rect 18061 9605 18095 9639
rect 10609 9537 10643 9571
rect 34069 9537 34103 9571
rect 47593 9537 47627 9571
rect 1961 9469 1995 9503
rect 3729 9469 3763 9503
rect 3985 9469 4019 9503
rect 5641 9469 5675 9503
rect 8953 9469 8987 9503
rect 11161 9469 11195 9503
rect 14013 9469 14047 9503
rect 16405 9469 16439 9503
rect 17601 9469 17635 9503
rect 7389 9401 7423 9435
rect 15301 9401 15335 9435
rect 31493 9401 31527 9435
rect 5089 9333 5123 9367
rect 6469 9333 6503 9367
rect 7849 9333 7883 9367
rect 8493 9333 8527 9367
rect 9597 9333 9631 9367
rect 12081 9333 12115 9367
rect 12817 9333 12851 9367
rect 13369 9333 13403 9367
rect 14749 9333 14783 9367
rect 15853 9333 15887 9367
rect 7481 9129 7515 9163
rect 13645 8993 13679 9027
rect 14749 8993 14783 9027
rect 15393 8993 15427 9027
rect 17601 8993 17635 9027
rect 12449 8925 12483 8959
rect 4445 8857 4479 8891
rect 11897 8857 11931 8891
rect 16957 8857 16991 8891
rect 1409 8789 1443 8823
rect 1961 8789 1995 8823
rect 2513 8789 2547 8823
rect 3249 8789 3283 8823
rect 3985 8789 4019 8823
rect 5365 8789 5399 8823
rect 6101 8789 6135 8823
rect 7021 8789 7055 8823
rect 8309 8789 8343 8823
rect 9137 8789 9171 8823
rect 10057 8789 10091 8823
rect 10701 8789 10735 8823
rect 11161 8789 11195 8823
rect 13001 8789 13035 8823
rect 16405 8789 16439 8823
rect 18245 8789 18279 8823
rect 4445 8585 4479 8619
rect 6929 8585 6963 8619
rect 15025 8585 15059 8619
rect 15393 8585 15427 8619
rect 3157 8517 3191 8551
rect 14914 8517 14948 8551
rect 12541 8449 12575 8483
rect 15117 8449 15151 8483
rect 1777 8381 1811 8415
rect 2697 8381 2731 8415
rect 13185 8381 13219 8415
rect 14289 8381 14323 8415
rect 14749 8381 14783 8415
rect 16405 8381 16439 8415
rect 17509 8381 17543 8415
rect 18153 8381 18187 8415
rect 1961 8313 1995 8347
rect 3709 8313 3743 8347
rect 5549 8313 5583 8347
rect 7481 8313 7515 8347
rect 8125 8313 8159 8347
rect 9321 8313 9355 8347
rect 9965 8313 9999 8347
rect 10793 8313 10827 8347
rect 4905 8245 4939 8279
rect 8769 8245 8803 8279
rect 11989 8245 12023 8279
rect 6285 8041 6319 8075
rect 11069 7905 11103 7939
rect 11897 7905 11931 7939
rect 12541 7905 12575 7939
rect 13001 7905 13035 7939
rect 13829 7905 13863 7939
rect 15393 7905 15427 7939
rect 16037 7905 16071 7939
rect 16681 7905 16715 7939
rect 17141 7905 17175 7939
rect 18245 7905 18279 7939
rect 2789 7769 2823 7803
rect 1501 7701 1535 7735
rect 1961 7701 1995 7735
rect 3249 7701 3283 7735
rect 3893 7701 3927 7735
rect 4537 7701 4571 7735
rect 5181 7701 5215 7735
rect 5733 7701 5767 7735
rect 6929 7701 6963 7735
rect 7573 7701 7607 7735
rect 8309 7701 8343 7735
rect 9137 7701 9171 7735
rect 9689 7701 9723 7735
rect 10425 7701 10459 7735
rect 14749 7701 14783 7735
rect 4169 7497 4203 7531
rect 6929 7497 6963 7531
rect 2605 7361 2639 7395
rect 2881 7361 2915 7395
rect 9137 7361 9171 7395
rect 1593 7293 1627 7327
rect 7113 7293 7147 7327
rect 7389 7293 7423 7327
rect 10885 7293 10919 7327
rect 12265 7293 12299 7327
rect 13093 7293 13127 7327
rect 13553 7293 13587 7327
rect 14473 7293 14507 7327
rect 15117 7293 15151 7327
rect 15761 7293 15795 7327
rect 16405 7293 16439 7327
rect 17601 7293 17635 7327
rect 18245 7293 18279 7327
rect 7297 7225 7331 7259
rect 9689 7225 9723 7259
rect 2145 7157 2179 7191
rect 4721 7157 4755 7191
rect 5365 7157 5399 7191
rect 5825 7157 5859 7191
rect 8033 7157 8067 7191
rect 10241 7157 10275 7191
rect 1593 6817 1627 6851
rect 2053 6817 2087 6851
rect 10241 6817 10275 6851
rect 11161 6817 11195 6851
rect 11805 6817 11839 6851
rect 12449 6817 12483 6851
rect 12909 6817 12943 6851
rect 13829 6817 13863 6851
rect 15393 6817 15427 6851
rect 16037 6817 16071 6851
rect 16957 6817 16991 6851
rect 17601 6817 17635 6851
rect 18245 6817 18279 6851
rect 4445 6681 4479 6715
rect 6193 6681 6227 6715
rect 2605 6613 2639 6647
rect 3157 6613 3191 6647
rect 3893 6613 3927 6647
rect 5089 6613 5123 6647
rect 5733 6613 5767 6647
rect 6929 6613 6963 6647
rect 7481 6613 7515 6647
rect 8217 6613 8251 6647
rect 9597 6613 9631 6647
rect 14749 6613 14783 6647
rect 1409 6205 1443 6239
rect 2053 6205 2087 6239
rect 3157 6205 3191 6239
rect 8585 6205 8619 6239
rect 9413 6205 9447 6239
rect 9873 6205 9907 6239
rect 11161 6205 11195 6239
rect 12541 6205 12575 6239
rect 13185 6205 13219 6239
rect 13829 6205 13863 6239
rect 14473 6205 14507 6239
rect 15117 6205 15151 6239
rect 15761 6205 15795 6239
rect 16405 6205 16439 6239
rect 17601 6205 17635 6239
rect 18245 6205 18279 6239
rect 4261 6137 4295 6171
rect 7389 6137 7423 6171
rect 3617 6069 3651 6103
rect 4721 6069 4755 6103
rect 5273 6069 5307 6103
rect 5825 6069 5859 6103
rect 6745 6069 6779 6103
rect 7941 6069 7975 6103
rect 11897 6069 11931 6103
rect 1777 5797 1811 5831
rect 1961 5797 1995 5831
rect 2697 5729 2731 5763
rect 3341 5729 3375 5763
rect 5089 5729 5123 5763
rect 5733 5729 5767 5763
rect 8401 5729 8435 5763
rect 10149 5729 10183 5763
rect 10793 5729 10827 5763
rect 11897 5729 11931 5763
rect 12541 5729 12575 5763
rect 13185 5729 13219 5763
rect 13829 5729 13863 5763
rect 14933 5729 14967 5763
rect 15393 5729 15427 5763
rect 16313 5729 16347 5763
rect 16957 5729 16991 5763
rect 17601 5729 17635 5763
rect 9505 5661 9539 5695
rect 7389 5593 7423 5627
rect 3893 5525 3927 5559
rect 6285 5525 6319 5559
rect 6837 5525 6871 5559
rect 7941 5525 7975 5559
rect 18061 5525 18095 5559
rect 24501 5525 24535 5559
rect 1409 5117 1443 5151
rect 2053 5117 2087 5151
rect 2881 5117 2915 5151
rect 3525 5117 3559 5151
rect 4169 5117 4203 5151
rect 4813 5117 4847 5151
rect 5457 5117 5491 5151
rect 6837 5117 6871 5151
rect 7573 5117 7607 5151
rect 8217 5117 8251 5151
rect 9045 5117 9079 5151
rect 9505 5117 9539 5151
rect 10149 5117 10183 5151
rect 11161 5117 11195 5151
rect 12725 5117 12759 5151
rect 13369 5117 13403 5151
rect 14013 5117 14047 5151
rect 15393 5117 15427 5151
rect 16405 5117 16439 5151
rect 17877 5117 17911 5151
rect 12081 5049 12115 5083
rect 14473 5049 14507 5083
rect 14657 5049 14691 5083
rect 16957 5049 16991 5083
rect 17693 5049 17727 5083
rect 24501 4845 24535 4879
rect 25237 5525 25271 5559
rect 1961 4709 1995 4743
rect 14933 4709 14967 4743
rect 2697 4641 2731 4675
rect 3157 4641 3191 4675
rect 4629 4641 4663 4675
rect 5273 4641 5307 4675
rect 5733 4641 5767 4675
rect 6377 4641 6411 4675
rect 7021 4641 7055 4675
rect 7665 4641 7699 4675
rect 8585 4641 8619 4675
rect 9689 4641 9723 4675
rect 10609 4641 10643 4675
rect 11253 4641 11287 4675
rect 11897 4641 11931 4675
rect 12541 4641 12575 4675
rect 13185 4641 13219 4675
rect 13829 4641 13863 4675
rect 15669 4641 15703 4675
rect 16405 4641 16439 4675
rect 17049 4641 17083 4675
rect 18061 4641 18095 4675
rect 14749 4505 14783 4539
rect 15485 4505 15519 4539
rect 16865 4505 16899 4539
rect 18245 4505 18279 4539
rect 1869 4437 1903 4471
rect 3893 4437 3927 4471
rect 19257 4437 19291 4471
rect 5917 4165 5951 4199
rect 19073 4097 19107 4131
rect 1593 4029 1627 4063
rect 2697 4029 2731 4063
rect 3341 4029 3375 4063
rect 3801 4029 3835 4063
rect 5181 4029 5215 4063
rect 6837 4029 6871 4063
rect 7481 4029 7515 4063
rect 8401 4029 8435 4063
rect 9045 4029 9079 4063
rect 9873 4029 9907 4063
rect 10517 4029 10551 4063
rect 11161 4029 11195 4063
rect 13001 4029 13035 4063
rect 15393 4029 15427 4063
rect 16221 4029 16255 4063
rect 17509 4029 17543 4063
rect 18061 4029 18095 4063
rect 4997 3961 5031 3995
rect 12081 3961 12115 3995
rect 12265 3961 12299 3995
rect 12817 3961 12851 3995
rect 13553 3961 13587 3995
rect 13737 3961 13771 3995
rect 14473 3961 14507 3995
rect 16037 3961 16071 3995
rect 18245 3961 18279 3995
rect 4537 3893 4571 3927
rect 14381 3893 14415 3927
rect 15485 3893 15519 3927
rect 10609 3689 10643 3723
rect 14565 3689 14599 3723
rect 4445 3621 4479 3655
rect 5641 3621 5675 3655
rect 6377 3621 6411 3655
rect 9321 3621 9355 3655
rect 12633 3621 12667 3655
rect 13369 3621 13403 3655
rect 15301 3621 15335 3655
rect 15853 3621 15887 3655
rect 16589 3621 16623 3655
rect 18061 3621 18095 3655
rect 1593 3553 1627 3587
rect 2237 3553 2271 3587
rect 2881 3553 2915 3587
rect 6929 3553 6963 3587
rect 7573 3553 7607 3587
rect 8217 3553 8251 3587
rect 9965 3553 9999 3587
rect 11722 3553 11756 3587
rect 15117 3553 15151 3587
rect 17325 3553 17359 3587
rect 18245 3553 18279 3587
rect 11989 3485 12023 3519
rect 12449 3485 12483 3519
rect 16773 3485 16807 3519
rect 4261 3417 4295 3451
rect 5457 3417 5491 3451
rect 16037 3417 16071 3451
rect 6285 3349 6319 3383
rect 9873 3349 9907 3383
rect 13277 3349 13311 3383
rect 17417 3349 17451 3383
rect 2513 3145 2547 3179
rect 5641 3145 5675 3179
rect 19165 4029 19199 4063
rect 19165 3145 19199 3179
rect 4813 3077 4847 3111
rect 14197 3077 14231 3111
rect 16405 3077 16439 3111
rect 19073 3077 19107 3111
rect 4077 3009 4111 3043
rect 10701 3009 10735 3043
rect 3341 2941 3375 2975
rect 3525 2941 3559 2975
rect 4997 2941 5031 2975
rect 6837 2941 6871 2975
rect 7021 2941 7055 2975
rect 8033 2941 8067 2975
rect 8677 2941 8711 2975
rect 9965 2941 9999 2975
rect 12081 2941 12115 2975
rect 13001 2941 13035 2975
rect 14013 2941 14047 2975
rect 14749 2941 14783 2975
rect 15577 2941 15611 2975
rect 16221 2941 16255 2975
rect 17509 2941 17543 2975
rect 1961 2873 1995 2907
rect 2513 2873 2547 2907
rect 2789 2873 2823 2907
rect 4261 2873 4295 2907
rect 5733 2873 5767 2907
rect 8493 2873 8527 2907
rect 9229 2873 9263 2907
rect 9413 2873 9447 2907
rect 10149 2873 10183 2907
rect 10885 2873 10919 2907
rect 12265 2873 12299 2907
rect 14933 2873 14967 2907
rect 18061 2873 18095 2907
rect 18245 2873 18279 2907
rect 1869 2805 1903 2839
rect 2697 2805 2731 2839
rect 12909 2805 12943 2839
rect 15485 2805 15519 2839
rect 15945 2601 15979 2635
rect 16589 2601 16623 2635
rect 19165 2601 19199 2635
rect 4997 2533 5031 2567
rect 5181 2533 5215 2567
rect 5917 2533 5951 2567
rect 7113 2533 7147 2567
rect 7849 2533 7883 2567
rect 8585 2533 8619 2567
rect 9781 2533 9815 2567
rect 10517 2533 10551 2567
rect 12357 2533 12391 2567
rect 13093 2533 13127 2567
rect 13829 2533 13863 2567
rect 15301 2533 15335 2567
rect 16497 2533 16531 2567
rect 18061 2533 18095 2567
rect 1501 2465 1535 2499
rect 4445 2465 4479 2499
rect 9597 2465 9631 2499
rect 11161 2465 11195 2499
rect 11345 2465 11379 2499
rect 14657 2465 14691 2499
rect 2053 2397 2087 2431
rect 2605 2397 2639 2431
rect 3249 2397 3283 2431
rect 4261 2329 4295 2363
rect 6929 2329 6963 2363
rect 8401 2329 8435 2363
rect 12541 2329 12575 2363
rect 15117 2329 15151 2363
rect 5825 2261 5859 2295
rect 7757 2261 7791 2295
rect 10425 2261 10459 2295
rect 13185 2261 13219 2295
rect 13921 2261 13955 2295
rect 17509 2261 17543 2295
rect 18153 2261 18187 2295
rect 22937 3689 22971 3723
rect 22569 3553 22603 3587
rect 20729 3485 20763 3519
rect 20729 3145 20763 3179
rect 21741 3213 21775 3247
rect 21741 2873 21775 2907
rect 22109 3213 22143 3247
rect 19257 2533 19291 2567
rect 22109 1921 22143 1955
rect 22477 3077 22511 3111
rect 19165 1785 19199 1819
rect 22569 2669 22603 2703
rect 23397 2805 23431 2839
rect 23397 2669 23431 2703
rect 22937 2125 22971 2159
rect 28641 4505 28675 4539
rect 26893 4029 26927 4063
rect 26525 3757 26559 3791
rect 25881 3417 25915 3451
rect 25789 3281 25823 3315
rect 25329 2941 25363 2975
rect 25329 1853 25363 1887
rect 25605 2805 25639 2839
rect 25605 1853 25639 1887
rect 25789 1853 25823 1887
rect 26341 3145 26375 3179
rect 25881 1853 25915 1887
rect 26065 3077 26099 3111
rect 26341 1921 26375 1955
rect 26525 1921 26559 1955
rect 26617 3009 26651 3043
rect 26617 1921 26651 1955
rect 26801 2873 26835 2907
rect 26065 1853 26099 1887
rect 27905 3893 27939 3927
rect 26893 1921 26927 1955
rect 27169 3621 27203 3655
rect 27169 1921 27203 1955
rect 27353 3621 27387 3655
rect 26801 1853 26835 1887
rect 27445 3281 27479 3315
rect 27445 1921 27479 1955
rect 27629 2805 27663 2839
rect 27629 1921 27663 1955
rect 27905 1921 27939 1955
rect 27353 1853 27387 1887
rect 25237 1785 25271 1819
rect 30573 4097 30607 4131
rect 29009 3961 29043 3995
rect 28733 3689 28767 3723
rect 28733 1921 28767 1955
rect 30297 3825 30331 3859
rect 29009 1921 29043 1955
rect 29193 3349 29227 3383
rect 29193 1921 29227 1955
rect 29469 3145 29503 3179
rect 28641 1717 28675 1751
rect 29561 3077 29595 3111
rect 29561 1717 29595 1751
rect 29469 1513 29503 1547
rect 30297 1513 30331 1547
rect 30481 3417 30515 3451
rect 22477 1445 22511 1479
rect 31125 3757 31159 3791
rect 30849 3553 30883 3587
rect 30573 1513 30607 1547
rect 30757 3485 30791 3519
rect 30481 1309 30515 1343
rect 30941 1989 30975 2023
rect 30941 1649 30975 1683
rect 31125 1649 31159 1683
rect 31309 2873 31343 2907
rect 31309 1649 31343 1683
rect 30849 1513 30883 1547
rect 33609 8517 33643 8551
rect 31585 6205 31619 6239
rect 31953 5593 31987 5627
rect 31769 5525 31803 5559
rect 31769 4845 31803 4879
rect 32045 5525 32079 5559
rect 32045 4845 32079 4879
rect 32321 5525 32355 5559
rect 32321 4845 32355 4879
rect 32505 5525 32539 5559
rect 32505 4845 32539 4879
rect 32965 5185 32999 5219
rect 31953 4641 31987 4675
rect 31585 3621 31619 3655
rect 32689 4165 32723 4199
rect 32689 3485 32723 3519
rect 31585 3213 31619 3247
rect 33425 5049 33459 5083
rect 32137 2805 32171 2839
rect 32321 2805 32355 2839
rect 32965 2805 32999 2839
rect 33333 3757 33367 3791
rect 33333 2669 33367 2703
rect 33425 2533 33459 2567
rect 33885 3689 33919 3723
rect 33885 3077 33919 3111
rect 33977 3213 34011 3247
rect 33977 2533 34011 2567
rect 33609 2329 33643 2363
rect 31585 1649 31619 1683
rect 31493 1513 31527 1547
rect 30757 1309 30791 1343
rect 37933 9469 37967 9503
rect 38761 9469 38795 9503
rect 39405 9469 39439 9503
rect 40049 9469 40083 9503
rect 40969 9469 41003 9503
rect 43085 9469 43119 9503
rect 44189 9401 44223 9435
rect 47041 9401 47075 9435
rect 48697 9401 48731 9435
rect 65717 9401 65751 9435
rect 41521 9333 41555 9367
rect 42073 9333 42107 9367
rect 43545 9333 43579 9367
rect 44741 9333 44775 9367
rect 45201 9333 45235 9367
rect 45845 9333 45879 9367
rect 46581 9333 46615 9367
rect 49157 9333 49191 9367
rect 49709 9333 49743 9367
rect 50261 9333 50295 9367
rect 63325 9333 63359 9367
rect 63969 9333 64003 9367
rect 64521 9333 64555 9367
rect 65165 9333 65199 9367
rect 66269 9333 66303 9367
rect 66729 9333 66763 9367
rect 67649 9333 67683 9367
rect 64521 9129 64555 9163
rect 50905 9061 50939 9095
rect 38117 8993 38151 9027
rect 38945 8993 38979 9027
rect 39589 8993 39623 9027
rect 41153 8993 41187 9027
rect 68109 8993 68143 9027
rect 48973 8925 49007 8959
rect 62405 8857 62439 8891
rect 66913 8857 66947 8891
rect 40417 8789 40451 8823
rect 41797 8789 41831 8823
rect 42349 8789 42383 8823
rect 42901 8789 42935 8823
rect 43453 8789 43487 8823
rect 44005 8789 44039 8823
rect 44557 8789 44591 8823
rect 45661 8789 45695 8823
rect 46213 8789 46247 8823
rect 46765 8789 46799 8823
rect 47317 8789 47351 8823
rect 47869 8789 47903 8823
rect 48421 8789 48455 8823
rect 49617 8789 49651 8823
rect 50169 8789 50203 8823
rect 51549 8789 51583 8823
rect 52009 8789 52043 8823
rect 52561 8789 52595 8823
rect 53205 8789 53239 8823
rect 54125 8789 54159 8823
rect 62957 8789 62991 8823
rect 63509 8789 63543 8823
rect 64061 8789 64095 8823
rect 65073 8789 65107 8823
rect 65717 8789 65751 8823
rect 67465 8789 67499 8823
rect 34437 8585 34471 8619
rect 50353 8585 50387 8619
rect 50813 8585 50847 8619
rect 51549 8585 51583 8619
rect 52009 8585 52043 8619
rect 54125 8585 54159 8619
rect 61393 8585 61427 8619
rect 34345 4437 34379 4471
rect 34161 3689 34195 3723
rect 34161 1921 34195 1955
rect 38117 8381 38151 8415
rect 38761 8381 38795 8415
rect 39405 8381 39439 8415
rect 40049 8381 40083 8415
rect 40509 8381 40543 8415
rect 41429 8381 41463 8415
rect 42257 8381 42291 8415
rect 43545 8381 43579 8415
rect 44649 8381 44683 8415
rect 66269 8381 66303 8415
rect 67465 8381 67499 8415
rect 68109 8381 68143 8415
rect 45753 8313 45787 8347
rect 46765 8313 46799 8347
rect 47317 8313 47351 8347
rect 48329 8313 48363 8347
rect 48789 8313 48823 8347
rect 49341 8313 49375 8347
rect 52561 8313 52595 8347
rect 53481 8313 53515 8347
rect 54677 8313 54711 8347
rect 55229 8313 55263 8347
rect 55689 8313 55723 8347
rect 62221 8313 62255 8347
rect 62957 8313 62991 8347
rect 64521 8313 64555 8347
rect 65625 8313 65659 8347
rect 66729 8313 66763 8347
rect 44005 8245 44039 8279
rect 45201 8245 45235 8279
rect 46213 8245 46247 8279
rect 64981 8245 65015 8279
rect 55321 8041 55355 8075
rect 56701 8041 56735 8075
rect 57345 8041 57379 8075
rect 57989 8041 58023 8075
rect 38117 7905 38151 7939
rect 38761 7905 38795 7939
rect 39405 7905 39439 7939
rect 40969 7905 41003 7939
rect 41613 7905 41647 7939
rect 42257 7905 42291 7939
rect 42901 7905 42935 7939
rect 43545 7905 43579 7939
rect 44005 7905 44039 7939
rect 44649 7905 44683 7939
rect 67373 7905 67407 7939
rect 68017 7905 68051 7939
rect 37473 7837 37507 7871
rect 48973 7837 49007 7871
rect 37381 6817 37415 6851
rect 37381 6205 37415 6239
rect 34989 5185 35023 5219
rect 34989 4505 35023 4539
rect 35817 4029 35851 4063
rect 35725 3893 35759 3927
rect 34897 3485 34931 3519
rect 34989 3485 35023 3519
rect 34989 3349 35023 3383
rect 35817 3621 35851 3655
rect 37289 3961 37323 3995
rect 49525 7769 49559 7803
rect 63693 7769 63727 7803
rect 65441 7769 65475 7803
rect 45661 7701 45695 7735
rect 46213 7701 46247 7735
rect 46857 7701 46891 7735
rect 47317 7701 47351 7735
rect 47869 7701 47903 7735
rect 48421 7701 48455 7735
rect 50169 7701 50203 7735
rect 50905 7701 50939 7735
rect 51457 7701 51491 7735
rect 52101 7701 52135 7735
rect 52561 7701 52595 7735
rect 53113 7701 53147 7735
rect 53665 7701 53699 7735
rect 54585 7701 54619 7735
rect 56149 7701 56183 7735
rect 60841 7701 60875 7735
rect 61945 7701 61979 7735
rect 62497 7701 62531 7735
rect 63049 7701 63083 7735
rect 64153 7701 64187 7735
rect 64889 7701 64923 7735
rect 65901 7701 65935 7735
rect 66637 7701 66671 7735
rect 56793 7497 56827 7531
rect 57437 7497 57471 7531
rect 57989 7497 58023 7531
rect 60197 7497 60231 7531
rect 60749 7497 60783 7531
rect 61669 7497 61703 7531
rect 38117 7293 38151 7327
rect 38761 7293 38795 7327
rect 39405 7293 39439 7327
rect 40049 7293 40083 7327
rect 40785 7293 40819 7327
rect 41429 7293 41463 7327
rect 42257 7293 42291 7327
rect 43361 7293 43395 7327
rect 44189 7293 44223 7327
rect 44833 7293 44867 7327
rect 45477 7293 45511 7327
rect 47133 7293 47167 7327
rect 50997 7293 51031 7327
rect 65441 7293 65475 7327
rect 66085 7293 66119 7327
rect 66729 7293 66763 7327
rect 67189 7293 67223 7327
rect 67925 7293 67959 7327
rect 51549 7225 51583 7259
rect 52653 7225 52687 7259
rect 54585 7225 54619 7259
rect 68109 7225 68143 7259
rect 45937 7157 45971 7191
rect 46489 7157 46523 7191
rect 47593 7157 47627 7191
rect 48237 7157 48271 7191
rect 48881 7157 48915 7191
rect 49341 7157 49375 7191
rect 49893 7157 49927 7191
rect 50537 7157 50571 7191
rect 52193 7157 52227 7191
rect 53481 7157 53515 7191
rect 54033 7157 54067 7191
rect 55229 7157 55263 7191
rect 55689 7157 55723 7191
rect 56241 7157 56275 7191
rect 59645 7157 59679 7191
rect 62313 7157 62347 7191
rect 62773 7157 62807 7191
rect 63325 7157 63359 7191
rect 63969 7157 64003 7191
rect 64797 7157 64831 7191
rect 38117 6817 38151 6851
rect 38577 6817 38611 6851
rect 39405 6817 39439 6851
rect 41337 6817 41371 6851
rect 42165 6817 42199 6851
rect 42809 6817 42843 6851
rect 43545 6817 43579 6851
rect 44005 6817 44039 6851
rect 44833 6817 44867 6851
rect 46029 6817 46063 6851
rect 46673 6817 46707 6851
rect 47501 6817 47535 6851
rect 59369 6817 59403 6851
rect 64981 6817 65015 6851
rect 65625 6817 65659 6851
rect 67465 6817 67499 6851
rect 67925 6817 67959 6851
rect 48513 6749 48547 6783
rect 49065 6681 49099 6715
rect 58357 6681 58391 6715
rect 40417 6613 40451 6647
rect 47961 6613 47995 6647
rect 49709 6613 49743 6647
rect 50169 6613 50203 6647
rect 50905 6613 50939 6647
rect 51457 6613 51491 6647
rect 52009 6613 52043 6647
rect 52561 6613 52595 6647
rect 53205 6613 53239 6647
rect 53941 6613 53975 6647
rect 54585 6613 54619 6647
rect 55045 6613 55079 6647
rect 56149 6613 56183 6647
rect 56701 6613 56735 6647
rect 57253 6613 57287 6647
rect 57897 6613 57931 6647
rect 59921 6613 59955 6647
rect 60381 6613 60415 6647
rect 61393 6613 61427 6647
rect 62037 6613 62071 6647
rect 62865 6613 62899 6647
rect 63417 6613 63451 6647
rect 64153 6613 64187 6647
rect 66821 6613 66855 6647
rect 39589 6409 39623 6443
rect 40049 6409 40083 6443
rect 37933 6273 37967 6307
rect 38761 6273 38795 6307
rect 48789 6273 48823 6307
rect 40693 6205 40727 6239
rect 41429 6205 41463 6239
rect 42073 6205 42107 6239
rect 43361 6205 43395 6239
rect 44005 6205 44039 6239
rect 44833 6205 44867 6239
rect 45477 6205 45511 6239
rect 46121 6205 46155 6239
rect 46765 6205 46799 6239
rect 47225 6205 47259 6239
rect 50261 6205 50295 6239
rect 50905 6205 50939 6239
rect 52009 6205 52043 6239
rect 64797 6205 64831 6239
rect 65257 6205 65291 6239
rect 66637 6205 66671 6239
rect 67097 6205 67131 6239
rect 68109 6205 68143 6239
rect 49341 6137 49375 6171
rect 58081 6137 58115 6171
rect 60749 6137 60783 6171
rect 48237 6069 48271 6103
rect 52561 6069 52595 6103
rect 53665 6069 53699 6103
rect 54401 6069 54435 6103
rect 55045 6069 55079 6103
rect 55597 6069 55631 6103
rect 56149 6069 56183 6103
rect 56977 6069 57011 6103
rect 57529 6069 57563 6103
rect 58909 6069 58943 6103
rect 59645 6069 59679 6103
rect 60105 6069 60139 6103
rect 61669 6069 61703 6103
rect 62313 6069 62347 6103
rect 62957 6069 62991 6103
rect 64061 6069 64095 6103
rect 65901 6069 65935 6103
rect 38485 5797 38519 5831
rect 67189 5797 67223 5831
rect 67925 5797 67959 5831
rect 39865 5729 39899 5763
rect 41061 5729 41095 5763
rect 41705 5729 41739 5763
rect 42349 5729 42383 5763
rect 42809 5729 42843 5763
rect 43637 5729 43671 5763
rect 44281 5729 44315 5763
rect 44925 5729 44959 5763
rect 46765 5729 46799 5763
rect 47225 5729 47259 5763
rect 48053 5729 48087 5763
rect 48697 5729 48731 5763
rect 49341 5729 49375 5763
rect 49985 5729 50019 5763
rect 51457 5729 51491 5763
rect 52101 5729 52135 5763
rect 52745 5729 52779 5763
rect 53205 5729 53239 5763
rect 54033 5729 54067 5763
rect 54677 5729 54711 5763
rect 55321 5729 55355 5763
rect 56701 5729 56735 5763
rect 62865 5729 62899 5763
rect 63509 5729 63543 5763
rect 64337 5729 64371 5763
rect 65441 5729 65475 5763
rect 66085 5729 66119 5763
rect 68109 5729 68143 5763
rect 38301 5593 38335 5627
rect 39221 5593 39255 5627
rect 60749 5593 60783 5627
rect 67373 5593 67407 5627
rect 45661 5525 45695 5559
rect 57161 5525 57195 5559
rect 57713 5525 57747 5559
rect 58817 5525 58851 5559
rect 59369 5525 59403 5559
rect 60289 5525 60323 5559
rect 61393 5525 61427 5559
rect 61945 5525 61979 5559
rect 39865 5321 39899 5355
rect 51181 5253 51215 5287
rect 49433 5185 49467 5219
rect 39221 5117 39255 5151
rect 41245 5117 41279 5151
rect 41429 5117 41463 5151
rect 42165 5117 42199 5151
rect 43545 5117 43579 5151
rect 44189 5117 44223 5151
rect 44649 5117 44683 5151
rect 45477 5117 45511 5151
rect 46121 5117 46155 5151
rect 46765 5117 46799 5151
rect 47409 5117 47443 5151
rect 48789 5117 48823 5151
rect 50077 5117 50111 5151
rect 51733 5117 51767 5151
rect 52193 5117 52227 5151
rect 54033 5117 54067 5151
rect 54493 5117 54527 5151
rect 55321 5117 55355 5151
rect 55965 5117 55999 5151
rect 56425 5117 56459 5151
rect 57253 5117 57287 5151
rect 57897 5117 57931 5151
rect 60105 5117 60139 5151
rect 60565 5117 60599 5151
rect 61393 5117 61427 5151
rect 61853 5117 61887 5151
rect 62681 5117 62715 5151
rect 63141 5117 63175 5151
rect 64337 5117 64371 5151
rect 65165 5117 65199 5151
rect 65809 5117 65843 5151
rect 66453 5117 66487 5151
rect 67925 5117 67959 5151
rect 38301 5049 38335 5083
rect 38485 5049 38519 5083
rect 39957 5049 39991 5083
rect 40693 5049 40727 5083
rect 51365 5049 51399 5083
rect 67189 5049 67223 5083
rect 68109 5049 68143 5083
rect 39129 4981 39163 5015
rect 40601 4981 40635 5015
rect 51457 4981 51491 5015
rect 51549 4981 51583 5015
rect 52837 4981 52871 5015
rect 58725 4981 58759 5015
rect 59369 4981 59403 5015
rect 67281 4981 67315 5015
rect 67189 4709 67223 4743
rect 68017 4709 68051 4743
rect 38485 4641 38519 4675
rect 39221 4641 39255 4675
rect 39865 4641 39899 4675
rect 40969 4641 41003 4675
rect 42165 4641 42199 4675
rect 42901 4641 42935 4675
rect 44741 4641 44775 4675
rect 46213 4641 46247 4675
rect 46673 4641 46707 4675
rect 47409 4641 47443 4675
rect 48053 4641 48087 4675
rect 48513 4641 48547 4675
rect 49157 4641 49191 4675
rect 49985 4641 50019 4675
rect 51457 4641 51491 4675
rect 52101 4641 52135 4675
rect 53389 4641 53423 4675
rect 54033 4641 54067 4675
rect 54677 4641 54711 4675
rect 55597 4641 55631 4675
rect 56885 4641 56919 4675
rect 57529 4641 57563 4675
rect 57989 4641 58023 4675
rect 58817 4641 58851 4675
rect 59737 4641 59771 4675
rect 62405 4641 62439 4675
rect 63233 4641 63267 4675
rect 64061 4641 64095 4675
rect 64705 4641 64739 4675
rect 65165 4641 65199 4675
rect 65993 4641 66027 4675
rect 44097 4573 44131 4607
rect 38301 4505 38335 4539
rect 40785 4505 40819 4539
rect 43361 4505 43395 4539
rect 61761 4505 61795 4539
rect 67833 4505 67867 4539
rect 39129 4437 39163 4471
rect 42073 4437 42107 4471
rect 52745 4437 52779 4471
rect 56241 4437 56275 4471
rect 60197 4437 60231 4471
rect 67281 4437 67315 4471
rect 39037 4165 39071 4199
rect 58081 4165 58115 4199
rect 41981 4097 42015 4131
rect 39221 4029 39255 4063
rect 39773 4029 39807 4063
rect 40693 4029 40727 4063
rect 42165 4029 42199 4063
rect 44649 4029 44683 4063
rect 45385 4029 45419 4063
rect 46029 4029 46063 4063
rect 46673 4029 46707 4063
rect 47317 4029 47351 4063
rect 48789 4029 48823 4063
rect 49249 4029 49283 4063
rect 49893 4029 49927 4063
rect 50721 4029 50755 4063
rect 51365 4029 51399 4063
rect 52009 4029 52043 4063
rect 52469 4029 52503 4063
rect 53849 4029 53883 4063
rect 54493 4029 54527 4063
rect 55137 4029 55171 4063
rect 55781 4029 55815 4063
rect 56609 4029 56643 4063
rect 57253 4029 57287 4063
rect 59093 4029 59127 4063
rect 59737 4029 59771 4063
rect 60657 4029 60691 4063
rect 61577 4029 61611 4063
rect 62773 4029 62807 4063
rect 63417 4029 63451 4063
rect 64337 4029 64371 4063
rect 65441 4029 65475 4063
rect 65993 4029 66027 4063
rect 66821 4029 66855 4063
rect 38301 3961 38335 3995
rect 38485 3961 38519 3995
rect 39957 3961 39991 3995
rect 41245 3961 41279 3995
rect 41429 3961 41463 3995
rect 43545 3961 43579 3995
rect 44465 3961 44499 3995
rect 66637 3961 66671 3995
rect 67465 3961 67499 3995
rect 67649 3961 67683 3995
rect 40601 3893 40635 3927
rect 43453 3893 43487 3927
rect 62037 3893 62071 3927
rect 66085 3893 66119 3927
rect 44925 3689 44959 3723
rect 37473 3621 37507 3655
rect 38485 3621 38519 3655
rect 40969 3621 41003 3655
rect 42165 3621 42199 3655
rect 42717 3621 42751 3655
rect 44373 3621 44407 3655
rect 45661 3621 45695 3655
rect 47685 3621 47719 3655
rect 52745 3621 52779 3655
rect 54493 3621 54527 3655
rect 55321 3621 55355 3655
rect 56701 3621 56735 3655
rect 57437 3621 57471 3655
rect 64245 3621 64279 3655
rect 65073 3621 65107 3655
rect 65901 3621 65935 3655
rect 67189 3621 67223 3655
rect 67925 3621 67959 3655
rect 39037 3553 39071 3587
rect 39221 3553 39255 3587
rect 42901 3553 42935 3587
rect 43637 3553 43671 3587
rect 46765 3553 46799 3587
rect 48237 3553 48271 3587
rect 48881 3553 48915 3587
rect 49709 3553 49743 3587
rect 50353 3553 50387 3587
rect 51457 3553 51491 3587
rect 51917 3553 51951 3587
rect 53573 3553 53607 3587
rect 58173 3553 58207 3587
rect 59001 3553 59035 3587
rect 59461 3553 59495 3587
rect 60289 3553 60323 3587
rect 61945 3553 61979 3587
rect 62405 3553 62439 3587
rect 63049 3553 63083 3587
rect 66085 3553 66119 3587
rect 37289 3485 37323 3519
rect 37381 3485 37415 3519
rect 41981 3485 42015 3519
rect 40785 3417 40819 3451
rect 43453 3417 43487 3451
rect 46581 3417 46615 3451
rect 47501 3417 47535 3451
rect 52561 3417 52595 3451
rect 53389 3417 53423 3451
rect 54309 3417 54343 3451
rect 55137 3417 55171 3451
rect 56517 3417 56551 3451
rect 57253 3417 57287 3451
rect 64061 3417 64095 3451
rect 64889 3417 64923 3451
rect 67741 3417 67775 3451
rect 38393 3349 38427 3383
rect 39773 3349 39807 3383
rect 44281 3349 44315 3383
rect 60749 3349 60783 3383
rect 67097 3349 67131 3383
rect 37381 3281 37415 3315
rect 34897 3145 34931 3179
rect 35633 3145 35667 3179
rect 35725 3145 35759 3179
rect 39129 3145 39163 3179
rect 44189 3145 44223 3179
rect 67281 3145 67315 3179
rect 39773 3077 39807 3111
rect 41245 3077 41279 3111
rect 68109 3077 68143 3111
rect 38301 3009 38335 3043
rect 40509 3009 40543 3043
rect 43361 3009 43395 3043
rect 45569 3009 45603 3043
rect 47041 3009 47075 3043
rect 51549 3009 51583 3043
rect 52285 3009 52319 3043
rect 54585 3009 54619 3043
rect 56057 3009 56091 3043
rect 61761 3009 61795 3043
rect 63417 3009 63451 3043
rect 38485 2941 38519 2975
rect 39221 2941 39255 2975
rect 39957 2941 39991 2975
rect 40693 2941 40727 2975
rect 41429 2941 41463 2975
rect 41981 2941 42015 2975
rect 43545 2941 43579 2975
rect 44281 2941 44315 2975
rect 46489 2941 46523 2975
rect 47225 2941 47259 2975
rect 48789 2941 48823 2975
rect 49341 2941 49375 2975
rect 50261 2941 50295 2975
rect 50997 2941 51031 2975
rect 52469 2941 52503 2975
rect 54033 2941 54067 2975
rect 54769 2941 54803 2975
rect 57529 2941 57563 2975
rect 59277 2941 59311 2975
rect 59921 2941 59955 2975
rect 60381 2941 60415 2975
rect 61209 2941 61243 2975
rect 62497 2941 62531 2975
rect 64521 2941 64555 2975
rect 65257 2941 65291 2975
rect 65993 2941 66027 2975
rect 66729 2941 66763 2975
rect 35725 2873 35759 2907
rect 42165 2873 42199 2907
rect 44833 2873 44867 2907
rect 45017 2873 45051 2907
rect 45753 2873 45787 2907
rect 48605 2873 48639 2907
rect 49525 2873 49559 2907
rect 50077 2873 50111 2907
rect 51733 2873 51767 2907
rect 53849 2873 53883 2907
rect 55505 2873 55539 2907
rect 56241 2873 56275 2907
rect 56977 2873 57011 2907
rect 57713 2873 57747 2907
rect 61025 2873 61059 2907
rect 62313 2873 62347 2907
rect 63233 2873 63267 2907
rect 64337 2873 64371 2907
rect 65073 2873 65107 2907
rect 65809 2873 65843 2907
rect 67925 2873 67959 2907
rect 36001 2805 36035 2839
rect 46397 2805 46431 2839
rect 50905 2805 50939 2839
rect 55413 2805 55447 2839
rect 56885 2805 56919 2839
rect 66637 2805 66671 2839
rect 34437 1921 34471 1955
rect 35449 2397 35483 2431
rect 35449 1785 35483 1819
rect 44281 2601 44315 2635
rect 49617 2601 49651 2635
rect 51549 2601 51583 2635
rect 54217 2601 54251 2635
rect 63693 2601 63727 2635
rect 39221 2533 39255 2567
rect 40969 2533 41003 2567
rect 42441 2533 42475 2567
rect 43637 2533 43671 2567
rect 44373 2533 44407 2567
rect 45109 2533 45143 2567
rect 46305 2533 46339 2567
rect 47041 2533 47075 2567
rect 47777 2533 47811 2567
rect 48789 2533 48823 2567
rect 48973 2533 49007 2567
rect 49709 2533 49743 2567
rect 50261 2533 50295 2567
rect 50445 2533 50479 2567
rect 51641 2533 51675 2567
rect 52929 2533 52963 2567
rect 53113 2533 53147 2567
rect 54309 2533 54343 2567
rect 54861 2533 54895 2567
rect 55045 2533 55079 2567
rect 55781 2533 55815 2567
rect 56977 2533 57011 2567
rect 57805 2533 57839 2567
rect 59645 2533 59679 2567
rect 60381 2533 60415 2567
rect 61117 2533 61151 2567
rect 62313 2533 62347 2567
rect 63785 2533 63819 2567
rect 64981 2533 65015 2567
rect 65717 2533 65751 2567
rect 66269 2533 66303 2567
rect 66453 2533 66487 2567
rect 67925 2533 67959 2567
rect 38485 2465 38519 2499
rect 41705 2465 41739 2499
rect 52193 2465 52227 2499
rect 52377 2465 52411 2499
rect 57161 2465 57195 2499
rect 58549 2465 58583 2499
rect 63049 2465 63083 2499
rect 67097 2465 67131 2499
rect 39037 2397 39071 2431
rect 39865 2397 39899 2431
rect 60933 2397 60967 2431
rect 62865 2397 62899 2431
rect 65533 2397 65567 2431
rect 37289 2329 37323 2363
rect 38301 2329 38335 2363
rect 40785 2329 40819 2363
rect 46857 2329 46891 2363
rect 55597 2329 55631 2363
rect 57621 2329 57655 2363
rect 59461 2329 59495 2363
rect 62129 2329 62163 2363
rect 64797 2329 64831 2363
rect 68109 2329 68143 2363
rect 41613 2261 41647 2295
rect 42349 2261 42383 2295
rect 43545 2261 43579 2295
rect 45017 2261 45051 2295
rect 46213 2261 46247 2295
rect 47685 2261 47719 2295
rect 60289 2261 60323 2295
rect 37289 1989 37323 2023
rect 39773 2057 39807 2091
rect 36461 1921 36495 1955
rect 36553 1853 36587 1887
rect 36553 1581 36587 1615
rect 36461 1445 36495 1479
rect 36001 1309 36035 1343
rect 34345 1241 34379 1275
rect 39773 1037 39807 1071
rect 34069 969 34103 1003
<< metal1 >>
rect 1104 67482 68816 67504
rect 1104 67430 4246 67482
rect 4298 67430 4310 67482
rect 4362 67430 4374 67482
rect 4426 67430 4438 67482
rect 4490 67430 14246 67482
rect 14298 67430 14310 67482
rect 14362 67430 14374 67482
rect 14426 67430 14438 67482
rect 14490 67430 24246 67482
rect 24298 67430 24310 67482
rect 24362 67430 24374 67482
rect 24426 67430 24438 67482
rect 24490 67430 34246 67482
rect 34298 67430 34310 67482
rect 34362 67430 34374 67482
rect 34426 67430 34438 67482
rect 34490 67430 44246 67482
rect 44298 67430 44310 67482
rect 44362 67430 44374 67482
rect 44426 67430 44438 67482
rect 44490 67430 54246 67482
rect 54298 67430 54310 67482
rect 54362 67430 54374 67482
rect 54426 67430 54438 67482
rect 54490 67430 64246 67482
rect 64298 67430 64310 67482
rect 64362 67430 64374 67482
rect 64426 67430 64438 67482
rect 64490 67430 68816 67482
rect 1104 67408 68816 67430
rect 16482 67368 16488 67380
rect 16443 67340 16488 67368
rect 16482 67328 16488 67340
rect 16540 67328 16546 67380
rect 934 67260 940 67312
rect 992 67300 998 67312
rect 1765 67303 1823 67309
rect 1765 67300 1777 67303
rect 992 67272 1777 67300
rect 992 67260 998 67272
rect 1765 67269 1777 67272
rect 1811 67269 1823 67303
rect 2866 67300 2872 67312
rect 2827 67272 2872 67300
rect 1765 67263 1823 67269
rect 2866 67260 2872 67272
rect 2924 67260 2930 67312
rect 8662 67300 8668 67312
rect 8623 67272 8668 67300
rect 8662 67260 8668 67272
rect 8720 67260 8726 67312
rect 10594 67300 10600 67312
rect 10555 67272 10600 67300
rect 10594 67260 10600 67272
rect 10652 67260 10658 67312
rect 18414 67300 18420 67312
rect 18375 67272 18420 67300
rect 18414 67260 18420 67272
rect 18472 67260 18478 67312
rect 24118 67260 24124 67312
rect 24176 67300 24182 67312
rect 24213 67303 24271 67309
rect 24213 67300 24225 67303
rect 24176 67272 24225 67300
rect 24176 67260 24182 67272
rect 24213 67269 24225 67272
rect 24259 67269 24271 67303
rect 26142 67300 26148 67312
rect 26103 67272 26148 67300
rect 24213 67263 24271 67269
rect 26142 67260 26148 67272
rect 26200 67260 26206 67312
rect 32030 67300 32036 67312
rect 31991 67272 32036 67300
rect 32030 67260 32036 67272
rect 32088 67260 32094 67312
rect 33962 67300 33968 67312
rect 33923 67272 33968 67300
rect 33962 67260 33968 67272
rect 34020 67260 34026 67312
rect 39758 67300 39764 67312
rect 39719 67272 39764 67300
rect 39758 67260 39764 67272
rect 39816 67260 39822 67312
rect 41690 67300 41696 67312
rect 41651 67272 41696 67300
rect 41690 67260 41696 67272
rect 41748 67260 41754 67312
rect 47578 67300 47584 67312
rect 47539 67272 47584 67300
rect 47578 67260 47584 67272
rect 47636 67260 47642 67312
rect 49510 67260 49516 67312
rect 49568 67300 49574 67312
rect 49605 67303 49663 67309
rect 49605 67300 49617 67303
rect 49568 67272 49617 67300
rect 49568 67260 49574 67272
rect 49605 67269 49617 67272
rect 49651 67269 49663 67303
rect 55306 67300 55312 67312
rect 55267 67272 55312 67300
rect 49605 67263 49663 67269
rect 55306 67260 55312 67272
rect 55364 67260 55370 67312
rect 57330 67260 57336 67312
rect 57388 67300 57394 67312
rect 57609 67303 57667 67309
rect 57609 67300 57621 67303
rect 57388 67272 57621 67300
rect 57388 67260 57394 67272
rect 57609 67269 57621 67272
rect 57655 67269 57667 67303
rect 63126 67300 63132 67312
rect 63087 67272 63132 67300
rect 57609 67263 57667 67269
rect 63126 67260 63132 67272
rect 63184 67260 63190 67312
rect 65058 67260 65064 67312
rect 65116 67300 65122 67312
rect 65613 67303 65671 67309
rect 65613 67300 65625 67303
rect 65116 67272 65625 67300
rect 65116 67260 65122 67272
rect 65613 67269 65625 67272
rect 65659 67269 65671 67303
rect 67358 67300 67364 67312
rect 67319 67272 67364 67300
rect 65613 67263 65671 67269
rect 67358 67260 67364 67272
rect 67416 67260 67422 67312
rect 4798 67124 4804 67176
rect 4856 67164 4862 67176
rect 4985 67167 5043 67173
rect 4985 67164 4997 67167
rect 4856 67136 4997 67164
rect 4856 67124 4862 67136
rect 4985 67133 4997 67136
rect 5031 67164 5043 67167
rect 5445 67167 5503 67173
rect 5445 67164 5457 67167
rect 5031 67136 5457 67164
rect 5031 67133 5043 67136
rect 4985 67127 5043 67133
rect 5445 67133 5457 67136
rect 5491 67133 5503 67167
rect 5445 67127 5503 67133
rect 12526 67124 12532 67176
rect 12584 67164 12590 67176
rect 12713 67167 12771 67173
rect 12713 67164 12725 67167
rect 12584 67136 12725 67164
rect 12584 67124 12590 67136
rect 12713 67133 12725 67136
rect 12759 67164 12771 67167
rect 13173 67167 13231 67173
rect 13173 67164 13185 67167
rect 12759 67136 13185 67164
rect 12759 67133 12771 67136
rect 12713 67127 12771 67133
rect 13173 67133 13185 67136
rect 13219 67133 13231 67167
rect 13173 67127 13231 67133
rect 20346 67124 20352 67176
rect 20404 67164 20410 67176
rect 20533 67167 20591 67173
rect 20533 67164 20545 67167
rect 20404 67136 20545 67164
rect 20404 67124 20410 67136
rect 20533 67133 20545 67136
rect 20579 67164 20591 67167
rect 20993 67167 21051 67173
rect 20993 67164 21005 67167
rect 20579 67136 21005 67164
rect 20579 67133 20591 67136
rect 20533 67127 20591 67133
rect 20993 67133 21005 67136
rect 21039 67133 21051 67167
rect 20993 67127 21051 67133
rect 24397 67167 24455 67173
rect 24397 67133 24409 67167
rect 24443 67164 24455 67167
rect 26970 67164 26976 67176
rect 24443 67136 26976 67164
rect 24443 67133 24455 67136
rect 24397 67127 24455 67133
rect 26970 67124 26976 67136
rect 27028 67124 27034 67176
rect 28074 67124 28080 67176
rect 28132 67164 28138 67176
rect 28445 67167 28503 67173
rect 28445 67164 28457 67167
rect 28132 67136 28457 67164
rect 28132 67124 28138 67136
rect 28445 67133 28457 67136
rect 28491 67164 28503 67167
rect 28905 67167 28963 67173
rect 28905 67164 28917 67167
rect 28491 67136 28917 67164
rect 28491 67133 28503 67136
rect 28445 67127 28503 67133
rect 28905 67133 28917 67136
rect 28951 67133 28963 67167
rect 28905 67127 28963 67133
rect 35894 67124 35900 67176
rect 35952 67164 35958 67176
rect 36449 67167 36507 67173
rect 36449 67164 36461 67167
rect 35952 67136 36461 67164
rect 35952 67124 35958 67136
rect 36449 67133 36461 67136
rect 36495 67164 36507 67167
rect 36909 67167 36967 67173
rect 36909 67164 36921 67167
rect 36495 67136 36921 67164
rect 36495 67133 36507 67136
rect 36449 67127 36507 67133
rect 36909 67133 36921 67136
rect 36955 67133 36967 67167
rect 36909 67127 36967 67133
rect 43714 67124 43720 67176
rect 43772 67164 43778 67176
rect 44453 67167 44511 67173
rect 44453 67164 44465 67167
rect 43772 67136 44465 67164
rect 43772 67124 43778 67136
rect 44453 67133 44465 67136
rect 44499 67164 44511 67167
rect 44913 67167 44971 67173
rect 44913 67164 44925 67167
rect 44499 67136 44925 67164
rect 44499 67133 44511 67136
rect 44453 67127 44511 67133
rect 44913 67133 44925 67136
rect 44959 67133 44971 67167
rect 44913 67127 44971 67133
rect 51442 67124 51448 67176
rect 51500 67164 51506 67176
rect 52457 67167 52515 67173
rect 52457 67164 52469 67167
rect 51500 67136 52469 67164
rect 51500 67124 51506 67136
rect 52457 67133 52469 67136
rect 52503 67164 52515 67167
rect 52917 67167 52975 67173
rect 52917 67164 52929 67167
rect 52503 67136 52929 67164
rect 52503 67133 52515 67136
rect 52457 67127 52515 67133
rect 52917 67133 52929 67136
rect 52963 67133 52975 67167
rect 59354 67164 59360 67176
rect 59315 67136 59360 67164
rect 52917 67127 52975 67133
rect 59354 67124 59360 67136
rect 59412 67164 59418 67176
rect 59909 67167 59967 67173
rect 59909 67164 59921 67167
rect 59412 67136 59921 67164
rect 59412 67124 59418 67136
rect 59909 67133 59921 67136
rect 59955 67133 59967 67167
rect 59909 67127 59967 67133
rect 64782 67124 64788 67176
rect 64840 67164 64846 67176
rect 66625 67167 66683 67173
rect 64840 67136 66576 67164
rect 64840 67124 64846 67136
rect 1949 67099 2007 67105
rect 1949 67065 1961 67099
rect 1995 67065 2007 67099
rect 1949 67059 2007 67065
rect 3053 67099 3111 67105
rect 3053 67065 3065 67099
rect 3099 67096 3111 67099
rect 3970 67096 3976 67108
rect 3099 67068 3976 67096
rect 3099 67065 3111 67068
rect 3053 67059 3111 67065
rect 1964 67028 1992 67059
rect 3970 67056 3976 67068
rect 4028 67056 4034 67108
rect 8481 67099 8539 67105
rect 8481 67065 8493 67099
rect 8527 67065 8539 67099
rect 8481 67059 8539 67065
rect 10781 67099 10839 67105
rect 10781 67065 10793 67099
rect 10827 67096 10839 67099
rect 11054 67096 11060 67108
rect 10827 67068 11060 67096
rect 10827 67065 10839 67068
rect 10781 67059 10839 67065
rect 3878 67028 3884 67040
rect 1964 67000 3884 67028
rect 3878 66988 3884 67000
rect 3936 66988 3942 67040
rect 8496 67028 8524 67059
rect 11054 67056 11060 67068
rect 11112 67056 11118 67108
rect 16574 67056 16580 67108
rect 16632 67096 16638 67108
rect 17221 67099 17279 67105
rect 17221 67096 17233 67099
rect 16632 67068 17233 67096
rect 16632 67056 16638 67068
rect 17221 67065 17233 67068
rect 17267 67065 17279 67099
rect 17221 67059 17279 67065
rect 18601 67099 18659 67105
rect 18601 67065 18613 67099
rect 18647 67096 18659 67099
rect 26329 67099 26387 67105
rect 26329 67096 26341 67099
rect 18647 67068 19104 67096
rect 18647 67065 18659 67068
rect 18601 67059 18659 67065
rect 19076 67040 19104 67068
rect 26206 67068 26341 67096
rect 9309 67031 9367 67037
rect 9309 67028 9321 67031
rect 8496 67000 9321 67028
rect 9309 66997 9321 67000
rect 9355 67028 9367 67031
rect 11698 67028 11704 67040
rect 9355 67000 11704 67028
rect 9355 66997 9367 67000
rect 9309 66991 9367 66997
rect 11698 66988 11704 67000
rect 11756 66988 11762 67040
rect 19058 66988 19064 67040
rect 19116 67028 19122 67040
rect 19153 67031 19211 67037
rect 19153 67028 19165 67031
rect 19116 67000 19165 67028
rect 19116 66988 19122 67000
rect 19153 66997 19165 67000
rect 19199 66997 19211 67031
rect 25590 67028 25596 67040
rect 25551 67000 25596 67028
rect 19153 66991 19211 66997
rect 25590 66988 25596 67000
rect 25648 67028 25654 67040
rect 26206 67028 26234 67068
rect 26329 67065 26341 67068
rect 26375 67065 26387 67099
rect 26329 67059 26387 67065
rect 32217 67099 32275 67105
rect 32217 67065 32229 67099
rect 32263 67065 32275 67099
rect 34146 67096 34152 67108
rect 34107 67068 34152 67096
rect 32217 67059 32275 67065
rect 25648 67000 26234 67028
rect 32232 67028 32260 67059
rect 34146 67056 34152 67068
rect 34204 67056 34210 67108
rect 39945 67099 40003 67105
rect 39945 67065 39957 67099
rect 39991 67065 40003 67099
rect 39945 67059 40003 67065
rect 33226 67028 33232 67040
rect 32232 67000 33232 67028
rect 25648 66988 25654 67000
rect 33226 66988 33232 67000
rect 33284 66988 33290 67040
rect 36538 66988 36544 67040
rect 36596 67028 36602 67040
rect 39209 67031 39267 67037
rect 39209 67028 39221 67031
rect 36596 67000 39221 67028
rect 36596 66988 36602 67000
rect 39209 66997 39221 67000
rect 39255 67028 39267 67031
rect 39960 67028 39988 67059
rect 41506 67056 41512 67108
rect 41564 67096 41570 67108
rect 41877 67099 41935 67105
rect 41877 67096 41889 67099
rect 41564 67068 41889 67096
rect 41564 67056 41570 67068
rect 41877 67065 41889 67068
rect 41923 67065 41935 67099
rect 47762 67096 47768 67108
rect 47723 67068 47768 67096
rect 41877 67059 41935 67065
rect 47762 67056 47768 67068
rect 47820 67056 47826 67108
rect 49789 67099 49847 67105
rect 49789 67065 49801 67099
rect 49835 67096 49847 67099
rect 55493 67099 55551 67105
rect 55493 67096 55505 67099
rect 49835 67068 50476 67096
rect 49835 67065 49847 67068
rect 49789 67059 49847 67065
rect 50448 67037 50476 67068
rect 55186 67068 55505 67096
rect 39255 67000 39988 67028
rect 50433 67031 50491 67037
rect 39255 66997 39267 67000
rect 39209 66991 39267 66997
rect 50433 66997 50445 67031
rect 50479 67028 50491 67031
rect 50798 67028 50804 67040
rect 50479 67000 50804 67028
rect 50479 66997 50491 67000
rect 50433 66991 50491 66997
rect 50798 66988 50804 67000
rect 50856 66988 50862 67040
rect 54754 67028 54760 67040
rect 54715 67000 54760 67028
rect 54754 66988 54760 67000
rect 54812 67028 54818 67040
rect 55186 67028 55214 67068
rect 55493 67065 55505 67068
rect 55539 67065 55551 67099
rect 57790 67096 57796 67108
rect 57751 67068 57796 67096
rect 55493 67059 55551 67065
rect 57790 67056 57796 67068
rect 57848 67056 57854 67108
rect 63313 67099 63371 67105
rect 63313 67065 63325 67099
rect 63359 67065 63371 67099
rect 65797 67099 65855 67105
rect 65797 67096 65809 67099
rect 63313 67059 63371 67065
rect 64846 67068 65809 67096
rect 62574 67028 62580 67040
rect 54812 67000 55214 67028
rect 62535 67000 62580 67028
rect 54812 66988 54818 67000
rect 62574 66988 62580 67000
rect 62632 67028 62638 67040
rect 63328 67028 63356 67059
rect 62632 67000 63356 67028
rect 62632 66988 62638 67000
rect 64598 66988 64604 67040
rect 64656 67028 64662 67040
rect 64693 67031 64751 67037
rect 64693 67028 64705 67031
rect 64656 67000 64705 67028
rect 64656 66988 64662 67000
rect 64693 66997 64705 67000
rect 64739 67028 64751 67031
rect 64846 67028 64874 67068
rect 65797 67065 65809 67068
rect 65843 67065 65855 67099
rect 66548 67096 66576 67136
rect 66625 67133 66637 67167
rect 66671 67164 66683 67167
rect 66990 67164 66996 67176
rect 66671 67136 66996 67164
rect 66671 67133 66683 67136
rect 66625 67127 66683 67133
rect 66990 67124 66996 67136
rect 67048 67124 67054 67176
rect 67177 67099 67235 67105
rect 67177 67096 67189 67099
rect 66548 67068 67189 67096
rect 65797 67059 65855 67065
rect 67177 67065 67189 67068
rect 67223 67096 67235 67099
rect 67913 67099 67971 67105
rect 67913 67096 67925 67099
rect 67223 67068 67925 67096
rect 67223 67065 67235 67068
rect 67177 67059 67235 67065
rect 67913 67065 67925 67068
rect 67959 67065 67971 67099
rect 67913 67059 67971 67065
rect 64739 67000 64874 67028
rect 64739 66997 64751 67000
rect 64693 66991 64751 66997
rect 1104 66938 68816 66960
rect 1104 66886 9246 66938
rect 9298 66886 9310 66938
rect 9362 66886 9374 66938
rect 9426 66886 9438 66938
rect 9490 66886 19246 66938
rect 19298 66886 19310 66938
rect 19362 66886 19374 66938
rect 19426 66886 19438 66938
rect 19490 66886 29246 66938
rect 29298 66886 29310 66938
rect 29362 66886 29374 66938
rect 29426 66886 29438 66938
rect 29490 66886 39246 66938
rect 39298 66886 39310 66938
rect 39362 66886 39374 66938
rect 39426 66886 39438 66938
rect 39490 66886 49246 66938
rect 49298 66886 49310 66938
rect 49362 66886 49374 66938
rect 49426 66886 49438 66938
rect 49490 66886 59246 66938
rect 59298 66886 59310 66938
rect 59362 66886 59374 66938
rect 59426 66886 59438 66938
rect 59490 66886 68816 66938
rect 1104 66864 68816 66886
rect 13538 66784 13544 66836
rect 13596 66824 13602 66836
rect 33781 66827 33839 66833
rect 33781 66824 33793 66827
rect 13596 66796 33793 66824
rect 13596 66784 13602 66796
rect 33781 66793 33793 66796
rect 33827 66824 33839 66827
rect 34146 66824 34152 66836
rect 33827 66796 34152 66824
rect 33827 66793 33839 66796
rect 33781 66787 33839 66793
rect 34146 66784 34152 66796
rect 34204 66784 34210 66836
rect 47762 66784 47768 66836
rect 47820 66824 47826 66836
rect 56502 66824 56508 66836
rect 47820 66796 56508 66824
rect 47820 66784 47826 66796
rect 56502 66784 56508 66796
rect 56560 66784 56566 66836
rect 66901 66827 66959 66833
rect 66901 66793 66913 66827
rect 66947 66824 66959 66827
rect 66990 66824 66996 66836
rect 66947 66796 66996 66824
rect 66947 66793 66959 66796
rect 66901 66787 66959 66793
rect 66990 66784 66996 66796
rect 67048 66784 67054 66836
rect 67542 66784 67548 66836
rect 67600 66824 67606 66836
rect 68005 66827 68063 66833
rect 68005 66824 68017 66827
rect 67600 66796 68017 66824
rect 67600 66784 67606 66796
rect 68005 66793 68017 66796
rect 68051 66793 68063 66827
rect 68005 66787 68063 66793
rect 1762 66756 1768 66768
rect 1723 66728 1768 66756
rect 1762 66716 1768 66728
rect 1820 66716 1826 66768
rect 1946 66688 1952 66700
rect 1907 66660 1952 66688
rect 1946 66648 1952 66660
rect 2004 66648 2010 66700
rect 2685 66691 2743 66697
rect 2685 66657 2697 66691
rect 2731 66688 2743 66691
rect 2774 66688 2780 66700
rect 2731 66660 2780 66688
rect 2731 66657 2743 66660
rect 2685 66651 2743 66657
rect 2774 66648 2780 66660
rect 2832 66688 2838 66700
rect 3145 66691 3203 66697
rect 3145 66688 3157 66691
rect 2832 66660 3157 66688
rect 2832 66648 2838 66660
rect 3145 66657 3157 66660
rect 3191 66657 3203 66691
rect 3145 66651 3203 66657
rect 10134 66648 10140 66700
rect 10192 66688 10198 66700
rect 57425 66691 57483 66697
rect 57425 66688 57437 66691
rect 10192 66660 57437 66688
rect 10192 66648 10198 66660
rect 57425 66657 57437 66660
rect 57471 66688 57483 66691
rect 57790 66688 57796 66700
rect 57471 66660 57796 66688
rect 57471 66657 57483 66660
rect 57425 66651 57483 66657
rect 57790 66648 57796 66660
rect 57848 66648 57854 66700
rect 66257 66691 66315 66697
rect 66257 66657 66269 66691
rect 66303 66688 66315 66691
rect 66346 66688 66352 66700
rect 66303 66660 66352 66688
rect 66303 66657 66315 66660
rect 66257 66651 66315 66657
rect 66346 66648 66352 66660
rect 66404 66688 66410 66700
rect 67913 66691 67971 66697
rect 67913 66688 67925 66691
rect 66404 66660 67925 66688
rect 66404 66648 66410 66660
rect 67913 66657 67925 66660
rect 67959 66657 67971 66691
rect 67913 66651 67971 66657
rect 3878 66580 3884 66632
rect 3936 66620 3942 66632
rect 18046 66620 18052 66632
rect 3936 66592 18052 66620
rect 3936 66580 3942 66592
rect 18046 66580 18052 66592
rect 18104 66580 18110 66632
rect 26878 66580 26884 66632
rect 26936 66620 26942 66632
rect 62574 66620 62580 66632
rect 26936 66592 62580 66620
rect 26936 66580 26942 66592
rect 62574 66580 62580 66592
rect 62632 66580 62638 66632
rect 3970 66484 3976 66496
rect 3931 66456 3976 66484
rect 3970 66444 3976 66456
rect 4028 66444 4034 66496
rect 11054 66484 11060 66496
rect 11015 66456 11060 66484
rect 11054 66444 11060 66456
rect 11112 66444 11118 66496
rect 30466 66484 30472 66496
rect 30427 66456 30472 66484
rect 30466 66444 30472 66456
rect 30524 66444 30530 66496
rect 41506 66484 41512 66496
rect 41467 66456 41512 66484
rect 41506 66444 41512 66456
rect 41564 66444 41570 66496
rect 65337 66487 65395 66493
rect 65337 66453 65349 66487
rect 65383 66484 65395 66487
rect 65702 66484 65708 66496
rect 65383 66456 65708 66484
rect 65383 66453 65395 66456
rect 65337 66447 65395 66453
rect 65702 66444 65708 66456
rect 65760 66484 65766 66496
rect 66070 66484 66076 66496
rect 65760 66456 66076 66484
rect 65760 66444 65766 66456
rect 66070 66444 66076 66456
rect 66128 66444 66134 66496
rect 1104 66394 68816 66416
rect 1104 66342 4246 66394
rect 4298 66342 4310 66394
rect 4362 66342 4374 66394
rect 4426 66342 4438 66394
rect 4490 66342 14246 66394
rect 14298 66342 14310 66394
rect 14362 66342 14374 66394
rect 14426 66342 14438 66394
rect 14490 66342 24246 66394
rect 24298 66342 24310 66394
rect 24362 66342 24374 66394
rect 24426 66342 24438 66394
rect 24490 66342 34246 66394
rect 34298 66342 34310 66394
rect 34362 66342 34374 66394
rect 34426 66342 34438 66394
rect 34490 66342 44246 66394
rect 44298 66342 44310 66394
rect 44362 66342 44374 66394
rect 44426 66342 44438 66394
rect 44490 66342 54246 66394
rect 54298 66342 54310 66394
rect 54362 66342 54374 66394
rect 54426 66342 54438 66394
rect 54490 66342 64246 66394
rect 64298 66342 64310 66394
rect 64362 66342 64374 66394
rect 64426 66342 64438 66394
rect 64490 66342 68816 66394
rect 1104 66320 68816 66342
rect 11054 66240 11060 66292
rect 11112 66280 11118 66292
rect 61470 66280 61476 66292
rect 11112 66252 61476 66280
rect 11112 66240 11118 66252
rect 61470 66240 61476 66252
rect 61528 66240 61534 66292
rect 1946 66104 1952 66156
rect 2004 66144 2010 66156
rect 2225 66147 2283 66153
rect 2225 66144 2237 66147
rect 2004 66116 2237 66144
rect 2004 66104 2010 66116
rect 2225 66113 2237 66116
rect 2271 66144 2283 66147
rect 2271 66116 16574 66144
rect 2271 66113 2283 66116
rect 2225 66107 2283 66113
rect 1581 66079 1639 66085
rect 1581 66045 1593 66079
rect 1627 66076 1639 66079
rect 4246 66076 4252 66088
rect 1627 66048 4252 66076
rect 1627 66045 1639 66048
rect 1581 66039 1639 66045
rect 4246 66036 4252 66048
rect 4304 66036 4310 66088
rect 14550 66036 14556 66088
rect 14608 66076 14614 66088
rect 14829 66079 14887 66085
rect 14829 66076 14841 66079
rect 14608 66048 14841 66076
rect 14608 66036 14614 66048
rect 14829 66045 14841 66048
rect 14875 66045 14887 66079
rect 16546 66076 16574 66116
rect 34256 66116 36492 66144
rect 30282 66076 30288 66088
rect 16546 66048 30288 66076
rect 14829 66039 14887 66045
rect 30282 66036 30288 66048
rect 30340 66036 30346 66088
rect 30190 65900 30196 65952
rect 30248 65940 30254 65952
rect 34256 65949 34284 66116
rect 36464 66088 36492 66116
rect 65518 66104 65524 66156
rect 65576 66144 65582 66156
rect 66257 66147 66315 66153
rect 66257 66144 66269 66147
rect 65576 66116 66269 66144
rect 65576 66104 65582 66116
rect 66257 66113 66269 66116
rect 66303 66113 66315 66147
rect 66257 66107 66315 66113
rect 36170 66076 36176 66088
rect 36131 66048 36176 66076
rect 36170 66036 36176 66048
rect 36228 66036 36234 66088
rect 36446 66076 36452 66088
rect 36407 66048 36452 66076
rect 36446 66036 36452 66048
rect 36504 66036 36510 66088
rect 65337 66079 65395 66085
rect 65337 66045 65349 66079
rect 65383 66076 65395 66079
rect 65794 66076 65800 66088
rect 65383 66048 65800 66076
rect 65383 66045 65395 66048
rect 65337 66039 65395 66045
rect 65794 66036 65800 66048
rect 65852 66036 65858 66088
rect 65981 66079 66039 66085
rect 65981 66045 65993 66079
rect 66027 66045 66039 66079
rect 65981 66039 66039 66045
rect 64690 66008 64696 66020
rect 64603 65980 64696 66008
rect 64690 65968 64696 65980
rect 64748 66008 64754 66020
rect 65996 66008 66024 66039
rect 66070 66036 66076 66088
rect 66128 66076 66134 66088
rect 66349 66079 66407 66085
rect 66349 66076 66361 66079
rect 66128 66048 66361 66076
rect 66128 66036 66134 66048
rect 66349 66045 66361 66048
rect 66395 66045 66407 66079
rect 68094 66076 68100 66088
rect 68055 66048 68100 66076
rect 66349 66039 66407 66045
rect 68094 66036 68100 66048
rect 68152 66036 68158 66088
rect 64748 65980 66024 66008
rect 64748 65968 64754 65980
rect 34241 65943 34299 65949
rect 34241 65940 34253 65943
rect 30248 65912 34253 65940
rect 30248 65900 30254 65912
rect 34241 65909 34253 65912
rect 34287 65909 34299 65943
rect 34882 65940 34888 65952
rect 34843 65912 34888 65940
rect 34241 65903 34299 65909
rect 34882 65900 34888 65912
rect 34940 65900 34946 65952
rect 36170 65900 36176 65952
rect 36228 65940 36234 65952
rect 36906 65940 36912 65952
rect 36228 65912 36912 65940
rect 36228 65900 36234 65912
rect 36906 65900 36912 65912
rect 36964 65900 36970 65952
rect 66714 65940 66720 65952
rect 66675 65912 66720 65940
rect 66714 65900 66720 65912
rect 66772 65900 66778 65952
rect 1104 65850 68816 65872
rect 1104 65798 9246 65850
rect 9298 65798 9310 65850
rect 9362 65798 9374 65850
rect 9426 65798 9438 65850
rect 9490 65798 19246 65850
rect 19298 65798 19310 65850
rect 19362 65798 19374 65850
rect 19426 65798 19438 65850
rect 19490 65798 29246 65850
rect 29298 65798 29310 65850
rect 29362 65798 29374 65850
rect 29426 65798 29438 65850
rect 29490 65798 39246 65850
rect 39298 65798 39310 65850
rect 39362 65798 39374 65850
rect 39426 65798 39438 65850
rect 39490 65798 49246 65850
rect 49298 65798 49310 65850
rect 49362 65798 49374 65850
rect 49426 65798 49438 65850
rect 49490 65798 59246 65850
rect 59298 65798 59310 65850
rect 59362 65798 59374 65850
rect 59426 65798 59438 65850
rect 59490 65798 68816 65850
rect 1104 65776 68816 65798
rect 16666 65696 16672 65748
rect 16724 65736 16730 65748
rect 30190 65736 30196 65748
rect 16724 65708 30196 65736
rect 16724 65696 16730 65708
rect 30190 65696 30196 65708
rect 30248 65696 30254 65748
rect 30282 65696 30288 65748
rect 30340 65736 30346 65748
rect 37918 65736 37924 65748
rect 30340 65708 37924 65736
rect 30340 65696 30346 65708
rect 37918 65696 37924 65708
rect 37976 65696 37982 65748
rect 65518 65736 65524 65748
rect 65479 65708 65524 65736
rect 65518 65696 65524 65708
rect 65576 65696 65582 65748
rect 68094 65736 68100 65748
rect 68055 65708 68100 65736
rect 68094 65696 68100 65708
rect 68152 65696 68158 65748
rect 1949 65603 2007 65609
rect 1949 65569 1961 65603
rect 1995 65600 2007 65603
rect 1995 65572 2636 65600
rect 1995 65569 2007 65572
rect 1949 65563 2007 65569
rect 1854 65396 1860 65408
rect 1815 65368 1860 65396
rect 1854 65356 1860 65368
rect 1912 65356 1918 65408
rect 2608 65405 2636 65572
rect 4614 65560 4620 65612
rect 4672 65600 4678 65612
rect 66714 65600 66720 65612
rect 4672 65572 66720 65600
rect 4672 65560 4678 65572
rect 66714 65560 66720 65572
rect 66772 65560 66778 65612
rect 4246 65492 4252 65544
rect 4304 65532 4310 65544
rect 67634 65532 67640 65544
rect 4304 65504 67640 65532
rect 4304 65492 4310 65504
rect 67634 65492 67640 65504
rect 67692 65492 67698 65544
rect 19058 65424 19064 65476
rect 19116 65464 19122 65476
rect 44637 65467 44695 65473
rect 44637 65464 44649 65467
rect 19116 65436 44649 65464
rect 19116 65424 19122 65436
rect 44637 65433 44649 65436
rect 44683 65433 44695 65467
rect 44637 65427 44695 65433
rect 2593 65399 2651 65405
rect 2593 65365 2605 65399
rect 2639 65396 2651 65399
rect 2682 65396 2688 65408
rect 2639 65368 2688 65396
rect 2639 65365 2651 65368
rect 2593 65359 2651 65365
rect 2682 65356 2688 65368
rect 2740 65356 2746 65408
rect 23014 65396 23020 65408
rect 22975 65368 23020 65396
rect 23014 65356 23020 65368
rect 23072 65356 23078 65408
rect 48685 65399 48743 65405
rect 48685 65365 48697 65399
rect 48731 65396 48743 65399
rect 56778 65396 56784 65408
rect 48731 65368 56784 65396
rect 48731 65365 48743 65368
rect 48685 65359 48743 65365
rect 56778 65356 56784 65368
rect 56836 65356 56842 65408
rect 65426 65356 65432 65408
rect 65484 65396 65490 65408
rect 66162 65396 66168 65408
rect 65484 65368 66168 65396
rect 65484 65356 65490 65368
rect 66162 65356 66168 65368
rect 66220 65396 66226 65408
rect 66809 65399 66867 65405
rect 66809 65396 66821 65399
rect 66220 65368 66821 65396
rect 66220 65356 66226 65368
rect 66809 65365 66821 65368
rect 66855 65365 66867 65399
rect 66809 65359 66867 65365
rect 1104 65306 68816 65328
rect 1104 65254 4246 65306
rect 4298 65254 4310 65306
rect 4362 65254 4374 65306
rect 4426 65254 4438 65306
rect 4490 65254 14246 65306
rect 14298 65254 14310 65306
rect 14362 65254 14374 65306
rect 14426 65254 14438 65306
rect 14490 65254 24246 65306
rect 24298 65254 24310 65306
rect 24362 65254 24374 65306
rect 24426 65254 24438 65306
rect 24490 65254 34246 65306
rect 34298 65254 34310 65306
rect 34362 65254 34374 65306
rect 34426 65254 34438 65306
rect 34490 65254 44246 65306
rect 44298 65254 44310 65306
rect 44362 65254 44374 65306
rect 44426 65254 44438 65306
rect 44490 65254 54246 65306
rect 54298 65254 54310 65306
rect 54362 65254 54374 65306
rect 54426 65254 54438 65306
rect 54490 65254 64246 65306
rect 64298 65254 64310 65306
rect 64362 65254 64374 65306
rect 64426 65254 64438 65306
rect 64490 65254 68816 65306
rect 1104 65232 68816 65254
rect 23014 65084 23020 65136
rect 23072 65124 23078 65136
rect 67174 65124 67180 65136
rect 23072 65096 67180 65124
rect 23072 65084 23078 65096
rect 67174 65084 67180 65096
rect 67232 65084 67238 65136
rect 66162 65016 66168 65068
rect 66220 65056 66226 65068
rect 66220 65028 67772 65056
rect 66220 65016 66226 65028
rect 17126 64948 17132 65000
rect 17184 64988 17190 65000
rect 17313 64991 17371 64997
rect 17313 64988 17325 64991
rect 17184 64960 17325 64988
rect 17184 64948 17190 64960
rect 17313 64957 17325 64960
rect 17359 64957 17371 64991
rect 17313 64951 17371 64957
rect 41325 64991 41383 64997
rect 41325 64957 41337 64991
rect 41371 64988 41383 64991
rect 55214 64988 55220 65000
rect 41371 64960 55220 64988
rect 41371 64957 41383 64960
rect 41325 64951 41383 64957
rect 55214 64948 55220 64960
rect 55272 64948 55278 65000
rect 66806 64948 66812 65000
rect 66864 64988 66870 65000
rect 67744 64997 67772 65028
rect 66901 64991 66959 64997
rect 66901 64988 66913 64991
rect 66864 64960 66913 64988
rect 66864 64948 66870 64960
rect 66901 64957 66913 64960
rect 66947 64988 66959 64991
rect 67505 64991 67563 64997
rect 67505 64988 67517 64991
rect 66947 64960 67517 64988
rect 66947 64957 66959 64960
rect 66901 64951 66959 64957
rect 67505 64957 67517 64960
rect 67551 64957 67563 64991
rect 67505 64951 67563 64957
rect 67729 64991 67787 64997
rect 67729 64957 67741 64991
rect 67775 64957 67787 64991
rect 67729 64951 67787 64957
rect 66254 64880 66260 64932
rect 66312 64920 66318 64932
rect 66349 64923 66407 64929
rect 66349 64920 66361 64923
rect 66312 64892 66361 64920
rect 66312 64880 66318 64892
rect 66349 64889 66361 64892
rect 66395 64920 66407 64923
rect 67361 64923 67419 64929
rect 67361 64920 67373 64923
rect 66395 64892 66668 64920
rect 66395 64889 66407 64892
rect 66349 64883 66407 64889
rect 66640 64852 66668 64892
rect 66916 64892 67373 64920
rect 66916 64852 66944 64892
rect 67361 64889 67373 64892
rect 67407 64889 67419 64923
rect 67361 64883 67419 64889
rect 67818 64880 67824 64932
rect 67876 64920 67882 64932
rect 67913 64923 67971 64929
rect 67913 64920 67925 64923
rect 67876 64892 67925 64920
rect 67876 64880 67882 64892
rect 67913 64889 67925 64892
rect 67959 64889 67971 64923
rect 67913 64883 67971 64889
rect 67634 64852 67640 64864
rect 66640 64824 66944 64852
rect 67595 64824 67640 64852
rect 67634 64812 67640 64824
rect 67692 64812 67698 64864
rect 1104 64762 68816 64784
rect 1104 64710 9246 64762
rect 9298 64710 9310 64762
rect 9362 64710 9374 64762
rect 9426 64710 9438 64762
rect 9490 64710 19246 64762
rect 19298 64710 19310 64762
rect 19362 64710 19374 64762
rect 19426 64710 19438 64762
rect 19490 64710 29246 64762
rect 29298 64710 29310 64762
rect 29362 64710 29374 64762
rect 29426 64710 29438 64762
rect 29490 64710 39246 64762
rect 39298 64710 39310 64762
rect 39362 64710 39374 64762
rect 39426 64710 39438 64762
rect 39490 64710 49246 64762
rect 49298 64710 49310 64762
rect 49362 64710 49374 64762
rect 49426 64710 49438 64762
rect 49490 64710 59246 64762
rect 59298 64710 59310 64762
rect 59362 64710 59374 64762
rect 59426 64710 59438 64762
rect 59490 64710 68816 64762
rect 1104 64688 68816 64710
rect 27522 64336 27528 64388
rect 27580 64376 27586 64388
rect 64690 64376 64696 64388
rect 27580 64348 64696 64376
rect 27580 64336 27586 64348
rect 64690 64336 64696 64348
rect 64748 64336 64754 64388
rect 2222 64308 2228 64320
rect 2183 64280 2228 64308
rect 2222 64268 2228 64280
rect 2280 64268 2286 64320
rect 6730 64268 6736 64320
rect 6788 64308 6794 64320
rect 52457 64311 52515 64317
rect 52457 64308 52469 64311
rect 6788 64280 52469 64308
rect 6788 64268 6794 64280
rect 52457 64277 52469 64280
rect 52503 64277 52515 64311
rect 52457 64271 52515 64277
rect 66162 64268 66168 64320
rect 66220 64308 66226 64320
rect 66993 64311 67051 64317
rect 66993 64308 67005 64311
rect 66220 64280 67005 64308
rect 66220 64268 66226 64280
rect 66993 64277 67005 64280
rect 67039 64308 67051 64311
rect 67634 64308 67640 64320
rect 67039 64280 67640 64308
rect 67039 64277 67051 64280
rect 66993 64271 67051 64277
rect 67634 64268 67640 64280
rect 67692 64268 67698 64320
rect 1104 64218 68816 64240
rect 1104 64166 4246 64218
rect 4298 64166 4310 64218
rect 4362 64166 4374 64218
rect 4426 64166 4438 64218
rect 4490 64166 14246 64218
rect 14298 64166 14310 64218
rect 14362 64166 14374 64218
rect 14426 64166 14438 64218
rect 14490 64166 24246 64218
rect 24298 64166 24310 64218
rect 24362 64166 24374 64218
rect 24426 64166 24438 64218
rect 24490 64166 34246 64218
rect 34298 64166 34310 64218
rect 34362 64166 34374 64218
rect 34426 64166 34438 64218
rect 34490 64166 44246 64218
rect 44298 64166 44310 64218
rect 44362 64166 44374 64218
rect 44426 64166 44438 64218
rect 44490 64166 54246 64218
rect 54298 64166 54310 64218
rect 54362 64166 54374 64218
rect 54426 64166 54438 64218
rect 54490 64166 64246 64218
rect 64298 64166 64310 64218
rect 64362 64166 64374 64218
rect 64426 64166 64438 64218
rect 64490 64166 68816 64218
rect 1104 64144 68816 64166
rect 2222 64064 2228 64116
rect 2280 64104 2286 64116
rect 38102 64104 38108 64116
rect 2280 64076 38108 64104
rect 2280 64064 2286 64076
rect 38102 64064 38108 64076
rect 38160 64064 38166 64116
rect 15381 64039 15439 64045
rect 15381 64036 15393 64039
rect 14292 64008 15393 64036
rect 14292 63977 14320 64008
rect 15381 64005 15393 64008
rect 15427 64036 15439 64039
rect 16666 64036 16672 64048
rect 15427 64008 16672 64036
rect 15427 64005 15439 64008
rect 15381 63999 15439 64005
rect 16666 63996 16672 64008
rect 16724 63996 16730 64048
rect 14277 63971 14335 63977
rect 14277 63937 14289 63971
rect 14323 63937 14335 63971
rect 68094 63968 68100 63980
rect 68055 63940 68100 63968
rect 14277 63931 14335 63937
rect 68094 63928 68100 63940
rect 68152 63928 68158 63980
rect 13998 63900 14004 63912
rect 13959 63872 14004 63900
rect 13998 63860 14004 63872
rect 14056 63900 14062 63912
rect 14737 63903 14795 63909
rect 14737 63900 14749 63903
rect 14056 63872 14749 63900
rect 14056 63860 14062 63872
rect 14737 63869 14749 63872
rect 14783 63869 14795 63903
rect 14737 63863 14795 63869
rect 67913 63835 67971 63841
rect 67913 63832 67925 63835
rect 67284 63804 67925 63832
rect 67284 63776 67312 63804
rect 67913 63801 67925 63804
rect 67959 63801 67971 63835
rect 67913 63795 67971 63801
rect 12894 63764 12900 63776
rect 12855 63736 12900 63764
rect 12894 63724 12900 63736
rect 12952 63724 12958 63776
rect 67266 63764 67272 63776
rect 67227 63736 67272 63764
rect 67266 63724 67272 63736
rect 67324 63724 67330 63776
rect 1104 63674 68816 63696
rect 1104 63622 9246 63674
rect 9298 63622 9310 63674
rect 9362 63622 9374 63674
rect 9426 63622 9438 63674
rect 9490 63622 19246 63674
rect 19298 63622 19310 63674
rect 19362 63622 19374 63674
rect 19426 63622 19438 63674
rect 19490 63622 29246 63674
rect 29298 63622 29310 63674
rect 29362 63622 29374 63674
rect 29426 63622 29438 63674
rect 29490 63622 39246 63674
rect 39298 63622 39310 63674
rect 39362 63622 39374 63674
rect 39426 63622 39438 63674
rect 39490 63622 49246 63674
rect 49298 63622 49310 63674
rect 49362 63622 49374 63674
rect 49426 63622 49438 63674
rect 49490 63622 59246 63674
rect 59298 63622 59310 63674
rect 59362 63622 59374 63674
rect 59426 63622 59438 63674
rect 59490 63622 68816 63674
rect 1104 63600 68816 63622
rect 12894 63520 12900 63572
rect 12952 63560 12958 63572
rect 27522 63560 27528 63572
rect 12952 63532 27528 63560
rect 12952 63520 12958 63532
rect 27522 63520 27528 63532
rect 27580 63520 27586 63572
rect 11333 63427 11391 63433
rect 11333 63393 11345 63427
rect 11379 63393 11391 63427
rect 11333 63387 11391 63393
rect 11977 63427 12035 63433
rect 11977 63393 11989 63427
rect 12023 63424 12035 63427
rect 12710 63424 12716 63436
rect 12023 63396 12716 63424
rect 12023 63393 12035 63396
rect 11977 63387 12035 63393
rect 11348 63356 11376 63387
rect 12710 63384 12716 63396
rect 12768 63384 12774 63436
rect 67913 63427 67971 63433
rect 67913 63424 67925 63427
rect 67284 63396 67925 63424
rect 13170 63356 13176 63368
rect 11348 63328 13176 63356
rect 13170 63316 13176 63328
rect 13228 63316 13234 63368
rect 11885 63291 11943 63297
rect 11885 63257 11897 63291
rect 11931 63288 11943 63291
rect 11931 63260 16574 63288
rect 11931 63257 11943 63260
rect 11885 63251 11943 63257
rect 12710 63220 12716 63232
rect 12671 63192 12716 63220
rect 12710 63180 12716 63192
rect 12768 63180 12774 63232
rect 13170 63220 13176 63232
rect 13131 63192 13176 63220
rect 13170 63180 13176 63192
rect 13228 63180 13234 63232
rect 16546 63220 16574 63260
rect 32398 63220 32404 63232
rect 16546 63192 32404 63220
rect 32398 63180 32404 63192
rect 32456 63180 32462 63232
rect 48869 63223 48927 63229
rect 48869 63189 48881 63223
rect 48915 63220 48927 63223
rect 50062 63220 50068 63232
rect 48915 63192 50068 63220
rect 48915 63189 48927 63192
rect 48869 63183 48927 63189
rect 50062 63180 50068 63192
rect 50120 63180 50126 63232
rect 66622 63180 66628 63232
rect 66680 63220 66686 63232
rect 67284 63229 67312 63396
rect 67913 63393 67925 63396
rect 67959 63393 67971 63427
rect 67913 63387 67971 63393
rect 68094 63288 68100 63300
rect 68055 63260 68100 63288
rect 68094 63248 68100 63260
rect 68152 63248 68158 63300
rect 67269 63223 67327 63229
rect 67269 63220 67281 63223
rect 66680 63192 67281 63220
rect 66680 63180 66686 63192
rect 67269 63189 67281 63192
rect 67315 63189 67327 63223
rect 67269 63183 67327 63189
rect 1104 63130 68816 63152
rect 1104 63078 4246 63130
rect 4298 63078 4310 63130
rect 4362 63078 4374 63130
rect 4426 63078 4438 63130
rect 4490 63078 14246 63130
rect 14298 63078 14310 63130
rect 14362 63078 14374 63130
rect 14426 63078 14438 63130
rect 14490 63078 24246 63130
rect 24298 63078 24310 63130
rect 24362 63078 24374 63130
rect 24426 63078 24438 63130
rect 24490 63078 34246 63130
rect 34298 63078 34310 63130
rect 34362 63078 34374 63130
rect 34426 63078 34438 63130
rect 34490 63078 44246 63130
rect 44298 63078 44310 63130
rect 44362 63078 44374 63130
rect 44426 63078 44438 63130
rect 44490 63078 54246 63130
rect 54298 63078 54310 63130
rect 54362 63078 54374 63130
rect 54426 63078 54438 63130
rect 54490 63078 64246 63130
rect 64298 63078 64310 63130
rect 64362 63078 64374 63130
rect 64426 63078 64438 63130
rect 64490 63078 68816 63130
rect 1104 63056 68816 63078
rect 12710 62976 12716 63028
rect 12768 63016 12774 63028
rect 19978 63016 19984 63028
rect 12768 62988 19984 63016
rect 12768 62976 12774 62988
rect 19978 62976 19984 62988
rect 20036 62976 20042 63028
rect 62758 62976 62764 63028
rect 62816 63016 62822 63028
rect 67361 63019 67419 63025
rect 67361 63016 67373 63019
rect 62816 62988 67373 63016
rect 62816 62976 62822 62988
rect 67361 62985 67373 62988
rect 67407 62985 67419 63019
rect 67361 62979 67419 62985
rect 2038 62908 2044 62960
rect 2096 62948 2102 62960
rect 7009 62951 7067 62957
rect 7009 62948 7021 62951
rect 2096 62920 7021 62948
rect 2096 62908 2102 62920
rect 7009 62917 7021 62920
rect 7055 62917 7067 62951
rect 7009 62911 7067 62917
rect 36446 62908 36452 62960
rect 36504 62948 36510 62960
rect 48958 62948 48964 62960
rect 36504 62920 48964 62948
rect 36504 62908 36510 62920
rect 48958 62908 48964 62920
rect 49016 62948 49022 62960
rect 49016 62920 49372 62948
rect 49016 62908 49022 62920
rect 3970 62840 3976 62892
rect 4028 62880 4034 62892
rect 49344 62889 49372 62920
rect 36817 62883 36875 62889
rect 36817 62880 36829 62883
rect 4028 62852 36829 62880
rect 4028 62840 4034 62852
rect 36817 62849 36829 62852
rect 36863 62849 36875 62883
rect 36817 62843 36875 62849
rect 49329 62883 49387 62889
rect 49329 62849 49341 62883
rect 49375 62849 49387 62883
rect 49329 62843 49387 62849
rect 1578 62812 1584 62824
rect 1539 62784 1584 62812
rect 1578 62772 1584 62784
rect 1636 62812 1642 62824
rect 2041 62815 2099 62821
rect 2041 62812 2053 62815
rect 1636 62784 2053 62812
rect 1636 62772 1642 62784
rect 2041 62781 2053 62784
rect 2087 62781 2099 62815
rect 9766 62812 9772 62824
rect 9727 62784 9772 62812
rect 2041 62775 2099 62781
rect 9766 62772 9772 62784
rect 9824 62772 9830 62824
rect 47397 62815 47455 62821
rect 47397 62781 47409 62815
rect 47443 62812 47455 62815
rect 49142 62812 49148 62824
rect 47443 62784 49148 62812
rect 47443 62781 47455 62784
rect 47397 62775 47455 62781
rect 49142 62772 49148 62784
rect 49200 62772 49206 62824
rect 66898 62772 66904 62824
rect 66956 62812 66962 62824
rect 67269 62815 67327 62821
rect 67269 62812 67281 62815
rect 66956 62784 67281 62812
rect 66956 62772 66962 62784
rect 67269 62781 67281 62784
rect 67315 62781 67327 62815
rect 67269 62775 67327 62781
rect 49605 62747 49663 62753
rect 49605 62713 49617 62747
rect 49651 62713 49663 62747
rect 49605 62707 49663 62713
rect 17770 62636 17776 62688
rect 17828 62676 17834 62688
rect 48777 62679 48835 62685
rect 48777 62676 48789 62679
rect 17828 62648 48789 62676
rect 17828 62636 17834 62648
rect 48777 62645 48789 62648
rect 48823 62676 48835 62679
rect 49620 62676 49648 62707
rect 50062 62704 50068 62756
rect 50120 62704 50126 62756
rect 67085 62747 67143 62753
rect 67085 62744 67097 62747
rect 66548 62716 67097 62744
rect 66548 62688 66576 62716
rect 67085 62713 67097 62716
rect 67131 62713 67143 62747
rect 67085 62707 67143 62713
rect 48823 62648 49648 62676
rect 51077 62679 51135 62685
rect 48823 62645 48835 62648
rect 48777 62639 48835 62645
rect 51077 62645 51089 62679
rect 51123 62676 51135 62679
rect 51442 62676 51448 62688
rect 51123 62648 51448 62676
rect 51123 62645 51135 62648
rect 51077 62639 51135 62645
rect 51442 62636 51448 62648
rect 51500 62636 51506 62688
rect 66530 62676 66536 62688
rect 66491 62648 66536 62676
rect 66530 62636 66536 62648
rect 66588 62636 66594 62688
rect 1104 62586 68816 62608
rect 1104 62534 9246 62586
rect 9298 62534 9310 62586
rect 9362 62534 9374 62586
rect 9426 62534 9438 62586
rect 9490 62534 19246 62586
rect 19298 62534 19310 62586
rect 19362 62534 19374 62586
rect 19426 62534 19438 62586
rect 19490 62534 29246 62586
rect 29298 62534 29310 62586
rect 29362 62534 29374 62586
rect 29426 62534 29438 62586
rect 29490 62534 39246 62586
rect 39298 62534 39310 62586
rect 39362 62534 39374 62586
rect 39426 62534 39438 62586
rect 39490 62534 49246 62586
rect 49298 62534 49310 62586
rect 49362 62534 49374 62586
rect 49426 62534 49438 62586
rect 49490 62534 59246 62586
rect 59298 62534 59310 62586
rect 59362 62534 59374 62586
rect 59426 62534 59438 62586
rect 59490 62534 68816 62586
rect 1104 62512 68816 62534
rect 9766 62432 9772 62484
rect 9824 62472 9830 62484
rect 64690 62472 64696 62484
rect 9824 62444 64696 62472
rect 9824 62432 9830 62444
rect 64690 62432 64696 62444
rect 64748 62432 64754 62484
rect 65058 62432 65064 62484
rect 65116 62472 65122 62484
rect 66898 62472 66904 62484
rect 65116 62444 66904 62472
rect 65116 62432 65122 62444
rect 66898 62432 66904 62444
rect 66956 62432 66962 62484
rect 48958 62404 48964 62416
rect 48919 62376 48964 62404
rect 48958 62364 48964 62376
rect 49016 62364 49022 62416
rect 49602 62364 49608 62416
rect 49660 62404 49666 62416
rect 66530 62404 66536 62416
rect 49660 62376 66536 62404
rect 49660 62364 49666 62376
rect 66530 62364 66536 62376
rect 66588 62364 66594 62416
rect 20257 62339 20315 62345
rect 20257 62305 20269 62339
rect 20303 62305 20315 62339
rect 20257 62299 20315 62305
rect 20349 62339 20407 62345
rect 20349 62305 20361 62339
rect 20395 62336 20407 62339
rect 20395 62308 25176 62336
rect 20395 62305 20407 62308
rect 20349 62299 20407 62305
rect 20272 62268 20300 62299
rect 20993 62271 21051 62277
rect 20993 62268 21005 62271
rect 20272 62240 21005 62268
rect 20993 62237 21005 62240
rect 21039 62268 21051 62271
rect 25148 62268 25176 62308
rect 32490 62268 32496 62280
rect 21039 62240 22232 62268
rect 25148 62240 32496 62268
rect 21039 62237 21051 62240
rect 20993 62231 21051 62237
rect 13541 62203 13599 62209
rect 13541 62169 13553 62203
rect 13587 62200 13599 62203
rect 22204 62200 22232 62240
rect 32490 62228 32496 62240
rect 32548 62228 32554 62280
rect 33134 62200 33140 62212
rect 13587 62172 21128 62200
rect 22204 62172 33140 62200
rect 13587 62169 13599 62172
rect 13541 62163 13599 62169
rect 21100 62132 21128 62172
rect 33134 62160 33140 62172
rect 33192 62160 33198 62212
rect 55030 62132 55036 62144
rect 21100 62104 55036 62132
rect 55030 62092 55036 62104
rect 55088 62092 55094 62144
rect 1104 62042 68816 62064
rect 1104 61990 4246 62042
rect 4298 61990 4310 62042
rect 4362 61990 4374 62042
rect 4426 61990 4438 62042
rect 4490 61990 14246 62042
rect 14298 61990 14310 62042
rect 14362 61990 14374 62042
rect 14426 61990 14438 62042
rect 14490 61990 24246 62042
rect 24298 61990 24310 62042
rect 24362 61990 24374 62042
rect 24426 61990 24438 62042
rect 24490 61990 34246 62042
rect 34298 61990 34310 62042
rect 34362 61990 34374 62042
rect 34426 61990 34438 62042
rect 34490 61990 44246 62042
rect 44298 61990 44310 62042
rect 44362 61990 44374 62042
rect 44426 61990 44438 62042
rect 44490 61990 54246 62042
rect 54298 61990 54310 62042
rect 54362 61990 54374 62042
rect 54426 61990 54438 62042
rect 54490 61990 64246 62042
rect 64298 61990 64310 62042
rect 64362 61990 64374 62042
rect 64426 61990 64438 62042
rect 64490 61990 68816 62042
rect 1104 61968 68816 61990
rect 36909 61863 36967 61869
rect 36909 61829 36921 61863
rect 36955 61860 36967 61863
rect 67266 61860 67272 61872
rect 36955 61832 67272 61860
rect 36955 61829 36967 61832
rect 36909 61823 36967 61829
rect 67266 61820 67272 61832
rect 67324 61820 67330 61872
rect 17497 61727 17555 61733
rect 17497 61693 17509 61727
rect 17543 61724 17555 61727
rect 67266 61724 67272 61736
rect 17543 61696 26234 61724
rect 17543 61693 17555 61696
rect 17497 61687 17555 61693
rect 1949 61659 2007 61665
rect 1949 61625 1961 61659
rect 1995 61656 2007 61659
rect 26206 61656 26234 61696
rect 45526 61696 67272 61724
rect 45526 61656 45554 61696
rect 67266 61684 67272 61696
rect 67324 61684 67330 61736
rect 1995 61628 2360 61656
rect 26206 61628 45554 61656
rect 1995 61625 2007 61628
rect 1949 61619 2007 61625
rect 2332 61600 2360 61628
rect 1854 61588 1860 61600
rect 1815 61560 1860 61588
rect 1854 61548 1860 61560
rect 1912 61548 1918 61600
rect 2314 61548 2320 61600
rect 2372 61588 2378 61600
rect 2501 61591 2559 61597
rect 2501 61588 2513 61591
rect 2372 61560 2513 61588
rect 2372 61548 2378 61560
rect 2501 61557 2513 61560
rect 2547 61557 2559 61591
rect 2501 61551 2559 61557
rect 1104 61498 68816 61520
rect 1104 61446 9246 61498
rect 9298 61446 9310 61498
rect 9362 61446 9374 61498
rect 9426 61446 9438 61498
rect 9490 61446 19246 61498
rect 19298 61446 19310 61498
rect 19362 61446 19374 61498
rect 19426 61446 19438 61498
rect 19490 61446 29246 61498
rect 29298 61446 29310 61498
rect 29362 61446 29374 61498
rect 29426 61446 29438 61498
rect 29490 61446 39246 61498
rect 39298 61446 39310 61498
rect 39362 61446 39374 61498
rect 39426 61446 39438 61498
rect 39490 61446 49246 61498
rect 49298 61446 49310 61498
rect 49362 61446 49374 61498
rect 49426 61446 49438 61498
rect 49490 61446 59246 61498
rect 59298 61446 59310 61498
rect 59362 61446 59374 61498
rect 59426 61446 59438 61498
rect 59490 61446 68816 61498
rect 1104 61424 68816 61446
rect 67453 61251 67511 61257
rect 67453 61217 67465 61251
rect 67499 61248 67511 61251
rect 68094 61248 68100 61260
rect 67499 61220 68100 61248
rect 67499 61217 67511 61220
rect 67453 61211 67511 61217
rect 68094 61208 68100 61220
rect 68152 61208 68158 61260
rect 1104 60954 68816 60976
rect 1104 60902 4246 60954
rect 4298 60902 4310 60954
rect 4362 60902 4374 60954
rect 4426 60902 4438 60954
rect 4490 60902 14246 60954
rect 14298 60902 14310 60954
rect 14362 60902 14374 60954
rect 14426 60902 14438 60954
rect 14490 60902 24246 60954
rect 24298 60902 24310 60954
rect 24362 60902 24374 60954
rect 24426 60902 24438 60954
rect 24490 60902 34246 60954
rect 34298 60902 34310 60954
rect 34362 60902 34374 60954
rect 34426 60902 34438 60954
rect 34490 60902 44246 60954
rect 44298 60902 44310 60954
rect 44362 60902 44374 60954
rect 44426 60902 44438 60954
rect 44490 60902 54246 60954
rect 54298 60902 54310 60954
rect 54362 60902 54374 60954
rect 54426 60902 54438 60954
rect 54490 60902 64246 60954
rect 64298 60902 64310 60954
rect 64362 60902 64374 60954
rect 64426 60902 64438 60954
rect 64490 60902 68816 60954
rect 1104 60880 68816 60902
rect 51442 60704 51448 60716
rect 51403 60676 51448 60704
rect 51442 60664 51448 60676
rect 51500 60664 51506 60716
rect 1104 60410 68816 60432
rect 1104 60358 9246 60410
rect 9298 60358 9310 60410
rect 9362 60358 9374 60410
rect 9426 60358 9438 60410
rect 9490 60358 19246 60410
rect 19298 60358 19310 60410
rect 19362 60358 19374 60410
rect 19426 60358 19438 60410
rect 19490 60358 29246 60410
rect 29298 60358 29310 60410
rect 29362 60358 29374 60410
rect 29426 60358 29438 60410
rect 29490 60358 39246 60410
rect 39298 60358 39310 60410
rect 39362 60358 39374 60410
rect 39426 60358 39438 60410
rect 39490 60358 49246 60410
rect 49298 60358 49310 60410
rect 49362 60358 49374 60410
rect 49426 60358 49438 60410
rect 49490 60358 59246 60410
rect 59298 60358 59310 60410
rect 59362 60358 59374 60410
rect 59426 60358 59438 60410
rect 59490 60358 68816 60410
rect 1104 60336 68816 60358
rect 51442 60188 51448 60240
rect 51500 60228 51506 60240
rect 51500 60200 52684 60228
rect 51500 60188 51506 60200
rect 1762 60160 1768 60172
rect 1723 60132 1768 60160
rect 1762 60120 1768 60132
rect 1820 60120 1826 60172
rect 1854 60120 1860 60172
rect 1912 60160 1918 60172
rect 1949 60163 2007 60169
rect 1949 60160 1961 60163
rect 1912 60132 1961 60160
rect 1912 60120 1918 60132
rect 1949 60129 1961 60132
rect 1995 60160 2007 60163
rect 2501 60163 2559 60169
rect 2501 60160 2513 60163
rect 1995 60132 2513 60160
rect 1995 60129 2007 60132
rect 1949 60123 2007 60129
rect 2501 60129 2513 60132
rect 2547 60129 2559 60163
rect 2501 60123 2559 60129
rect 50982 60120 50988 60172
rect 51040 60160 51046 60172
rect 52221 60163 52279 60169
rect 52221 60160 52233 60163
rect 51040 60132 52233 60160
rect 51040 60120 51046 60132
rect 52221 60129 52233 60132
rect 52267 60129 52279 60163
rect 52362 60160 52368 60172
rect 52323 60132 52368 60160
rect 52221 60123 52279 60129
rect 52362 60120 52368 60132
rect 52420 60120 52426 60172
rect 52656 60169 52684 60200
rect 52457 60163 52515 60169
rect 52457 60129 52469 60163
rect 52503 60129 52515 60163
rect 52457 60123 52515 60129
rect 52641 60163 52699 60169
rect 52641 60129 52653 60163
rect 52687 60160 52699 60163
rect 52687 60132 55214 60160
rect 52687 60129 52699 60132
rect 52641 60123 52699 60129
rect 2130 60052 2136 60104
rect 2188 60092 2194 60104
rect 15657 60095 15715 60101
rect 15657 60092 15669 60095
rect 2188 60064 15669 60092
rect 2188 60052 2194 60064
rect 15657 60061 15669 60064
rect 15703 60061 15715 60095
rect 15657 60055 15715 60061
rect 44082 60052 44088 60104
rect 44140 60092 44146 60104
rect 49602 60092 49608 60104
rect 44140 60064 49608 60092
rect 44140 60052 44146 60064
rect 49602 60052 49608 60064
rect 49660 60052 49666 60104
rect 51626 60052 51632 60104
rect 51684 60092 51690 60104
rect 52472 60092 52500 60123
rect 51684 60064 52500 60092
rect 55186 60092 55214 60132
rect 56502 60120 56508 60172
rect 56560 60160 56566 60172
rect 57149 60163 57207 60169
rect 57149 60160 57161 60163
rect 56560 60132 57161 60160
rect 56560 60120 56566 60132
rect 57149 60129 57161 60132
rect 57195 60129 57207 60163
rect 57149 60123 57207 60129
rect 58618 60092 58624 60104
rect 55186 60064 58624 60092
rect 51684 60052 51690 60064
rect 58618 60052 58624 60064
rect 58676 60052 58682 60104
rect 30282 59984 30288 60036
rect 30340 60024 30346 60036
rect 66806 60024 66812 60036
rect 30340 59996 66812 60024
rect 30340 59984 30346 59996
rect 66806 59984 66812 59996
rect 66864 59984 66870 60036
rect 2590 59916 2596 59968
rect 2648 59956 2654 59968
rect 44361 59959 44419 59965
rect 44361 59956 44373 59959
rect 2648 59928 44373 59956
rect 2648 59916 2654 59928
rect 44361 59925 44373 59928
rect 44407 59925 44419 59959
rect 47394 59956 47400 59968
rect 47355 59928 47400 59956
rect 44361 59919 44419 59925
rect 47394 59916 47400 59928
rect 47452 59916 47458 59968
rect 50430 59916 50436 59968
rect 50488 59956 50494 59968
rect 50982 59956 50988 59968
rect 50488 59928 50988 59956
rect 50488 59916 50494 59928
rect 50982 59916 50988 59928
rect 51040 59956 51046 59968
rect 51445 59959 51503 59965
rect 51445 59956 51457 59959
rect 51040 59928 51457 59956
rect 51040 59916 51046 59928
rect 51445 59925 51457 59928
rect 51491 59925 51503 59959
rect 52086 59956 52092 59968
rect 52047 59928 52092 59956
rect 51445 59919 51503 59925
rect 52086 59916 52092 59928
rect 52144 59916 52150 59968
rect 53190 59956 53196 59968
rect 53151 59928 53196 59956
rect 53190 59916 53196 59928
rect 53248 59916 53254 59968
rect 1104 59866 68816 59888
rect 1104 59814 4246 59866
rect 4298 59814 4310 59866
rect 4362 59814 4374 59866
rect 4426 59814 4438 59866
rect 4490 59814 14246 59866
rect 14298 59814 14310 59866
rect 14362 59814 14374 59866
rect 14426 59814 14438 59866
rect 14490 59814 24246 59866
rect 24298 59814 24310 59866
rect 24362 59814 24374 59866
rect 24426 59814 24438 59866
rect 24490 59814 34246 59866
rect 34298 59814 34310 59866
rect 34362 59814 34374 59866
rect 34426 59814 34438 59866
rect 34490 59814 44246 59866
rect 44298 59814 44310 59866
rect 44362 59814 44374 59866
rect 44426 59814 44438 59866
rect 44490 59814 54246 59866
rect 54298 59814 54310 59866
rect 54362 59814 54374 59866
rect 54426 59814 54438 59866
rect 54490 59814 64246 59866
rect 64298 59814 64310 59866
rect 64362 59814 64374 59866
rect 64426 59814 64438 59866
rect 64490 59814 68816 59866
rect 1104 59792 68816 59814
rect 14826 59576 14832 59628
rect 14884 59616 14890 59628
rect 66254 59616 66260 59628
rect 14884 59588 66260 59616
rect 14884 59576 14890 59588
rect 66254 59576 66260 59588
rect 66312 59576 66318 59628
rect 16117 59551 16175 59557
rect 16117 59517 16129 59551
rect 16163 59548 16175 59551
rect 16393 59551 16451 59557
rect 16163 59520 16344 59548
rect 16163 59517 16175 59520
rect 16117 59511 16175 59517
rect 16316 59480 16344 59520
rect 16393 59517 16405 59551
rect 16439 59548 16451 59551
rect 16666 59548 16672 59560
rect 16439 59520 16672 59548
rect 16439 59517 16451 59520
rect 16393 59511 16451 59517
rect 16666 59508 16672 59520
rect 16724 59548 16730 59560
rect 17218 59548 17224 59560
rect 16724 59520 17224 59548
rect 16724 59508 16730 59520
rect 17218 59508 17224 59520
rect 17276 59508 17282 59560
rect 66714 59508 66720 59560
rect 66772 59548 66778 59560
rect 67085 59551 67143 59557
rect 67085 59548 67097 59551
rect 66772 59520 67097 59548
rect 66772 59508 66778 59520
rect 67085 59517 67097 59520
rect 67131 59517 67143 59551
rect 67085 59511 67143 59517
rect 17037 59483 17095 59489
rect 17037 59480 17049 59483
rect 16316 59452 17049 59480
rect 17037 59449 17049 59452
rect 17083 59480 17095 59483
rect 33502 59480 33508 59492
rect 17083 59452 33508 59480
rect 17083 59449 17095 59452
rect 17037 59443 17095 59449
rect 33502 59440 33508 59452
rect 33560 59440 33566 59492
rect 14826 59412 14832 59424
rect 14787 59384 14832 59412
rect 14826 59372 14832 59384
rect 14884 59372 14890 59424
rect 17218 59372 17224 59424
rect 17276 59412 17282 59424
rect 17497 59415 17555 59421
rect 17497 59412 17509 59415
rect 17276 59384 17509 59412
rect 17276 59372 17282 59384
rect 17497 59381 17509 59384
rect 17543 59381 17555 59415
rect 51626 59412 51632 59424
rect 51587 59384 51632 59412
rect 17497 59375 17555 59381
rect 51626 59372 51632 59384
rect 51684 59372 51690 59424
rect 52362 59372 52368 59424
rect 52420 59412 52426 59424
rect 52825 59415 52883 59421
rect 52825 59412 52837 59415
rect 52420 59384 52837 59412
rect 52420 59372 52426 59384
rect 52825 59381 52837 59384
rect 52871 59412 52883 59415
rect 58710 59412 58716 59424
rect 52871 59384 58716 59412
rect 52871 59381 52883 59384
rect 52825 59375 52883 59381
rect 58710 59372 58716 59384
rect 58768 59372 58774 59424
rect 1104 59322 68816 59344
rect 1104 59270 9246 59322
rect 9298 59270 9310 59322
rect 9362 59270 9374 59322
rect 9426 59270 9438 59322
rect 9490 59270 19246 59322
rect 19298 59270 19310 59322
rect 19362 59270 19374 59322
rect 19426 59270 19438 59322
rect 19490 59270 29246 59322
rect 29298 59270 29310 59322
rect 29362 59270 29374 59322
rect 29426 59270 29438 59322
rect 29490 59270 39246 59322
rect 39298 59270 39310 59322
rect 39362 59270 39374 59322
rect 39426 59270 39438 59322
rect 39490 59270 49246 59322
rect 49298 59270 49310 59322
rect 49362 59270 49374 59322
rect 49426 59270 49438 59322
rect 49490 59270 59246 59322
rect 59298 59270 59310 59322
rect 59362 59270 59374 59322
rect 59426 59270 59438 59322
rect 59490 59270 68816 59322
rect 1104 59248 68816 59270
rect 10505 59007 10563 59013
rect 10505 58973 10517 59007
rect 10551 59004 10563 59007
rect 66622 59004 66628 59016
rect 10551 58976 66628 59004
rect 10551 58973 10563 58976
rect 10505 58967 10563 58973
rect 66622 58964 66628 58976
rect 66680 58964 66686 59016
rect 33134 58896 33140 58948
rect 33192 58936 33198 58948
rect 33410 58936 33416 58948
rect 33192 58908 33416 58936
rect 33192 58896 33198 58908
rect 33410 58896 33416 58908
rect 33468 58936 33474 58948
rect 43257 58939 43315 58945
rect 43257 58936 43269 58939
rect 33468 58908 43269 58936
rect 33468 58896 33474 58908
rect 43257 58905 43269 58908
rect 43303 58936 43315 58939
rect 43990 58936 43996 58948
rect 43303 58908 43996 58936
rect 43303 58905 43315 58908
rect 43257 58899 43315 58905
rect 43990 58896 43996 58908
rect 44048 58896 44054 58948
rect 13446 58868 13452 58880
rect 13407 58840 13452 58868
rect 13446 58828 13452 58840
rect 13504 58828 13510 58880
rect 64138 58828 64144 58880
rect 64196 58868 64202 58880
rect 64325 58871 64383 58877
rect 64325 58868 64337 58871
rect 64196 58840 64337 58868
rect 64196 58828 64202 58840
rect 64325 58837 64337 58840
rect 64371 58837 64383 58871
rect 64325 58831 64383 58837
rect 1104 58778 68816 58800
rect 1104 58726 4246 58778
rect 4298 58726 4310 58778
rect 4362 58726 4374 58778
rect 4426 58726 4438 58778
rect 4490 58726 14246 58778
rect 14298 58726 14310 58778
rect 14362 58726 14374 58778
rect 14426 58726 14438 58778
rect 14490 58726 24246 58778
rect 24298 58726 24310 58778
rect 24362 58726 24374 58778
rect 24426 58726 24438 58778
rect 24490 58726 34246 58778
rect 34298 58726 34310 58778
rect 34362 58726 34374 58778
rect 34426 58726 34438 58778
rect 34490 58726 44246 58778
rect 44298 58726 44310 58778
rect 44362 58726 44374 58778
rect 44426 58726 44438 58778
rect 44490 58726 54246 58778
rect 54298 58726 54310 58778
rect 54362 58726 54374 58778
rect 54426 58726 54438 58778
rect 54490 58726 64246 58778
rect 64298 58726 64310 58778
rect 64362 58726 64374 58778
rect 64426 58726 64438 58778
rect 64490 58726 68816 58778
rect 1104 58704 68816 58726
rect 8202 58624 8208 58676
rect 8260 58664 8266 58676
rect 29086 58664 29092 58676
rect 8260 58636 29092 58664
rect 8260 58624 8266 58636
rect 29086 58624 29092 58636
rect 29144 58664 29150 58676
rect 30282 58664 30288 58676
rect 29144 58636 30288 58664
rect 29144 58624 29150 58636
rect 30282 58624 30288 58636
rect 30340 58624 30346 58676
rect 42518 58624 42524 58676
rect 42576 58664 42582 58676
rect 42576 58636 44312 58664
rect 42576 58624 42582 58636
rect 3878 58556 3884 58608
rect 3936 58596 3942 58608
rect 44174 58596 44180 58608
rect 3936 58568 44180 58596
rect 3936 58556 3942 58568
rect 44174 58556 44180 58568
rect 44232 58556 44238 58608
rect 2682 58488 2688 58540
rect 2740 58528 2746 58540
rect 23201 58531 23259 58537
rect 23201 58528 23213 58531
rect 2740 58500 23213 58528
rect 2740 58488 2746 58500
rect 23201 58497 23213 58500
rect 23247 58497 23259 58531
rect 43990 58528 43996 58540
rect 43951 58500 43996 58528
rect 23201 58491 23259 58497
rect 43990 58488 43996 58500
rect 44048 58488 44054 58540
rect 44082 58488 44088 58540
rect 44140 58528 44146 58540
rect 44284 58537 44312 58636
rect 44450 58556 44456 58608
rect 44508 58596 44514 58608
rect 48777 58599 48835 58605
rect 48777 58596 48789 58599
rect 44508 58568 48789 58596
rect 44508 58556 44514 58568
rect 48777 58565 48789 58568
rect 48823 58565 48835 58599
rect 68094 58596 68100 58608
rect 68055 58568 68100 58596
rect 48777 58559 48835 58565
rect 68094 58556 68100 58568
rect 68152 58556 68158 58608
rect 44269 58531 44327 58537
rect 44140 58500 44185 58528
rect 44140 58488 44146 58500
rect 44269 58497 44281 58531
rect 44315 58497 44327 58531
rect 44269 58491 44327 58497
rect 22741 58463 22799 58469
rect 22741 58429 22753 58463
rect 22787 58429 22799 58463
rect 27982 58460 27988 58472
rect 27943 58432 27988 58460
rect 22741 58423 22799 58429
rect 22756 58392 22784 58423
rect 27982 58420 27988 58432
rect 28040 58420 28046 58472
rect 34514 58460 34520 58472
rect 34475 58432 34520 58460
rect 34514 58420 34520 58432
rect 34572 58420 34578 58472
rect 43254 58420 43260 58472
rect 43312 58460 43318 58472
rect 44177 58463 44235 58469
rect 44177 58460 44189 58463
rect 43312 58432 44189 58460
rect 43312 58420 43318 58432
rect 44177 58429 44189 58432
rect 44223 58429 44235 58463
rect 44177 58423 44235 58429
rect 67358 58392 67364 58404
rect 22756 58364 67364 58392
rect 67358 58352 67364 58364
rect 67416 58352 67422 58404
rect 67913 58395 67971 58401
rect 67913 58361 67925 58395
rect 67959 58361 67971 58395
rect 67913 58355 67971 58361
rect 42518 58324 42524 58336
rect 42479 58296 42524 58324
rect 42518 58284 42524 58296
rect 42576 58284 42582 58336
rect 43254 58324 43260 58336
rect 43215 58296 43260 58324
rect 43254 58284 43260 58296
rect 43312 58284 43318 58336
rect 43806 58324 43812 58336
rect 43767 58296 43812 58324
rect 43806 58284 43812 58296
rect 43864 58284 43870 58336
rect 66990 58284 66996 58336
rect 67048 58324 67054 58336
rect 67269 58327 67327 58333
rect 67269 58324 67281 58327
rect 67048 58296 67281 58324
rect 67048 58284 67054 58296
rect 67269 58293 67281 58296
rect 67315 58324 67327 58327
rect 67928 58324 67956 58355
rect 67315 58296 67956 58324
rect 67315 58293 67327 58296
rect 67269 58287 67327 58293
rect 1104 58234 68816 58256
rect 1104 58182 9246 58234
rect 9298 58182 9310 58234
rect 9362 58182 9374 58234
rect 9426 58182 9438 58234
rect 9490 58182 19246 58234
rect 19298 58182 19310 58234
rect 19362 58182 19374 58234
rect 19426 58182 19438 58234
rect 19490 58182 29246 58234
rect 29298 58182 29310 58234
rect 29362 58182 29374 58234
rect 29426 58182 29438 58234
rect 29490 58182 39246 58234
rect 39298 58182 39310 58234
rect 39362 58182 39374 58234
rect 39426 58182 39438 58234
rect 39490 58182 49246 58234
rect 49298 58182 49310 58234
rect 49362 58182 49374 58234
rect 49426 58182 49438 58234
rect 49490 58182 59246 58234
rect 59298 58182 59310 58234
rect 59362 58182 59374 58234
rect 59426 58182 59438 58234
rect 59490 58182 68816 58234
rect 1104 58160 68816 58182
rect 6825 58123 6883 58129
rect 6825 58089 6837 58123
rect 6871 58120 6883 58123
rect 6914 58120 6920 58132
rect 6871 58092 6920 58120
rect 6871 58089 6883 58092
rect 6825 58083 6883 58089
rect 6914 58080 6920 58092
rect 6972 58120 6978 58132
rect 8202 58120 8208 58132
rect 6972 58092 8208 58120
rect 6972 58080 6978 58092
rect 8202 58080 8208 58092
rect 8260 58080 8266 58132
rect 34514 58080 34520 58132
rect 34572 58120 34578 58132
rect 46842 58120 46848 58132
rect 34572 58092 46848 58120
rect 34572 58080 34578 58092
rect 46842 58080 46848 58092
rect 46900 58080 46906 58132
rect 5997 58055 6055 58061
rect 5997 58021 6009 58055
rect 6043 58052 6055 58055
rect 65518 58052 65524 58064
rect 6043 58024 7512 58052
rect 65479 58024 65524 58052
rect 6043 58021 6055 58024
rect 5997 58015 6055 58021
rect 4706 57944 4712 57996
rect 4764 57984 4770 57996
rect 5629 57987 5687 57993
rect 5629 57984 5641 57987
rect 4764 57956 5641 57984
rect 4764 57944 4770 57956
rect 5629 57953 5641 57956
rect 5675 57953 5687 57987
rect 5629 57947 5687 57953
rect 6089 57987 6147 57993
rect 6089 57953 6101 57987
rect 6135 57984 6147 57987
rect 6914 57984 6920 57996
rect 6135 57956 6920 57984
rect 6135 57953 6147 57956
rect 6089 57947 6147 57953
rect 6914 57944 6920 57956
rect 6972 57944 6978 57996
rect 6362 57916 6368 57928
rect 6323 57888 6368 57916
rect 6362 57876 6368 57888
rect 6420 57876 6426 57928
rect 7484 57925 7512 58024
rect 65518 58012 65524 58024
rect 65576 58012 65582 58064
rect 27982 57944 27988 57996
rect 28040 57984 28046 57996
rect 48866 57984 48872 57996
rect 28040 57956 48872 57984
rect 28040 57944 28046 57956
rect 48866 57944 48872 57956
rect 48924 57944 48930 57996
rect 65058 57984 65064 57996
rect 65019 57956 65064 57984
rect 65058 57944 65064 57956
rect 65116 57944 65122 57996
rect 7469 57919 7527 57925
rect 7469 57885 7481 57919
rect 7515 57916 7527 57919
rect 50246 57916 50252 57928
rect 7515 57888 50252 57916
rect 7515 57885 7527 57888
rect 7469 57879 7527 57885
rect 50246 57876 50252 57888
rect 50304 57876 50310 57928
rect 5445 57851 5503 57857
rect 5445 57817 5457 57851
rect 5491 57848 5503 57851
rect 5491 57820 16574 57848
rect 5491 57817 5503 57820
rect 5445 57811 5503 57817
rect 4706 57780 4712 57792
rect 4667 57752 4712 57780
rect 4706 57740 4712 57752
rect 4764 57740 4770 57792
rect 8202 57780 8208 57792
rect 8163 57752 8208 57780
rect 8202 57740 8208 57752
rect 8260 57740 8266 57792
rect 16546 57780 16574 57820
rect 26970 57808 26976 57860
rect 27028 57848 27034 57860
rect 28077 57851 28135 57857
rect 28077 57848 28089 57851
rect 27028 57820 28089 57848
rect 27028 57808 27034 57820
rect 28077 57817 28089 57820
rect 28123 57817 28135 57851
rect 28077 57811 28135 57817
rect 27798 57780 27804 57792
rect 16546 57752 27804 57780
rect 27798 57740 27804 57752
rect 27856 57740 27862 57792
rect 36170 57780 36176 57792
rect 36131 57752 36176 57780
rect 36170 57740 36176 57752
rect 36228 57740 36234 57792
rect 43438 57780 43444 57792
rect 43399 57752 43444 57780
rect 43438 57740 43444 57752
rect 43496 57780 43502 57792
rect 44082 57780 44088 57792
rect 43496 57752 44088 57780
rect 43496 57740 43502 57752
rect 44082 57740 44088 57752
rect 44140 57740 44146 57792
rect 45278 57780 45284 57792
rect 45239 57752 45284 57780
rect 45278 57740 45284 57752
rect 45336 57740 45342 57792
rect 55122 57780 55128 57792
rect 55083 57752 55128 57780
rect 55122 57740 55128 57752
rect 55180 57740 55186 57792
rect 58618 57740 58624 57792
rect 58676 57780 58682 57792
rect 64417 57783 64475 57789
rect 64417 57780 64429 57783
rect 58676 57752 64429 57780
rect 58676 57740 58682 57752
rect 64417 57749 64429 57752
rect 64463 57780 64475 57783
rect 65058 57780 65064 57792
rect 64463 57752 65064 57780
rect 64463 57749 64475 57752
rect 64417 57743 64475 57749
rect 65058 57740 65064 57752
rect 65116 57740 65122 57792
rect 1104 57690 68816 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 14246 57690
rect 14298 57638 14310 57690
rect 14362 57638 14374 57690
rect 14426 57638 14438 57690
rect 14490 57638 24246 57690
rect 24298 57638 24310 57690
rect 24362 57638 24374 57690
rect 24426 57638 24438 57690
rect 24490 57638 34246 57690
rect 34298 57638 34310 57690
rect 34362 57638 34374 57690
rect 34426 57638 34438 57690
rect 34490 57638 44246 57690
rect 44298 57638 44310 57690
rect 44362 57638 44374 57690
rect 44426 57638 44438 57690
rect 44490 57638 54246 57690
rect 54298 57638 54310 57690
rect 54362 57638 54374 57690
rect 54426 57638 54438 57690
rect 54490 57638 64246 57690
rect 64298 57638 64310 57690
rect 64362 57638 64374 57690
rect 64426 57638 64438 57690
rect 64490 57638 68816 57690
rect 1104 57616 68816 57638
rect 8202 57536 8208 57588
rect 8260 57576 8266 57588
rect 44910 57576 44916 57588
rect 8260 57548 44916 57576
rect 8260 57536 8266 57548
rect 44910 57536 44916 57548
rect 44968 57536 44974 57588
rect 45278 57536 45284 57588
rect 45336 57576 45342 57588
rect 63954 57576 63960 57588
rect 45336 57548 63960 57576
rect 45336 57536 45342 57548
rect 63954 57536 63960 57548
rect 64012 57536 64018 57588
rect 67266 57576 67272 57588
rect 67227 57548 67272 57576
rect 67266 57536 67272 57548
rect 67324 57536 67330 57588
rect 11698 57468 11704 57520
rect 11756 57508 11762 57520
rect 17313 57511 17371 57517
rect 17313 57508 17325 57511
rect 11756 57480 17325 57508
rect 11756 57468 11762 57480
rect 17313 57477 17325 57480
rect 17359 57477 17371 57511
rect 17313 57471 17371 57477
rect 36170 57468 36176 57520
rect 36228 57508 36234 57520
rect 51442 57508 51448 57520
rect 36228 57480 51448 57508
rect 36228 57468 36234 57480
rect 51442 57468 51448 57480
rect 51500 57468 51506 57520
rect 8846 57400 8852 57452
rect 8904 57440 8910 57452
rect 35621 57443 35679 57449
rect 35621 57440 35633 57443
rect 8904 57412 35633 57440
rect 8904 57400 8910 57412
rect 35621 57409 35633 57412
rect 35667 57409 35679 57443
rect 35621 57403 35679 57409
rect 1578 57372 1584 57384
rect 1539 57344 1584 57372
rect 1578 57332 1584 57344
rect 1636 57372 1642 57384
rect 2041 57375 2099 57381
rect 2041 57372 2053 57375
rect 1636 57344 2053 57372
rect 1636 57332 1642 57344
rect 2041 57341 2053 57344
rect 2087 57341 2099 57375
rect 25498 57372 25504 57384
rect 25459 57344 25504 57372
rect 2041 57335 2099 57341
rect 25498 57332 25504 57344
rect 25556 57332 25562 57384
rect 67266 57332 67272 57384
rect 67324 57372 67330 57384
rect 67913 57375 67971 57381
rect 67913 57372 67925 57375
rect 67324 57344 67925 57372
rect 67324 57332 67330 57344
rect 67913 57341 67925 57344
rect 67959 57341 67971 57375
rect 67913 57335 67971 57341
rect 68094 57304 68100 57316
rect 68055 57276 68100 57304
rect 68094 57264 68100 57276
rect 68152 57264 68158 57316
rect 6362 57196 6368 57248
rect 6420 57236 6426 57248
rect 6917 57239 6975 57245
rect 6917 57236 6929 57239
rect 6420 57208 6929 57236
rect 6420 57196 6426 57208
rect 6917 57205 6929 57208
rect 6963 57236 6975 57239
rect 18322 57236 18328 57248
rect 6963 57208 18328 57236
rect 6963 57205 6975 57208
rect 6917 57199 6975 57205
rect 18322 57196 18328 57208
rect 18380 57196 18386 57248
rect 50246 57196 50252 57248
rect 50304 57236 50310 57248
rect 66162 57236 66168 57248
rect 50304 57208 66168 57236
rect 50304 57196 50310 57208
rect 66162 57196 66168 57208
rect 66220 57196 66226 57248
rect 1104 57146 68816 57168
rect 1104 57094 9246 57146
rect 9298 57094 9310 57146
rect 9362 57094 9374 57146
rect 9426 57094 9438 57146
rect 9490 57094 19246 57146
rect 19298 57094 19310 57146
rect 19362 57094 19374 57146
rect 19426 57094 19438 57146
rect 19490 57094 29246 57146
rect 29298 57094 29310 57146
rect 29362 57094 29374 57146
rect 29426 57094 29438 57146
rect 29490 57094 39246 57146
rect 39298 57094 39310 57146
rect 39362 57094 39374 57146
rect 39426 57094 39438 57146
rect 39490 57094 49246 57146
rect 49298 57094 49310 57146
rect 49362 57094 49374 57146
rect 49426 57094 49438 57146
rect 49490 57094 59246 57146
rect 59298 57094 59310 57146
rect 59362 57094 59374 57146
rect 59426 57094 59438 57146
rect 59490 57094 68816 57146
rect 1104 57072 68816 57094
rect 10781 56695 10839 56701
rect 10781 56661 10793 56695
rect 10827 56692 10839 56695
rect 12618 56692 12624 56704
rect 10827 56664 12624 56692
rect 10827 56661 10839 56664
rect 10781 56655 10839 56661
rect 12618 56652 12624 56664
rect 12676 56652 12682 56704
rect 1104 56602 68816 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 14246 56602
rect 14298 56550 14310 56602
rect 14362 56550 14374 56602
rect 14426 56550 14438 56602
rect 14490 56550 24246 56602
rect 24298 56550 24310 56602
rect 24362 56550 24374 56602
rect 24426 56550 24438 56602
rect 24490 56550 34246 56602
rect 34298 56550 34310 56602
rect 34362 56550 34374 56602
rect 34426 56550 34438 56602
rect 34490 56550 44246 56602
rect 44298 56550 44310 56602
rect 44362 56550 44374 56602
rect 44426 56550 44438 56602
rect 44490 56550 54246 56602
rect 54298 56550 54310 56602
rect 54362 56550 54374 56602
rect 54426 56550 54438 56602
rect 54490 56550 64246 56602
rect 64298 56550 64310 56602
rect 64362 56550 64374 56602
rect 64426 56550 64438 56602
rect 64490 56550 68816 56602
rect 1104 56528 68816 56550
rect 1762 56352 1768 56364
rect 1723 56324 1768 56352
rect 1762 56312 1768 56324
rect 1820 56312 1826 56364
rect 26206 56324 35894 56352
rect 18233 56287 18291 56293
rect 18233 56253 18245 56287
rect 18279 56284 18291 56287
rect 26206 56284 26234 56324
rect 30282 56284 30288 56296
rect 18279 56256 26234 56284
rect 30243 56256 30288 56284
rect 18279 56253 18291 56256
rect 18233 56247 18291 56253
rect 30282 56244 30288 56256
rect 30340 56244 30346 56296
rect 35866 56284 35894 56324
rect 44634 56284 44640 56296
rect 35866 56256 44640 56284
rect 44634 56244 44640 56256
rect 44692 56244 44698 56296
rect 67453 56287 67511 56293
rect 67453 56253 67465 56287
rect 67499 56284 67511 56287
rect 68094 56284 68100 56296
rect 67499 56256 68100 56284
rect 67499 56253 67511 56256
rect 67453 56247 67511 56253
rect 68094 56244 68100 56256
rect 68152 56244 68158 56296
rect 1949 56219 2007 56225
rect 1949 56185 1961 56219
rect 1995 56185 2007 56219
rect 1949 56179 2007 56185
rect 1964 56148 1992 56179
rect 2498 56148 2504 56160
rect 1964 56120 2504 56148
rect 2498 56108 2504 56120
rect 2556 56108 2562 56160
rect 1104 56058 68816 56080
rect 1104 56006 9246 56058
rect 9298 56006 9310 56058
rect 9362 56006 9374 56058
rect 9426 56006 9438 56058
rect 9490 56006 19246 56058
rect 19298 56006 19310 56058
rect 19362 56006 19374 56058
rect 19426 56006 19438 56058
rect 19490 56006 29246 56058
rect 29298 56006 29310 56058
rect 29362 56006 29374 56058
rect 29426 56006 29438 56058
rect 29490 56006 39246 56058
rect 39298 56006 39310 56058
rect 39362 56006 39374 56058
rect 39426 56006 39438 56058
rect 39490 56006 49246 56058
rect 49298 56006 49310 56058
rect 49362 56006 49374 56058
rect 49426 56006 49438 56058
rect 49490 56006 59246 56058
rect 59298 56006 59310 56058
rect 59362 56006 59374 56058
rect 59426 56006 59438 56058
rect 59490 56006 68816 56058
rect 1104 55984 68816 56006
rect 6886 55848 16574 55876
rect 2682 55632 2688 55684
rect 2740 55672 2746 55684
rect 6886 55672 6914 55848
rect 9950 55808 9956 55820
rect 9911 55780 9956 55808
rect 9950 55768 9956 55780
rect 10008 55768 10014 55820
rect 10045 55743 10103 55749
rect 10045 55709 10057 55743
rect 10091 55740 10103 55743
rect 10091 55712 13308 55740
rect 10091 55709 10103 55712
rect 10045 55703 10103 55709
rect 2740 55644 6914 55672
rect 2740 55632 2746 55644
rect 11054 55604 11060 55616
rect 11015 55576 11060 55604
rect 11054 55564 11060 55576
rect 11112 55564 11118 55616
rect 13078 55604 13084 55616
rect 13039 55576 13084 55604
rect 13078 55564 13084 55576
rect 13136 55564 13142 55616
rect 13280 55604 13308 55712
rect 16546 55672 16574 55848
rect 31294 55836 31300 55888
rect 31352 55876 31358 55888
rect 51626 55876 51632 55888
rect 31352 55848 51632 55876
rect 31352 55836 31358 55848
rect 51626 55836 51632 55848
rect 51684 55836 51690 55888
rect 25498 55672 25504 55684
rect 16546 55644 25504 55672
rect 25498 55632 25504 55644
rect 25556 55632 25562 55684
rect 47578 55672 47584 55684
rect 26206 55644 47584 55672
rect 26206 55604 26234 55644
rect 47578 55632 47584 55644
rect 47636 55632 47642 55684
rect 38010 55604 38016 55616
rect 13280 55576 26234 55604
rect 37971 55576 38016 55604
rect 38010 55564 38016 55576
rect 38068 55564 38074 55616
rect 1104 55514 68816 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 14246 55514
rect 14298 55462 14310 55514
rect 14362 55462 14374 55514
rect 14426 55462 14438 55514
rect 14490 55462 24246 55514
rect 24298 55462 24310 55514
rect 24362 55462 24374 55514
rect 24426 55462 24438 55514
rect 24490 55462 34246 55514
rect 34298 55462 34310 55514
rect 34362 55462 34374 55514
rect 34426 55462 34438 55514
rect 34490 55462 44246 55514
rect 44298 55462 44310 55514
rect 44362 55462 44374 55514
rect 44426 55462 44438 55514
rect 44490 55462 54246 55514
rect 54298 55462 54310 55514
rect 54362 55462 54374 55514
rect 54426 55462 54438 55514
rect 54490 55462 64246 55514
rect 64298 55462 64310 55514
rect 64362 55462 64374 55514
rect 64426 55462 64438 55514
rect 64490 55462 68816 55514
rect 1104 55440 68816 55462
rect 11054 55360 11060 55412
rect 11112 55400 11118 55412
rect 42334 55400 42340 55412
rect 11112 55372 42340 55400
rect 11112 55360 11118 55372
rect 42334 55360 42340 55372
rect 42392 55360 42398 55412
rect 9950 55292 9956 55344
rect 10008 55332 10014 55344
rect 10229 55335 10287 55341
rect 10229 55332 10241 55335
rect 10008 55304 10241 55332
rect 10008 55292 10014 55304
rect 10229 55301 10241 55304
rect 10275 55332 10287 55335
rect 31294 55332 31300 55344
rect 10275 55304 31300 55332
rect 10275 55301 10287 55304
rect 10229 55295 10287 55301
rect 31294 55292 31300 55304
rect 31352 55292 31358 55344
rect 37369 55335 37427 55341
rect 37369 55301 37381 55335
rect 37415 55332 37427 55335
rect 38749 55335 38807 55341
rect 38749 55332 38761 55335
rect 37415 55304 38761 55332
rect 37415 55301 37427 55304
rect 37369 55295 37427 55301
rect 38749 55301 38761 55304
rect 38795 55332 38807 55335
rect 39942 55332 39948 55344
rect 38795 55304 39948 55332
rect 38795 55301 38807 55304
rect 38749 55295 38807 55301
rect 39942 55292 39948 55304
rect 40000 55292 40006 55344
rect 61105 55335 61163 55341
rect 61105 55301 61117 55335
rect 61151 55332 61163 55335
rect 67450 55332 67456 55344
rect 61151 55304 67456 55332
rect 61151 55301 61163 55304
rect 61105 55295 61163 55301
rect 67450 55292 67456 55304
rect 67508 55292 67514 55344
rect 2593 55267 2651 55273
rect 2593 55264 2605 55267
rect 2503 55236 2605 55264
rect 2593 55233 2605 55236
rect 2639 55264 2651 55267
rect 2682 55264 2688 55276
rect 2639 55236 2688 55264
rect 2639 55233 2651 55236
rect 2593 55227 2651 55233
rect 1949 55199 2007 55205
rect 1949 55165 1961 55199
rect 1995 55196 2007 55199
rect 2608 55196 2636 55227
rect 2682 55224 2688 55236
rect 2740 55224 2746 55276
rect 38856 55236 39620 55264
rect 1995 55168 2636 55196
rect 1995 55165 2007 55168
rect 1949 55159 2007 55165
rect 38010 55156 38016 55208
rect 38068 55196 38074 55208
rect 38565 55199 38623 55205
rect 38565 55196 38577 55199
rect 38068 55168 38577 55196
rect 38068 55156 38074 55168
rect 38565 55165 38577 55168
rect 38611 55165 38623 55199
rect 38565 55159 38623 55165
rect 38657 55199 38715 55205
rect 38657 55165 38669 55199
rect 38703 55196 38715 55199
rect 38746 55196 38752 55208
rect 38703 55168 38752 55196
rect 38703 55165 38715 55168
rect 38657 55159 38715 55165
rect 38746 55156 38752 55168
rect 38804 55156 38810 55208
rect 38856 55205 38884 55236
rect 38841 55199 38899 55205
rect 38841 55165 38853 55199
rect 38887 55196 38899 55199
rect 39025 55199 39083 55205
rect 38887 55168 38921 55196
rect 38887 55165 38899 55168
rect 38841 55159 38899 55165
rect 39025 55165 39037 55199
rect 39071 55165 39083 55199
rect 39025 55159 39083 55165
rect 37458 55088 37464 55140
rect 37516 55128 37522 55140
rect 39040 55128 39068 55159
rect 39592 55137 39620 55236
rect 41690 55224 41696 55276
rect 41748 55264 41754 55276
rect 41969 55267 42027 55273
rect 41969 55264 41981 55267
rect 41748 55236 41981 55264
rect 41748 55224 41754 55236
rect 41969 55233 41981 55236
rect 42015 55233 42027 55267
rect 41969 55227 42027 55233
rect 67082 55224 67088 55276
rect 67140 55264 67146 55276
rect 67177 55267 67235 55273
rect 67177 55264 67189 55267
rect 67140 55236 67189 55264
rect 67140 55224 67146 55236
rect 67177 55233 67189 55236
rect 67223 55233 67235 55267
rect 67177 55227 67235 55233
rect 39577 55131 39635 55137
rect 39577 55128 39589 55131
rect 37516 55100 39068 55128
rect 39487 55100 39589 55128
rect 37516 55088 37522 55100
rect 39577 55097 39589 55100
rect 39623 55097 39635 55131
rect 39577 55091 39635 55097
rect 1854 55060 1860 55072
rect 1815 55032 1860 55060
rect 1854 55020 1860 55032
rect 1912 55020 1918 55072
rect 38378 55060 38384 55072
rect 38339 55032 38384 55060
rect 38378 55020 38384 55032
rect 38436 55020 38442 55072
rect 39592 55060 39620 55091
rect 62758 55060 62764 55072
rect 39592 55032 62764 55060
rect 62758 55020 62764 55032
rect 62816 55020 62822 55072
rect 1104 54970 68816 54992
rect 1104 54918 9246 54970
rect 9298 54918 9310 54970
rect 9362 54918 9374 54970
rect 9426 54918 9438 54970
rect 9490 54918 19246 54970
rect 19298 54918 19310 54970
rect 19362 54918 19374 54970
rect 19426 54918 19438 54970
rect 19490 54918 29246 54970
rect 29298 54918 29310 54970
rect 29362 54918 29374 54970
rect 29426 54918 29438 54970
rect 29490 54918 39246 54970
rect 39298 54918 39310 54970
rect 39362 54918 39374 54970
rect 39426 54918 39438 54970
rect 39490 54918 49246 54970
rect 49298 54918 49310 54970
rect 49362 54918 49374 54970
rect 49426 54918 49438 54970
rect 49490 54918 59246 54970
rect 59298 54918 59310 54970
rect 59362 54918 59374 54970
rect 59426 54918 59438 54970
rect 59490 54918 68816 54970
rect 1104 54896 68816 54918
rect 33870 54476 33876 54528
rect 33928 54516 33934 54528
rect 38105 54519 38163 54525
rect 38105 54516 38117 54519
rect 33928 54488 38117 54516
rect 33928 54476 33934 54488
rect 38105 54485 38117 54488
rect 38151 54516 38163 54519
rect 38746 54516 38752 54528
rect 38151 54488 38752 54516
rect 38151 54485 38163 54488
rect 38105 54479 38163 54485
rect 38746 54476 38752 54488
rect 38804 54476 38810 54528
rect 44818 54516 44824 54528
rect 44779 54488 44824 54516
rect 44818 54476 44824 54488
rect 44876 54476 44882 54528
rect 62114 54516 62120 54528
rect 62075 54488 62120 54516
rect 62114 54476 62120 54488
rect 62172 54476 62178 54528
rect 1104 54426 68816 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 14246 54426
rect 14298 54374 14310 54426
rect 14362 54374 14374 54426
rect 14426 54374 14438 54426
rect 14490 54374 24246 54426
rect 24298 54374 24310 54426
rect 24362 54374 24374 54426
rect 24426 54374 24438 54426
rect 24490 54374 34246 54426
rect 34298 54374 34310 54426
rect 34362 54374 34374 54426
rect 34426 54374 34438 54426
rect 34490 54374 44246 54426
rect 44298 54374 44310 54426
rect 44362 54374 44374 54426
rect 44426 54374 44438 54426
rect 44490 54374 54246 54426
rect 54298 54374 54310 54426
rect 54362 54374 54374 54426
rect 54426 54374 54438 54426
rect 54490 54374 64246 54426
rect 64298 54374 64310 54426
rect 64362 54374 64374 54426
rect 64426 54374 64438 54426
rect 64490 54374 68816 54426
rect 1104 54352 68816 54374
rect 2406 54272 2412 54324
rect 2464 54312 2470 54324
rect 44818 54312 44824 54324
rect 2464 54284 44824 54312
rect 2464 54272 2470 54284
rect 44818 54272 44824 54284
rect 44876 54272 44882 54324
rect 45526 54148 55214 54176
rect 5629 54111 5687 54117
rect 5629 54077 5641 54111
rect 5675 54108 5687 54111
rect 45526 54108 45554 54148
rect 48774 54108 48780 54120
rect 5675 54080 45554 54108
rect 48735 54080 48780 54108
rect 5675 54077 5687 54080
rect 5629 54071 5687 54077
rect 48774 54068 48780 54080
rect 48832 54068 48838 54120
rect 55186 54108 55214 54148
rect 66898 54108 66904 54120
rect 55186 54080 66904 54108
rect 66898 54068 66904 54080
rect 66956 54068 66962 54120
rect 1104 53882 68816 53904
rect 1104 53830 9246 53882
rect 9298 53830 9310 53882
rect 9362 53830 9374 53882
rect 9426 53830 9438 53882
rect 9490 53830 19246 53882
rect 19298 53830 19310 53882
rect 19362 53830 19374 53882
rect 19426 53830 19438 53882
rect 19490 53830 29246 53882
rect 29298 53830 29310 53882
rect 29362 53830 29374 53882
rect 29426 53830 29438 53882
rect 29490 53830 39246 53882
rect 39298 53830 39310 53882
rect 39362 53830 39374 53882
rect 39426 53830 39438 53882
rect 39490 53830 49246 53882
rect 49298 53830 49310 53882
rect 49362 53830 49374 53882
rect 49426 53830 49438 53882
rect 49490 53830 59246 53882
rect 59298 53830 59310 53882
rect 59362 53830 59374 53882
rect 59426 53830 59438 53882
rect 59490 53830 68816 53882
rect 1104 53808 68816 53830
rect 33321 53771 33379 53777
rect 33321 53737 33333 53771
rect 33367 53768 33379 53771
rect 37458 53768 37464 53780
rect 33367 53740 37464 53768
rect 33367 53737 33379 53740
rect 33321 53731 33379 53737
rect 37458 53728 37464 53740
rect 37516 53728 37522 53780
rect 32309 53703 32367 53709
rect 32309 53700 32321 53703
rect 28736 53672 32321 53700
rect 28736 53641 28764 53672
rect 32309 53669 32321 53672
rect 32355 53700 32367 53703
rect 32355 53672 35894 53700
rect 32355 53669 32367 53672
rect 32309 53663 32367 53669
rect 28077 53635 28135 53641
rect 28077 53632 28089 53635
rect 26206 53604 28089 53632
rect 7745 53431 7803 53437
rect 7745 53397 7757 53431
rect 7791 53428 7803 53431
rect 12158 53428 12164 53440
rect 7791 53400 12164 53428
rect 7791 53397 7803 53400
rect 7745 53391 7803 53397
rect 12158 53388 12164 53400
rect 12216 53388 12222 53440
rect 19978 53388 19984 53440
rect 20036 53428 20042 53440
rect 26206 53428 26234 53604
rect 28077 53601 28089 53604
rect 28123 53632 28135 53635
rect 28721 53635 28779 53641
rect 28721 53632 28733 53635
rect 28123 53604 28733 53632
rect 28123 53601 28135 53604
rect 28077 53595 28135 53601
rect 28721 53601 28733 53604
rect 28767 53601 28779 53635
rect 28721 53595 28779 53601
rect 29086 53524 29092 53576
rect 29144 53564 29150 53576
rect 29365 53567 29423 53573
rect 29365 53564 29377 53567
rect 29144 53536 29377 53564
rect 29144 53524 29150 53536
rect 29365 53533 29377 53536
rect 29411 53564 29423 53567
rect 29546 53564 29552 53576
rect 29411 53536 29552 53564
rect 29411 53533 29423 53536
rect 29365 53527 29423 53533
rect 29546 53524 29552 53536
rect 29604 53524 29610 53576
rect 32858 53564 32864 53576
rect 32819 53536 32864 53564
rect 32858 53524 32864 53536
rect 32916 53524 32922 53576
rect 32968 53573 32996 53672
rect 33045 53635 33103 53641
rect 33045 53601 33057 53635
rect 33091 53632 33103 53635
rect 35866 53632 35894 53672
rect 43254 53632 43260 53644
rect 33091 53604 33548 53632
rect 35866 53604 43260 53632
rect 33091 53601 33103 53604
rect 33045 53595 33103 53601
rect 32953 53567 33011 53573
rect 32953 53533 32965 53567
rect 32999 53533 33011 53567
rect 33134 53564 33140 53576
rect 33095 53536 33140 53564
rect 32953 53527 33011 53533
rect 33134 53524 33140 53536
rect 33192 53524 33198 53576
rect 31757 53499 31815 53505
rect 31757 53465 31769 53499
rect 31803 53496 31815 53499
rect 33244 53496 33272 53604
rect 33520 53564 33548 53604
rect 43254 53592 43260 53604
rect 43312 53592 43318 53644
rect 67913 53635 67971 53641
rect 67913 53632 67925 53635
rect 67284 53604 67925 53632
rect 33520 53536 35894 53564
rect 31803 53468 33272 53496
rect 31803 53465 31815 53468
rect 31757 53459 31815 53465
rect 20036 53400 26234 53428
rect 35866 53428 35894 53536
rect 37182 53428 37188 53440
rect 35866 53400 37188 53428
rect 20036 53388 20042 53400
rect 37182 53388 37188 53400
rect 37240 53428 37246 53440
rect 43438 53428 43444 53440
rect 37240 53400 43444 53428
rect 37240 53388 37246 53400
rect 43438 53388 43444 53400
rect 43496 53388 43502 53440
rect 53926 53428 53932 53440
rect 53887 53400 53932 53428
rect 53926 53388 53932 53400
rect 53984 53388 53990 53440
rect 55493 53431 55551 53437
rect 55493 53397 55505 53431
rect 55539 53428 55551 53431
rect 55582 53428 55588 53440
rect 55539 53400 55588 53428
rect 55539 53397 55551 53400
rect 55493 53391 55551 53397
rect 55582 53388 55588 53400
rect 55640 53388 55646 53440
rect 55858 53388 55864 53440
rect 55916 53428 55922 53440
rect 67284 53437 67312 53604
rect 67913 53601 67925 53604
rect 67959 53601 67971 53635
rect 67913 53595 67971 53601
rect 68094 53496 68100 53508
rect 68055 53468 68100 53496
rect 68094 53456 68100 53468
rect 68152 53456 68158 53508
rect 67269 53431 67327 53437
rect 67269 53428 67281 53431
rect 55916 53400 67281 53428
rect 55916 53388 55922 53400
rect 67269 53397 67281 53400
rect 67315 53397 67327 53431
rect 67269 53391 67327 53397
rect 1104 53338 68816 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 14246 53338
rect 14298 53286 14310 53338
rect 14362 53286 14374 53338
rect 14426 53286 14438 53338
rect 14490 53286 24246 53338
rect 24298 53286 24310 53338
rect 24362 53286 24374 53338
rect 24426 53286 24438 53338
rect 24490 53286 34246 53338
rect 34298 53286 34310 53338
rect 34362 53286 34374 53338
rect 34426 53286 34438 53338
rect 34490 53286 44246 53338
rect 44298 53286 44310 53338
rect 44362 53286 44374 53338
rect 44426 53286 44438 53338
rect 44490 53286 54246 53338
rect 54298 53286 54310 53338
rect 54362 53286 54374 53338
rect 54426 53286 54438 53338
rect 54490 53286 64246 53338
rect 64298 53286 64310 53338
rect 64362 53286 64374 53338
rect 64426 53286 64438 53338
rect 64490 53286 68816 53338
rect 1104 53264 68816 53286
rect 2682 53184 2688 53236
rect 2740 53224 2746 53236
rect 55769 53227 55827 53233
rect 55769 53224 55781 53227
rect 2740 53196 55781 53224
rect 2740 53184 2746 53196
rect 55769 53193 55781 53196
rect 55815 53193 55827 53227
rect 55769 53187 55827 53193
rect 53926 53116 53932 53168
rect 53984 53156 53990 53168
rect 54665 53159 54723 53165
rect 54665 53156 54677 53159
rect 53984 53128 54677 53156
rect 53984 53116 53990 53128
rect 54665 53125 54677 53128
rect 54711 53125 54723 53159
rect 54665 53119 54723 53125
rect 40681 53091 40739 53097
rect 40681 53057 40693 53091
rect 40727 53088 40739 53091
rect 66346 53088 66352 53100
rect 40727 53060 66352 53088
rect 40727 53057 40739 53060
rect 40681 53051 40739 53057
rect 66346 53048 66352 53060
rect 66404 53048 66410 53100
rect 41325 53023 41383 53029
rect 41325 52989 41337 53023
rect 41371 53020 41383 53023
rect 45094 53020 45100 53032
rect 41371 52992 45100 53020
rect 41371 52989 41383 52992
rect 41325 52983 41383 52989
rect 45094 52980 45100 52992
rect 45152 52980 45158 53032
rect 51077 53023 51135 53029
rect 51077 52989 51089 53023
rect 51123 53020 51135 53023
rect 51994 53020 52000 53032
rect 51123 52992 52000 53020
rect 51123 52989 51135 52992
rect 51077 52983 51135 52989
rect 51994 52980 52000 52992
rect 52052 52980 52058 53032
rect 53006 52980 53012 53032
rect 53064 53020 53070 53032
rect 54389 53023 54447 53029
rect 54389 53020 54401 53023
rect 53064 52992 54401 53020
rect 53064 52980 53070 52992
rect 54389 52989 54401 52992
rect 54435 52989 54447 53023
rect 54570 53020 54576 53032
rect 54531 52992 54576 53020
rect 54389 52983 54447 52989
rect 54570 52980 54576 52992
rect 54628 52980 54634 53032
rect 54662 52980 54668 53032
rect 54720 53020 54726 53032
rect 54757 53023 54815 53029
rect 54757 53020 54769 53023
rect 54720 52992 54769 53020
rect 54720 52980 54726 52992
rect 54757 52989 54769 52992
rect 54803 52989 54815 53023
rect 54757 52983 54815 52989
rect 54849 53023 54907 53029
rect 54849 52989 54861 53023
rect 54895 53020 54907 53023
rect 55582 53020 55588 53032
rect 54895 52992 55168 53020
rect 55543 52992 55588 53020
rect 54895 52989 54907 52992
rect 54849 52983 54907 52989
rect 32125 52955 32183 52961
rect 32125 52921 32137 52955
rect 32171 52952 32183 52955
rect 32858 52952 32864 52964
rect 32171 52924 32864 52952
rect 32171 52921 32183 52924
rect 32125 52915 32183 52921
rect 32858 52912 32864 52924
rect 32916 52912 32922 52964
rect 36906 52912 36912 52964
rect 36964 52952 36970 52964
rect 55033 52955 55091 52961
rect 55033 52952 55045 52955
rect 36964 52924 55045 52952
rect 36964 52912 36970 52924
rect 55033 52921 55045 52924
rect 55079 52921 55091 52955
rect 55033 52915 55091 52921
rect 32769 52887 32827 52893
rect 32769 52853 32781 52887
rect 32815 52884 32827 52887
rect 33134 52884 33140 52896
rect 32815 52856 33140 52884
rect 32815 52853 32827 52856
rect 32769 52847 32827 52853
rect 33134 52844 33140 52856
rect 33192 52844 33198 52896
rect 53006 52884 53012 52896
rect 52967 52856 53012 52884
rect 53006 52844 53012 52856
rect 53064 52844 53070 52896
rect 53834 52884 53840 52896
rect 53795 52856 53840 52884
rect 53834 52844 53840 52856
rect 53892 52884 53898 52896
rect 55140 52884 55168 52992
rect 55582 52980 55588 52992
rect 55640 52980 55646 53032
rect 62850 53020 62856 53032
rect 62811 52992 62856 53020
rect 62850 52980 62856 52992
rect 62908 52980 62914 53032
rect 65242 53020 65248 53032
rect 65203 52992 65248 53020
rect 65242 52980 65248 52992
rect 65300 52980 65306 53032
rect 62758 52952 62764 52964
rect 62719 52924 62764 52952
rect 62758 52912 62764 52924
rect 62816 52912 62822 52964
rect 53892 52856 55168 52884
rect 53892 52844 53898 52856
rect 1104 52794 68816 52816
rect 1104 52742 9246 52794
rect 9298 52742 9310 52794
rect 9362 52742 9374 52794
rect 9426 52742 9438 52794
rect 9490 52742 19246 52794
rect 19298 52742 19310 52794
rect 19362 52742 19374 52794
rect 19426 52742 19438 52794
rect 19490 52742 29246 52794
rect 29298 52742 29310 52794
rect 29362 52742 29374 52794
rect 29426 52742 29438 52794
rect 29490 52742 39246 52794
rect 39298 52742 39310 52794
rect 39362 52742 39374 52794
rect 39426 52742 39438 52794
rect 39490 52742 49246 52794
rect 49298 52742 49310 52794
rect 49362 52742 49374 52794
rect 49426 52742 49438 52794
rect 49490 52742 59246 52794
rect 59298 52742 59310 52794
rect 59362 52742 59374 52794
rect 59426 52742 59438 52794
rect 59490 52742 68816 52794
rect 1104 52720 68816 52742
rect 39942 52640 39948 52692
rect 40000 52680 40006 52692
rect 48222 52680 48228 52692
rect 40000 52652 48228 52680
rect 40000 52640 40006 52652
rect 48222 52640 48228 52652
rect 48280 52680 48286 52692
rect 55582 52680 55588 52692
rect 48280 52652 55588 52680
rect 48280 52640 48286 52652
rect 55582 52640 55588 52652
rect 55640 52640 55646 52692
rect 62390 52640 62396 52692
rect 62448 52680 62454 52692
rect 62850 52680 62856 52692
rect 62448 52652 62856 52680
rect 62448 52640 62454 52652
rect 62850 52640 62856 52652
rect 62908 52680 62914 52692
rect 63221 52683 63279 52689
rect 63221 52680 63233 52683
rect 62908 52652 63233 52680
rect 62908 52640 62914 52652
rect 63221 52649 63233 52652
rect 63267 52649 63279 52683
rect 63221 52643 63279 52649
rect 1578 52544 1584 52556
rect 1539 52516 1584 52544
rect 1578 52504 1584 52516
rect 1636 52544 1642 52556
rect 2041 52547 2099 52553
rect 2041 52544 2053 52547
rect 1636 52516 2053 52544
rect 1636 52504 1642 52516
rect 2041 52513 2053 52516
rect 2087 52513 2099 52547
rect 2041 52507 2099 52513
rect 11238 52504 11244 52556
rect 11296 52544 11302 52556
rect 53834 52544 53840 52556
rect 11296 52516 53840 52544
rect 11296 52504 11302 52516
rect 53834 52504 53840 52516
rect 53892 52504 53898 52556
rect 54662 52544 54668 52556
rect 54036 52516 54668 52544
rect 54036 52488 54064 52516
rect 54662 52504 54668 52516
rect 54720 52504 54726 52556
rect 19978 52436 19984 52488
rect 20036 52476 20042 52488
rect 20622 52476 20628 52488
rect 20036 52448 20628 52476
rect 20036 52436 20042 52448
rect 20622 52436 20628 52448
rect 20680 52436 20686 52488
rect 54018 52476 54024 52488
rect 53979 52448 54024 52476
rect 54018 52436 54024 52448
rect 54076 52436 54082 52488
rect 54570 52436 54576 52488
rect 54628 52476 54634 52488
rect 55306 52476 55312 52488
rect 54628 52448 55312 52476
rect 54628 52436 54634 52448
rect 55306 52436 55312 52448
rect 55364 52436 55370 52488
rect 65978 52408 65984 52420
rect 45526 52380 65984 52408
rect 27065 52343 27123 52349
rect 27065 52309 27077 52343
rect 27111 52340 27123 52343
rect 45526 52340 45554 52380
rect 65978 52368 65984 52380
rect 66036 52368 66042 52420
rect 27111 52312 45554 52340
rect 27111 52309 27123 52312
rect 27065 52303 27123 52309
rect 1104 52250 68816 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 14246 52250
rect 14298 52198 14310 52250
rect 14362 52198 14374 52250
rect 14426 52198 14438 52250
rect 14490 52198 24246 52250
rect 24298 52198 24310 52250
rect 24362 52198 24374 52250
rect 24426 52198 24438 52250
rect 24490 52198 34246 52250
rect 34298 52198 34310 52250
rect 34362 52198 34374 52250
rect 34426 52198 34438 52250
rect 34490 52198 44246 52250
rect 44298 52198 44310 52250
rect 44362 52198 44374 52250
rect 44426 52198 44438 52250
rect 44490 52198 54246 52250
rect 54298 52198 54310 52250
rect 54362 52198 54374 52250
rect 54426 52198 54438 52250
rect 54490 52198 64246 52250
rect 64298 52198 64310 52250
rect 64362 52198 64374 52250
rect 64426 52198 64438 52250
rect 64490 52198 68816 52250
rect 1104 52176 68816 52198
rect 67174 52096 67180 52148
rect 67232 52136 67238 52148
rect 67269 52139 67327 52145
rect 67269 52136 67281 52139
rect 67232 52108 67281 52136
rect 67232 52096 67238 52108
rect 67269 52105 67281 52108
rect 67315 52105 67327 52139
rect 67269 52099 67327 52105
rect 15838 51932 15844 51944
rect 15799 51904 15844 51932
rect 15838 51892 15844 51904
rect 15896 51892 15902 51944
rect 67284 51932 67312 52099
rect 68094 52000 68100 52012
rect 68055 51972 68100 52000
rect 68094 51960 68100 51972
rect 68152 51960 68158 52012
rect 67913 51935 67971 51941
rect 67913 51932 67925 51935
rect 67284 51904 67925 51932
rect 67913 51901 67925 51904
rect 67959 51901 67971 51935
rect 67913 51895 67971 51901
rect 31294 51756 31300 51808
rect 31352 51796 31358 51808
rect 32030 51796 32036 51808
rect 31352 51768 32036 51796
rect 31352 51756 31358 51768
rect 32030 51756 32036 51768
rect 32088 51796 32094 51808
rect 53926 51796 53932 51808
rect 32088 51768 53932 51796
rect 32088 51756 32094 51768
rect 53926 51756 53932 51768
rect 53984 51756 53990 51808
rect 1104 51706 68816 51728
rect 1104 51654 9246 51706
rect 9298 51654 9310 51706
rect 9362 51654 9374 51706
rect 9426 51654 9438 51706
rect 9490 51654 19246 51706
rect 19298 51654 19310 51706
rect 19362 51654 19374 51706
rect 19426 51654 19438 51706
rect 19490 51654 29246 51706
rect 29298 51654 29310 51706
rect 29362 51654 29374 51706
rect 29426 51654 29438 51706
rect 29490 51654 39246 51706
rect 39298 51654 39310 51706
rect 39362 51654 39374 51706
rect 39426 51654 39438 51706
rect 39490 51654 49246 51706
rect 49298 51654 49310 51706
rect 49362 51654 49374 51706
rect 49426 51654 49438 51706
rect 49490 51654 59246 51706
rect 59298 51654 59310 51706
rect 59362 51654 59374 51706
rect 59426 51654 59438 51706
rect 59490 51654 68816 51706
rect 1104 51632 68816 51654
rect 15289 51459 15347 51465
rect 15289 51425 15301 51459
rect 15335 51456 15347 51459
rect 15841 51459 15899 51465
rect 15841 51456 15853 51459
rect 15335 51428 15853 51456
rect 15335 51425 15347 51428
rect 15289 51419 15347 51425
rect 15841 51425 15853 51428
rect 15887 51456 15899 51459
rect 39942 51456 39948 51468
rect 15887 51428 39948 51456
rect 15887 51425 15899 51428
rect 15841 51419 15899 51425
rect 39942 51416 39948 51428
rect 40000 51416 40006 51468
rect 15105 51391 15163 51397
rect 15105 51357 15117 51391
rect 15151 51388 15163 51391
rect 31294 51388 31300 51400
rect 15151 51360 31300 51388
rect 15151 51357 15163 51360
rect 15105 51351 15163 51357
rect 31294 51348 31300 51360
rect 31352 51348 31358 51400
rect 31481 51391 31539 51397
rect 31481 51357 31493 51391
rect 31527 51388 31539 51391
rect 46198 51388 46204 51400
rect 31527 51360 35894 51388
rect 46159 51360 46204 51388
rect 31527 51357 31539 51360
rect 31481 51351 31539 51357
rect 35866 51320 35894 51360
rect 46198 51348 46204 51360
rect 46256 51348 46262 51400
rect 66438 51320 66444 51332
rect 6886 51292 16574 51320
rect 2498 51212 2504 51264
rect 2556 51252 2562 51264
rect 6886 51252 6914 51292
rect 2556 51224 6914 51252
rect 16546 51252 16574 51292
rect 26206 51292 31616 51320
rect 35866 51292 66444 51320
rect 26206 51252 26234 51292
rect 16546 51224 26234 51252
rect 31588 51252 31616 51292
rect 66438 51280 66444 51292
rect 66496 51280 66502 51332
rect 67361 51255 67419 51261
rect 67361 51252 67373 51255
rect 31588 51224 67373 51252
rect 2556 51212 2562 51224
rect 67361 51221 67373 51224
rect 67407 51221 67419 51255
rect 67361 51215 67419 51221
rect 1104 51162 68816 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 14246 51162
rect 14298 51110 14310 51162
rect 14362 51110 14374 51162
rect 14426 51110 14438 51162
rect 14490 51110 24246 51162
rect 24298 51110 24310 51162
rect 24362 51110 24374 51162
rect 24426 51110 24438 51162
rect 24490 51110 34246 51162
rect 34298 51110 34310 51162
rect 34362 51110 34374 51162
rect 34426 51110 34438 51162
rect 34490 51110 44246 51162
rect 44298 51110 44310 51162
rect 44362 51110 44374 51162
rect 44426 51110 44438 51162
rect 44490 51110 54246 51162
rect 54298 51110 54310 51162
rect 54362 51110 54374 51162
rect 54426 51110 54438 51162
rect 54490 51110 64246 51162
rect 64298 51110 64310 51162
rect 64362 51110 64374 51162
rect 64426 51110 64438 51162
rect 64490 51110 68816 51162
rect 1104 51088 68816 51110
rect 1854 51048 1860 51060
rect 1815 51020 1860 51048
rect 1854 51008 1860 51020
rect 1912 51008 1918 51060
rect 2593 51051 2651 51057
rect 2593 51017 2605 51051
rect 2639 51048 2651 51051
rect 2682 51048 2688 51060
rect 2639 51020 2688 51048
rect 2639 51017 2651 51020
rect 2593 51011 2651 51017
rect 1949 50847 2007 50853
rect 1949 50813 1961 50847
rect 1995 50844 2007 50847
rect 2608 50844 2636 51011
rect 2682 51008 2688 51020
rect 2740 51008 2746 51060
rect 16574 50872 16580 50924
rect 16632 50912 16638 50924
rect 34425 50915 34483 50921
rect 34425 50912 34437 50915
rect 16632 50884 34437 50912
rect 16632 50872 16638 50884
rect 34425 50881 34437 50884
rect 34471 50881 34483 50915
rect 34425 50875 34483 50881
rect 1995 50816 2636 50844
rect 17957 50847 18015 50853
rect 1995 50813 2007 50816
rect 1949 50807 2007 50813
rect 17957 50813 17969 50847
rect 18003 50844 18015 50847
rect 54205 50847 54263 50853
rect 18003 50816 18644 50844
rect 18003 50813 18015 50816
rect 17957 50807 18015 50813
rect 17589 50779 17647 50785
rect 17589 50745 17601 50779
rect 17635 50776 17647 50779
rect 17862 50776 17868 50788
rect 17635 50748 17868 50776
rect 17635 50745 17647 50748
rect 17589 50739 17647 50745
rect 17862 50736 17868 50748
rect 17920 50736 17926 50788
rect 18616 50717 18644 50816
rect 54205 50813 54217 50847
rect 54251 50844 54263 50847
rect 55950 50844 55956 50856
rect 54251 50816 55956 50844
rect 54251 50813 54263 50816
rect 54205 50807 54263 50813
rect 55950 50804 55956 50816
rect 56008 50804 56014 50856
rect 67453 50847 67511 50853
rect 67453 50813 67465 50847
rect 67499 50844 67511 50847
rect 68094 50844 68100 50856
rect 67499 50816 68100 50844
rect 67499 50813 67511 50816
rect 67453 50807 67511 50813
rect 68094 50804 68100 50816
rect 68152 50804 68158 50856
rect 18601 50711 18659 50717
rect 18601 50677 18613 50711
rect 18647 50708 18659 50711
rect 49602 50708 49608 50720
rect 18647 50680 49608 50708
rect 18647 50677 18659 50680
rect 18601 50671 18659 50677
rect 49602 50668 49608 50680
rect 49660 50708 49666 50720
rect 50430 50708 50436 50720
rect 49660 50680 50436 50708
rect 49660 50668 49666 50680
rect 50430 50668 50436 50680
rect 50488 50668 50494 50720
rect 1104 50618 68816 50640
rect 1104 50566 9246 50618
rect 9298 50566 9310 50618
rect 9362 50566 9374 50618
rect 9426 50566 9438 50618
rect 9490 50566 19246 50618
rect 19298 50566 19310 50618
rect 19362 50566 19374 50618
rect 19426 50566 19438 50618
rect 19490 50566 29246 50618
rect 29298 50566 29310 50618
rect 29362 50566 29374 50618
rect 29426 50566 29438 50618
rect 29490 50566 39246 50618
rect 39298 50566 39310 50618
rect 39362 50566 39374 50618
rect 39426 50566 39438 50618
rect 39490 50566 49246 50618
rect 49298 50566 49310 50618
rect 49362 50566 49374 50618
rect 49426 50566 49438 50618
rect 49490 50566 59246 50618
rect 59298 50566 59310 50618
rect 59362 50566 59374 50618
rect 59426 50566 59438 50618
rect 59490 50566 68816 50618
rect 1104 50544 68816 50566
rect 30926 50328 30932 50380
rect 30984 50368 30990 50380
rect 54018 50368 54024 50380
rect 30984 50340 54024 50368
rect 30984 50328 30990 50340
rect 54018 50328 54024 50340
rect 54076 50328 54082 50380
rect 34146 50192 34152 50244
rect 34204 50232 34210 50244
rect 34425 50235 34483 50241
rect 34425 50232 34437 50235
rect 34204 50204 34437 50232
rect 34204 50192 34210 50204
rect 34425 50201 34437 50204
rect 34471 50201 34483 50235
rect 34425 50195 34483 50201
rect 3142 50164 3148 50176
rect 3103 50136 3148 50164
rect 3142 50124 3148 50136
rect 3200 50124 3206 50176
rect 23290 50164 23296 50176
rect 23251 50136 23296 50164
rect 23290 50124 23296 50136
rect 23348 50124 23354 50176
rect 1104 50074 68816 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 14246 50074
rect 14298 50022 14310 50074
rect 14362 50022 14374 50074
rect 14426 50022 14438 50074
rect 14490 50022 24246 50074
rect 24298 50022 24310 50074
rect 24362 50022 24374 50074
rect 24426 50022 24438 50074
rect 24490 50022 34246 50074
rect 34298 50022 34310 50074
rect 34362 50022 34374 50074
rect 34426 50022 34438 50074
rect 34490 50022 44246 50074
rect 44298 50022 44310 50074
rect 44362 50022 44374 50074
rect 44426 50022 44438 50074
rect 44490 50022 54246 50074
rect 54298 50022 54310 50074
rect 54362 50022 54374 50074
rect 54426 50022 54438 50074
rect 54490 50022 64246 50074
rect 64298 50022 64310 50074
rect 64362 50022 64374 50074
rect 64426 50022 64438 50074
rect 64490 50022 68816 50074
rect 1104 50000 68816 50022
rect 23290 49920 23296 49972
rect 23348 49960 23354 49972
rect 65426 49960 65432 49972
rect 23348 49932 65432 49960
rect 23348 49920 23354 49932
rect 65426 49920 65432 49932
rect 65484 49920 65490 49972
rect 30926 49892 30932 49904
rect 20088 49864 30932 49892
rect 1762 49824 1768 49836
rect 1723 49796 1768 49824
rect 1762 49784 1768 49796
rect 1820 49784 1826 49836
rect 2593 49827 2651 49833
rect 2593 49824 2605 49827
rect 1964 49796 2605 49824
rect 1964 49765 1992 49796
rect 2593 49793 2605 49796
rect 2639 49824 2651 49827
rect 11790 49824 11796 49836
rect 2639 49796 11796 49824
rect 2639 49793 2651 49796
rect 2593 49787 2651 49793
rect 11790 49784 11796 49796
rect 11848 49784 11854 49836
rect 20088 49833 20116 49864
rect 30926 49852 30932 49864
rect 30984 49852 30990 49904
rect 34885 49895 34943 49901
rect 34885 49861 34897 49895
rect 34931 49892 34943 49895
rect 34974 49892 34980 49904
rect 34931 49864 34980 49892
rect 34931 49861 34943 49864
rect 34885 49855 34943 49861
rect 34974 49852 34980 49864
rect 35032 49852 35038 49904
rect 20073 49827 20131 49833
rect 20073 49793 20085 49827
rect 20119 49793 20131 49827
rect 21361 49827 21419 49833
rect 21361 49824 21373 49827
rect 20073 49787 20131 49793
rect 20824 49796 21373 49824
rect 1949 49759 2007 49765
rect 1949 49725 1961 49759
rect 1995 49725 2007 49759
rect 1949 49719 2007 49725
rect 6914 49716 6920 49768
rect 6972 49756 6978 49768
rect 20824 49765 20852 49796
rect 21361 49793 21373 49796
rect 21407 49824 21419 49827
rect 33870 49824 33876 49836
rect 21407 49796 33876 49824
rect 21407 49793 21419 49796
rect 21361 49787 21419 49793
rect 33870 49784 33876 49796
rect 33928 49784 33934 49836
rect 35437 49827 35495 49833
rect 35437 49824 35449 49827
rect 34348 49796 35449 49824
rect 34348 49765 34376 49796
rect 35437 49793 35449 49796
rect 35483 49824 35495 49827
rect 35483 49796 45554 49824
rect 35483 49793 35495 49796
rect 35437 49787 35495 49793
rect 20809 49759 20867 49765
rect 6972 49728 20760 49756
rect 6972 49716 6978 49728
rect 20732 49620 20760 49728
rect 20809 49725 20821 49759
rect 20855 49725 20867 49759
rect 34333 49759 34391 49765
rect 34333 49756 34345 49759
rect 20809 49719 20867 49725
rect 21008 49728 34345 49756
rect 21008 49620 21036 49728
rect 34333 49725 34345 49728
rect 34379 49725 34391 49759
rect 34517 49759 34575 49765
rect 34517 49756 34529 49759
rect 34333 49719 34391 49725
rect 34440 49728 34529 49756
rect 33962 49648 33968 49700
rect 34020 49688 34026 49700
rect 34440 49688 34468 49728
rect 34517 49725 34529 49728
rect 34563 49725 34575 49759
rect 34517 49719 34575 49725
rect 34698 49716 34704 49768
rect 34756 49765 34762 49768
rect 34756 49756 34764 49765
rect 35989 49759 36047 49765
rect 35989 49756 36001 49759
rect 34756 49728 36001 49756
rect 34756 49719 34764 49728
rect 35989 49725 36001 49728
rect 36035 49725 36047 49759
rect 45526 49756 45554 49796
rect 62758 49756 62764 49768
rect 45526 49728 62764 49756
rect 35989 49719 36047 49725
rect 34756 49716 34762 49719
rect 62758 49716 62764 49728
rect 62816 49716 62822 49768
rect 34020 49660 34468 49688
rect 34609 49691 34667 49697
rect 34020 49648 34026 49660
rect 34609 49657 34621 49691
rect 34655 49688 34667 49691
rect 40126 49688 40132 49700
rect 34655 49660 40132 49688
rect 34655 49657 34667 49660
rect 34609 49651 34667 49657
rect 20732 49592 21036 49620
rect 28258 49580 28264 49632
rect 28316 49620 28322 49632
rect 33781 49623 33839 49629
rect 33781 49620 33793 49623
rect 28316 49592 33793 49620
rect 28316 49580 28322 49592
rect 33781 49589 33793 49592
rect 33827 49620 33839 49623
rect 34624 49620 34652 49651
rect 40126 49648 40132 49660
rect 40184 49648 40190 49700
rect 33827 49592 34652 49620
rect 33827 49589 33839 49592
rect 33781 49583 33839 49589
rect 1104 49530 68816 49552
rect 1104 49478 9246 49530
rect 9298 49478 9310 49530
rect 9362 49478 9374 49530
rect 9426 49478 9438 49530
rect 9490 49478 19246 49530
rect 19298 49478 19310 49530
rect 19362 49478 19374 49530
rect 19426 49478 19438 49530
rect 19490 49478 29246 49530
rect 29298 49478 29310 49530
rect 29362 49478 29374 49530
rect 29426 49478 29438 49530
rect 29490 49478 39246 49530
rect 39298 49478 39310 49530
rect 39362 49478 39374 49530
rect 39426 49478 39438 49530
rect 39490 49478 49246 49530
rect 49298 49478 49310 49530
rect 49362 49478 49374 49530
rect 49426 49478 49438 49530
rect 49490 49478 59246 49530
rect 59298 49478 59310 49530
rect 59362 49478 59374 49530
rect 59426 49478 59438 49530
rect 59490 49478 68816 49530
rect 1104 49456 68816 49478
rect 33962 49076 33968 49088
rect 33923 49048 33968 49076
rect 33962 49036 33968 49048
rect 34020 49036 34026 49088
rect 40126 49036 40132 49088
rect 40184 49076 40190 49088
rect 65794 49076 65800 49088
rect 40184 49048 65800 49076
rect 40184 49036 40190 49048
rect 65794 49036 65800 49048
rect 65852 49036 65858 49088
rect 1104 48986 68816 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 14246 48986
rect 14298 48934 14310 48986
rect 14362 48934 14374 48986
rect 14426 48934 14438 48986
rect 14490 48934 24246 48986
rect 24298 48934 24310 48986
rect 24362 48934 24374 48986
rect 24426 48934 24438 48986
rect 24490 48934 34246 48986
rect 34298 48934 34310 48986
rect 34362 48934 34374 48986
rect 34426 48934 34438 48986
rect 34490 48934 44246 48986
rect 44298 48934 44310 48986
rect 44362 48934 44374 48986
rect 44426 48934 44438 48986
rect 44490 48934 54246 48986
rect 54298 48934 54310 48986
rect 54362 48934 54374 48986
rect 54426 48934 54438 48986
rect 54490 48934 64246 48986
rect 64298 48934 64310 48986
rect 64362 48934 64374 48986
rect 64426 48934 64438 48986
rect 64490 48934 68816 48986
rect 1104 48912 68816 48934
rect 1104 48442 68816 48464
rect 1104 48390 9246 48442
rect 9298 48390 9310 48442
rect 9362 48390 9374 48442
rect 9426 48390 9438 48442
rect 9490 48390 19246 48442
rect 19298 48390 19310 48442
rect 19362 48390 19374 48442
rect 19426 48390 19438 48442
rect 19490 48390 29246 48442
rect 29298 48390 29310 48442
rect 29362 48390 29374 48442
rect 29426 48390 29438 48442
rect 29490 48390 39246 48442
rect 39298 48390 39310 48442
rect 39362 48390 39374 48442
rect 39426 48390 39438 48442
rect 39490 48390 49246 48442
rect 49298 48390 49310 48442
rect 49362 48390 49374 48442
rect 49426 48390 49438 48442
rect 49490 48390 59246 48442
rect 59298 48390 59310 48442
rect 59362 48390 59374 48442
rect 59426 48390 59438 48442
rect 59490 48390 68816 48442
rect 1104 48368 68816 48390
rect 26326 48152 26332 48204
rect 26384 48192 26390 48204
rect 27522 48192 27528 48204
rect 26384 48164 27528 48192
rect 26384 48152 26390 48164
rect 27522 48152 27528 48164
rect 27580 48152 27586 48204
rect 66806 48152 66812 48204
rect 66864 48192 66870 48204
rect 67913 48195 67971 48201
rect 67913 48192 67925 48195
rect 66864 48164 67925 48192
rect 66864 48152 66870 48164
rect 67913 48161 67925 48164
rect 67959 48161 67971 48195
rect 67913 48155 67971 48161
rect 68094 48056 68100 48068
rect 68055 48028 68100 48056
rect 68094 48016 68100 48028
rect 68152 48016 68158 48068
rect 45002 47988 45008 48000
rect 44963 47960 45008 47988
rect 45002 47948 45008 47960
rect 45060 47948 45066 48000
rect 1104 47898 68816 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 14246 47898
rect 14298 47846 14310 47898
rect 14362 47846 14374 47898
rect 14426 47846 14438 47898
rect 14490 47846 24246 47898
rect 24298 47846 24310 47898
rect 24362 47846 24374 47898
rect 24426 47846 24438 47898
rect 24490 47846 34246 47898
rect 34298 47846 34310 47898
rect 34362 47846 34374 47898
rect 34426 47846 34438 47898
rect 34490 47846 44246 47898
rect 44298 47846 44310 47898
rect 44362 47846 44374 47898
rect 44426 47846 44438 47898
rect 44490 47846 54246 47898
rect 54298 47846 54310 47898
rect 54362 47846 54374 47898
rect 54426 47846 54438 47898
rect 54490 47846 64246 47898
rect 64298 47846 64310 47898
rect 64362 47846 64374 47898
rect 64426 47846 64438 47898
rect 64490 47846 68816 47898
rect 1104 47824 68816 47846
rect 33226 47608 33232 47660
rect 33284 47648 33290 47660
rect 40402 47648 40408 47660
rect 33284 47620 40408 47648
rect 33284 47608 33290 47620
rect 40402 47608 40408 47620
rect 40460 47608 40466 47660
rect 40310 47540 40316 47592
rect 40368 47580 40374 47592
rect 65334 47580 65340 47592
rect 40368 47552 65340 47580
rect 40368 47540 40374 47552
rect 65334 47540 65340 47552
rect 65392 47540 65398 47592
rect 1104 47354 68816 47376
rect 1104 47302 9246 47354
rect 9298 47302 9310 47354
rect 9362 47302 9374 47354
rect 9426 47302 9438 47354
rect 9490 47302 19246 47354
rect 19298 47302 19310 47354
rect 19362 47302 19374 47354
rect 19426 47302 19438 47354
rect 19490 47302 29246 47354
rect 29298 47302 29310 47354
rect 29362 47302 29374 47354
rect 29426 47302 29438 47354
rect 29490 47302 39246 47354
rect 39298 47302 39310 47354
rect 39362 47302 39374 47354
rect 39426 47302 39438 47354
rect 39490 47302 49246 47354
rect 49298 47302 49310 47354
rect 49362 47302 49374 47354
rect 49426 47302 49438 47354
rect 49490 47302 59246 47354
rect 59298 47302 59310 47354
rect 59362 47302 59374 47354
rect 59426 47302 59438 47354
rect 59490 47302 68816 47354
rect 1104 47280 68816 47302
rect 27522 47200 27528 47252
rect 27580 47240 27586 47252
rect 31757 47243 31815 47249
rect 31757 47240 31769 47243
rect 27580 47212 31769 47240
rect 27580 47200 27586 47212
rect 31757 47209 31769 47212
rect 31803 47209 31815 47243
rect 31757 47203 31815 47209
rect 1854 47172 1860 47184
rect 1815 47144 1860 47172
rect 1854 47132 1860 47144
rect 1912 47132 1918 47184
rect 31662 47172 31668 47184
rect 25424 47144 31668 47172
rect 25424 47113 25452 47144
rect 31662 47132 31668 47144
rect 31720 47132 31726 47184
rect 25409 47107 25467 47113
rect 25409 47073 25421 47107
rect 25455 47073 25467 47107
rect 31772 47104 31800 47203
rect 31846 47132 31852 47184
rect 31904 47172 31910 47184
rect 40770 47172 40776 47184
rect 31904 47144 40776 47172
rect 31904 47132 31910 47144
rect 40770 47132 40776 47144
rect 40828 47132 40834 47184
rect 32401 47107 32459 47113
rect 32401 47104 32413 47107
rect 31772 47076 32413 47104
rect 25409 47067 25467 47073
rect 32401 47073 32413 47076
rect 32447 47073 32459 47107
rect 67913 47107 67971 47113
rect 67913 47104 67925 47107
rect 32401 47067 32459 47073
rect 67284 47076 67925 47104
rect 26053 47039 26111 47045
rect 26053 47005 26065 47039
rect 26099 47036 26111 47039
rect 44818 47036 44824 47048
rect 26099 47008 44824 47036
rect 26099 47005 26111 47008
rect 26053 46999 26111 47005
rect 44818 46996 44824 47008
rect 44876 46996 44882 47048
rect 2041 46971 2099 46977
rect 2041 46937 2053 46971
rect 2087 46968 2099 46971
rect 32582 46968 32588 46980
rect 2087 46940 32444 46968
rect 32543 46940 32588 46968
rect 2087 46937 2099 46940
rect 2041 46931 2099 46937
rect 32416 46900 32444 46940
rect 32582 46928 32588 46940
rect 32640 46928 32646 46980
rect 33962 46968 33968 46980
rect 32692 46940 33968 46968
rect 32692 46900 32720 46940
rect 33962 46928 33968 46940
rect 34020 46928 34026 46980
rect 39669 46971 39727 46977
rect 39669 46937 39681 46971
rect 39715 46968 39727 46971
rect 46750 46968 46756 46980
rect 39715 46940 46756 46968
rect 39715 46937 39727 46940
rect 39669 46931 39727 46937
rect 46750 46928 46756 46940
rect 46808 46928 46814 46980
rect 48682 46928 48688 46980
rect 48740 46968 48746 46980
rect 49605 46971 49663 46977
rect 49605 46968 49617 46971
rect 48740 46940 49617 46968
rect 48740 46928 48746 46940
rect 49605 46937 49617 46940
rect 49651 46937 49663 46971
rect 49605 46931 49663 46937
rect 67174 46928 67180 46980
rect 67232 46968 67238 46980
rect 67284 46977 67312 47076
rect 67913 47073 67925 47076
rect 67959 47073 67971 47107
rect 67913 47067 67971 47073
rect 67269 46971 67327 46977
rect 67269 46968 67281 46971
rect 67232 46940 67281 46968
rect 67232 46928 67238 46940
rect 67269 46937 67281 46940
rect 67315 46937 67327 46971
rect 68094 46968 68100 46980
rect 68055 46940 68100 46968
rect 67269 46931 67327 46937
rect 68094 46928 68100 46940
rect 68152 46928 68158 46980
rect 32416 46872 32720 46900
rect 1104 46810 68816 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 14246 46810
rect 14298 46758 14310 46810
rect 14362 46758 14374 46810
rect 14426 46758 14438 46810
rect 14490 46758 24246 46810
rect 24298 46758 24310 46810
rect 24362 46758 24374 46810
rect 24426 46758 24438 46810
rect 24490 46758 34246 46810
rect 34298 46758 34310 46810
rect 34362 46758 34374 46810
rect 34426 46758 34438 46810
rect 34490 46758 44246 46810
rect 44298 46758 44310 46810
rect 44362 46758 44374 46810
rect 44426 46758 44438 46810
rect 44490 46758 54246 46810
rect 54298 46758 54310 46810
rect 54362 46758 54374 46810
rect 54426 46758 54438 46810
rect 54490 46758 64246 46810
rect 64298 46758 64310 46810
rect 64362 46758 64374 46810
rect 64426 46758 64438 46810
rect 64490 46758 68816 46810
rect 1104 46736 68816 46758
rect 1673 46699 1731 46705
rect 1673 46665 1685 46699
rect 1719 46696 1731 46699
rect 1854 46696 1860 46708
rect 1719 46668 1860 46696
rect 1719 46665 1731 46668
rect 1673 46659 1731 46665
rect 1854 46656 1860 46668
rect 1912 46656 1918 46708
rect 7561 46563 7619 46569
rect 7561 46529 7573 46563
rect 7607 46560 7619 46563
rect 7607 46532 26234 46560
rect 7607 46529 7619 46532
rect 7561 46523 7619 46529
rect 21269 46495 21327 46501
rect 21269 46461 21281 46495
rect 21315 46461 21327 46495
rect 26206 46492 26234 46532
rect 60734 46492 60740 46504
rect 26206 46464 60740 46492
rect 21269 46455 21327 46461
rect 21284 46424 21312 46455
rect 60734 46452 60740 46464
rect 60792 46452 60798 46504
rect 63678 46424 63684 46436
rect 21284 46396 63684 46424
rect 63678 46384 63684 46396
rect 63736 46384 63742 46436
rect 1104 46266 68816 46288
rect 1104 46214 9246 46266
rect 9298 46214 9310 46266
rect 9362 46214 9374 46266
rect 9426 46214 9438 46266
rect 9490 46214 19246 46266
rect 19298 46214 19310 46266
rect 19362 46214 19374 46266
rect 19426 46214 19438 46266
rect 19490 46214 29246 46266
rect 29298 46214 29310 46266
rect 29362 46214 29374 46266
rect 29426 46214 29438 46266
rect 29490 46214 39246 46266
rect 39298 46214 39310 46266
rect 39362 46214 39374 46266
rect 39426 46214 39438 46266
rect 39490 46214 49246 46266
rect 49298 46214 49310 46266
rect 49362 46214 49374 46266
rect 49426 46214 49438 46266
rect 49490 46214 59246 46266
rect 59298 46214 59310 46266
rect 59362 46214 59374 46266
rect 59426 46214 59438 46266
rect 59490 46214 68816 46266
rect 1104 46192 68816 46214
rect 2406 46112 2412 46164
rect 2464 46152 2470 46164
rect 2501 46155 2559 46161
rect 2501 46152 2513 46155
rect 2464 46124 2513 46152
rect 2464 46112 2470 46124
rect 2501 46121 2513 46124
rect 2547 46121 2559 46155
rect 2501 46115 2559 46121
rect 1949 46087 2007 46093
rect 1949 46053 1961 46087
rect 1995 46084 2007 46087
rect 2424 46084 2452 46112
rect 1995 46056 2452 46084
rect 1995 46053 2007 46056
rect 1949 46047 2007 46053
rect 1762 45948 1768 45960
rect 1723 45920 1768 45948
rect 1762 45908 1768 45920
rect 1820 45908 1826 45960
rect 39114 45772 39120 45824
rect 39172 45812 39178 45824
rect 39301 45815 39359 45821
rect 39301 45812 39313 45815
rect 39172 45784 39313 45812
rect 39172 45772 39178 45784
rect 39301 45781 39313 45784
rect 39347 45781 39359 45815
rect 39301 45775 39359 45781
rect 1104 45722 68816 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 14246 45722
rect 14298 45670 14310 45722
rect 14362 45670 14374 45722
rect 14426 45670 14438 45722
rect 14490 45670 24246 45722
rect 24298 45670 24310 45722
rect 24362 45670 24374 45722
rect 24426 45670 24438 45722
rect 24490 45670 34246 45722
rect 34298 45670 34310 45722
rect 34362 45670 34374 45722
rect 34426 45670 34438 45722
rect 34490 45670 44246 45722
rect 44298 45670 44310 45722
rect 44362 45670 44374 45722
rect 44426 45670 44438 45722
rect 44490 45670 54246 45722
rect 54298 45670 54310 45722
rect 54362 45670 54374 45722
rect 54426 45670 54438 45722
rect 54490 45670 64246 45722
rect 64298 45670 64310 45722
rect 64362 45670 64374 45722
rect 64426 45670 64438 45722
rect 64490 45670 68816 45722
rect 1104 45648 68816 45670
rect 39942 45540 39948 45552
rect 39903 45512 39948 45540
rect 39942 45500 39948 45512
rect 40000 45500 40006 45552
rect 58069 45543 58127 45549
rect 58069 45509 58081 45543
rect 58115 45540 58127 45543
rect 58618 45540 58624 45552
rect 58115 45512 58624 45540
rect 58115 45509 58127 45512
rect 58069 45503 58127 45509
rect 58618 45500 58624 45512
rect 58676 45500 58682 45552
rect 65610 45472 65616 45484
rect 40972 45444 65616 45472
rect 12986 45404 12992 45416
rect 12947 45376 12992 45404
rect 12986 45364 12992 45376
rect 13044 45364 13050 45416
rect 40126 45413 40132 45416
rect 39393 45407 39451 45413
rect 39393 45373 39405 45407
rect 39439 45404 39451 45407
rect 40077 45407 40132 45413
rect 40077 45404 40089 45407
rect 39439 45376 40089 45404
rect 39439 45373 39451 45376
rect 39393 45367 39451 45373
rect 40077 45373 40089 45376
rect 40123 45373 40132 45407
rect 40077 45367 40132 45373
rect 40126 45364 40132 45367
rect 40184 45404 40190 45416
rect 40310 45404 40316 45416
rect 40184 45376 40225 45404
rect 40271 45376 40316 45404
rect 40184 45364 40190 45376
rect 40310 45364 40316 45376
rect 40368 45364 40374 45416
rect 40497 45407 40555 45413
rect 40497 45373 40509 45407
rect 40543 45373 40555 45407
rect 40497 45367 40555 45373
rect 39114 45296 39120 45348
rect 39172 45336 39178 45348
rect 40221 45339 40279 45345
rect 40221 45336 40233 45339
rect 39172 45308 40233 45336
rect 39172 45296 39178 45308
rect 40221 45305 40233 45308
rect 40267 45305 40279 45339
rect 40221 45299 40279 45305
rect 39850 45228 39856 45280
rect 39908 45268 39914 45280
rect 40512 45268 40540 45367
rect 40972 45277 41000 45444
rect 65610 45432 65616 45444
rect 65668 45432 65674 45484
rect 67453 45407 67511 45413
rect 67453 45373 67465 45407
rect 67499 45404 67511 45407
rect 68094 45404 68100 45416
rect 67499 45376 68100 45404
rect 67499 45373 67511 45376
rect 67453 45367 67511 45373
rect 68094 45364 68100 45376
rect 68152 45364 68158 45416
rect 40957 45271 41015 45277
rect 40957 45268 40969 45271
rect 39908 45240 40969 45268
rect 39908 45228 39914 45240
rect 40957 45237 40969 45240
rect 41003 45237 41015 45271
rect 40957 45231 41015 45237
rect 1104 45178 68816 45200
rect 1104 45126 9246 45178
rect 9298 45126 9310 45178
rect 9362 45126 9374 45178
rect 9426 45126 9438 45178
rect 9490 45126 19246 45178
rect 19298 45126 19310 45178
rect 19362 45126 19374 45178
rect 19426 45126 19438 45178
rect 19490 45126 29246 45178
rect 29298 45126 29310 45178
rect 29362 45126 29374 45178
rect 29426 45126 29438 45178
rect 29490 45126 39246 45178
rect 39298 45126 39310 45178
rect 39362 45126 39374 45178
rect 39426 45126 39438 45178
rect 39490 45126 49246 45178
rect 49298 45126 49310 45178
rect 49362 45126 49374 45178
rect 49426 45126 49438 45178
rect 49490 45126 59246 45178
rect 59298 45126 59310 45178
rect 59362 45126 59374 45178
rect 59426 45126 59438 45178
rect 59490 45126 68816 45178
rect 1104 45104 68816 45126
rect 12986 45024 12992 45076
rect 13044 45064 13050 45076
rect 66530 45064 66536 45076
rect 13044 45036 66536 45064
rect 13044 45024 13050 45036
rect 66530 45024 66536 45036
rect 66588 45024 66594 45076
rect 1949 44999 2007 45005
rect 1949 44965 1961 44999
rect 1995 44996 2007 44999
rect 2130 44996 2136 45008
rect 1995 44968 2136 44996
rect 1995 44965 2007 44968
rect 1949 44959 2007 44965
rect 2130 44956 2136 44968
rect 2188 44996 2194 45008
rect 2501 44999 2559 45005
rect 2501 44996 2513 44999
rect 2188 44968 2513 44996
rect 2188 44956 2194 44968
rect 2501 44965 2513 44968
rect 2547 44965 2559 44999
rect 2501 44959 2559 44965
rect 13630 44956 13636 45008
rect 13688 44996 13694 45008
rect 13688 44968 18276 44996
rect 13688 44956 13694 44968
rect 17046 44931 17104 44937
rect 17046 44928 17058 44931
rect 16040 44900 17058 44928
rect 7282 44752 7288 44804
rect 7340 44792 7346 44804
rect 15933 44795 15991 44801
rect 15933 44792 15945 44795
rect 7340 44764 15945 44792
rect 7340 44752 7346 44764
rect 15933 44761 15945 44764
rect 15979 44761 15991 44795
rect 15933 44755 15991 44761
rect 1854 44724 1860 44736
rect 1815 44696 1860 44724
rect 1854 44684 1860 44696
rect 1912 44684 1918 44736
rect 7006 44684 7012 44736
rect 7064 44724 7070 44736
rect 15289 44727 15347 44733
rect 15289 44724 15301 44727
rect 7064 44696 15301 44724
rect 7064 44684 7070 44696
rect 15289 44693 15301 44696
rect 15335 44724 15347 44727
rect 16040 44724 16068 44900
rect 17046 44897 17058 44900
rect 17092 44897 17104 44931
rect 17046 44891 17104 44897
rect 17218 44888 17224 44940
rect 17276 44888 17282 44940
rect 17678 44888 17684 44940
rect 17736 44928 17742 44940
rect 17862 44928 17868 44940
rect 17736 44900 17868 44928
rect 17736 44888 17742 44900
rect 17862 44888 17868 44900
rect 17920 44888 17926 44940
rect 18248 44928 18276 44968
rect 21358 44956 21364 45008
rect 21416 44996 21422 45008
rect 30282 44996 30288 45008
rect 21416 44968 30288 44996
rect 21416 44956 21422 44968
rect 30282 44956 30288 44968
rect 30340 44956 30346 45008
rect 58710 44996 58716 45008
rect 58671 44968 58716 44996
rect 58710 44956 58716 44968
rect 58768 44996 58774 45008
rect 59541 44999 59599 45005
rect 59541 44996 59553 44999
rect 58768 44968 59553 44996
rect 58768 44956 58774 44968
rect 59541 44965 59553 44968
rect 59587 44965 59599 44999
rect 59541 44959 59599 44965
rect 34146 44928 34152 44940
rect 18248 44900 34152 44928
rect 34146 44888 34152 44900
rect 34204 44888 34210 44940
rect 58529 44931 58587 44937
rect 58529 44897 58541 44931
rect 58575 44928 58587 44931
rect 58618 44928 58624 44940
rect 58575 44900 58624 44928
rect 58575 44897 58587 44900
rect 58529 44891 58587 44897
rect 58618 44888 58624 44900
rect 58676 44888 58682 44940
rect 58802 44928 58808 44940
rect 58763 44900 58808 44928
rect 58802 44888 58808 44900
rect 58860 44888 58866 44940
rect 58897 44931 58955 44937
rect 58897 44897 58909 44931
rect 58943 44897 58955 44931
rect 58897 44891 58955 44897
rect 17236 44860 17264 44888
rect 17313 44863 17371 44869
rect 17313 44860 17325 44863
rect 17236 44832 17325 44860
rect 17313 44829 17325 44832
rect 17359 44860 17371 44863
rect 17359 44832 17908 44860
rect 17359 44829 17371 44832
rect 17313 44823 17371 44829
rect 17880 44736 17908 44832
rect 17862 44724 17868 44736
rect 15335 44696 16068 44724
rect 17823 44696 17868 44724
rect 15335 44693 15347 44696
rect 15289 44687 15347 44693
rect 17862 44684 17868 44696
rect 17920 44684 17926 44736
rect 39577 44727 39635 44733
rect 39577 44693 39589 44727
rect 39623 44724 39635 44727
rect 40310 44724 40316 44736
rect 39623 44696 40316 44724
rect 39623 44693 39635 44696
rect 39577 44687 39635 44693
rect 40310 44684 40316 44696
rect 40368 44684 40374 44736
rect 49602 44684 49608 44736
rect 49660 44724 49666 44736
rect 58069 44727 58127 44733
rect 58069 44724 58081 44727
rect 49660 44696 58081 44724
rect 49660 44684 49666 44696
rect 58069 44693 58081 44696
rect 58115 44724 58127 44727
rect 58912 44724 58940 44891
rect 59081 44795 59139 44801
rect 59081 44761 59093 44795
rect 59127 44792 59139 44795
rect 59998 44792 60004 44804
rect 59127 44764 60004 44792
rect 59127 44761 59139 44764
rect 59081 44755 59139 44761
rect 59998 44752 60004 44764
rect 60056 44752 60062 44804
rect 58115 44696 58940 44724
rect 58115 44693 58127 44696
rect 58069 44687 58127 44693
rect 1104 44634 68816 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 14246 44634
rect 14298 44582 14310 44634
rect 14362 44582 14374 44634
rect 14426 44582 14438 44634
rect 14490 44582 24246 44634
rect 24298 44582 24310 44634
rect 24362 44582 24374 44634
rect 24426 44582 24438 44634
rect 24490 44582 34246 44634
rect 34298 44582 34310 44634
rect 34362 44582 34374 44634
rect 34426 44582 34438 44634
rect 34490 44582 44246 44634
rect 44298 44582 44310 44634
rect 44362 44582 44374 44634
rect 44426 44582 44438 44634
rect 44490 44582 54246 44634
rect 54298 44582 54310 44634
rect 54362 44582 54374 44634
rect 54426 44582 54438 44634
rect 54490 44582 64246 44634
rect 64298 44582 64310 44634
rect 64362 44582 64374 44634
rect 64426 44582 64438 44634
rect 64490 44582 68816 44634
rect 1104 44560 68816 44582
rect 58069 44523 58127 44529
rect 58069 44489 58081 44523
rect 58115 44520 58127 44523
rect 58253 44523 58311 44529
rect 58253 44520 58265 44523
rect 58115 44492 58265 44520
rect 58115 44489 58127 44492
rect 58069 44483 58127 44489
rect 58253 44489 58265 44492
rect 58299 44520 58311 44523
rect 58802 44520 58808 44532
rect 58299 44492 58808 44520
rect 58299 44489 58311 44492
rect 58253 44483 58311 44489
rect 58802 44480 58808 44492
rect 58860 44480 58866 44532
rect 11698 44344 11704 44396
rect 11756 44384 11762 44396
rect 21358 44384 21364 44396
rect 11756 44356 21364 44384
rect 11756 44344 11762 44356
rect 21358 44344 21364 44356
rect 21416 44344 21422 44396
rect 10686 44316 10692 44328
rect 10647 44288 10692 44316
rect 10686 44276 10692 44288
rect 10744 44276 10750 44328
rect 48958 44208 48964 44260
rect 49016 44248 49022 44260
rect 49602 44248 49608 44260
rect 49016 44220 49608 44248
rect 49016 44208 49022 44220
rect 49602 44208 49608 44220
rect 49660 44208 49666 44260
rect 33134 44140 33140 44192
rect 33192 44180 33198 44192
rect 58069 44183 58127 44189
rect 58069 44180 58081 44183
rect 33192 44152 58081 44180
rect 33192 44140 33198 44152
rect 58069 44149 58081 44152
rect 58115 44149 58127 44183
rect 58069 44143 58127 44149
rect 1104 44090 68816 44112
rect 1104 44038 9246 44090
rect 9298 44038 9310 44090
rect 9362 44038 9374 44090
rect 9426 44038 9438 44090
rect 9490 44038 19246 44090
rect 19298 44038 19310 44090
rect 19362 44038 19374 44090
rect 19426 44038 19438 44090
rect 19490 44038 29246 44090
rect 29298 44038 29310 44090
rect 29362 44038 29374 44090
rect 29426 44038 29438 44090
rect 29490 44038 39246 44090
rect 39298 44038 39310 44090
rect 39362 44038 39374 44090
rect 39426 44038 39438 44090
rect 39490 44038 49246 44090
rect 49298 44038 49310 44090
rect 49362 44038 49374 44090
rect 49426 44038 49438 44090
rect 49490 44038 59246 44090
rect 59298 44038 59310 44090
rect 59362 44038 59374 44090
rect 59426 44038 59438 44090
rect 59490 44038 68816 44090
rect 1104 44016 68816 44038
rect 55306 43936 55312 43988
rect 55364 43976 55370 43988
rect 56042 43976 56048 43988
rect 55364 43948 56048 43976
rect 55364 43936 55370 43948
rect 56042 43936 56048 43948
rect 56100 43936 56106 43988
rect 30469 43843 30527 43849
rect 30469 43809 30481 43843
rect 30515 43840 30527 43843
rect 30558 43840 30564 43852
rect 30515 43812 30564 43840
rect 30515 43809 30527 43812
rect 30469 43803 30527 43809
rect 30558 43800 30564 43812
rect 30616 43840 30622 43852
rect 31113 43843 31171 43849
rect 31113 43840 31125 43843
rect 30616 43812 31125 43840
rect 30616 43800 30622 43812
rect 31113 43809 31125 43812
rect 31159 43809 31171 43843
rect 62390 43840 62396 43852
rect 62351 43812 62396 43840
rect 31113 43803 31171 43809
rect 62390 43800 62396 43812
rect 62448 43840 62454 43852
rect 62853 43843 62911 43849
rect 62853 43840 62865 43843
rect 62448 43812 62865 43840
rect 62448 43800 62454 43812
rect 62853 43809 62865 43812
rect 62899 43809 62911 43843
rect 62853 43803 62911 43809
rect 56042 43732 56048 43784
rect 56100 43772 56106 43784
rect 62117 43775 62175 43781
rect 62117 43772 62129 43775
rect 56100 43744 62129 43772
rect 56100 43732 56106 43744
rect 62117 43741 62129 43744
rect 62163 43741 62175 43775
rect 62117 43735 62175 43741
rect 17862 43596 17868 43648
rect 17920 43636 17926 43648
rect 30653 43639 30711 43645
rect 30653 43636 30665 43639
rect 17920 43608 30665 43636
rect 17920 43596 17926 43608
rect 30653 43605 30665 43608
rect 30699 43636 30711 43639
rect 30742 43636 30748 43648
rect 30699 43608 30748 43636
rect 30699 43605 30711 43608
rect 30653 43599 30711 43605
rect 30742 43596 30748 43608
rect 30800 43596 30806 43648
rect 35710 43636 35716 43648
rect 35671 43608 35716 43636
rect 35710 43596 35716 43608
rect 35768 43596 35774 43648
rect 65429 43639 65487 43645
rect 65429 43605 65441 43639
rect 65475 43636 65487 43639
rect 67542 43636 67548 43648
rect 65475 43608 67548 43636
rect 65475 43605 65487 43608
rect 65429 43599 65487 43605
rect 67542 43596 67548 43608
rect 67600 43596 67606 43648
rect 1104 43546 68816 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 14246 43546
rect 14298 43494 14310 43546
rect 14362 43494 14374 43546
rect 14426 43494 14438 43546
rect 14490 43494 24246 43546
rect 24298 43494 24310 43546
rect 24362 43494 24374 43546
rect 24426 43494 24438 43546
rect 24490 43494 34246 43546
rect 34298 43494 34310 43546
rect 34362 43494 34374 43546
rect 34426 43494 34438 43546
rect 34490 43494 44246 43546
rect 44298 43494 44310 43546
rect 44362 43494 44374 43546
rect 44426 43494 44438 43546
rect 44490 43494 54246 43546
rect 54298 43494 54310 43546
rect 54362 43494 54374 43546
rect 54426 43494 54438 43546
rect 54490 43494 64246 43546
rect 64298 43494 64310 43546
rect 64362 43494 64374 43546
rect 64426 43494 64438 43546
rect 64490 43494 68816 43546
rect 1104 43472 68816 43494
rect 2961 43299 3019 43305
rect 2961 43265 2973 43299
rect 3007 43296 3019 43299
rect 3694 43296 3700 43308
rect 3007 43268 3700 43296
rect 3007 43265 3019 43268
rect 2961 43259 3019 43265
rect 3694 43256 3700 43268
rect 3752 43256 3758 43308
rect 17862 43296 17868 43308
rect 6886 43268 17868 43296
rect 3237 43231 3295 43237
rect 3237 43197 3249 43231
rect 3283 43228 3295 43231
rect 4341 43231 4399 43237
rect 4341 43228 4353 43231
rect 3283 43200 4353 43228
rect 3283 43197 3295 43200
rect 3237 43191 3295 43197
rect 4341 43197 4353 43200
rect 4387 43228 4399 43231
rect 6886 43228 6914 43268
rect 17862 43256 17868 43268
rect 17920 43256 17926 43308
rect 12986 43228 12992 43240
rect 4387 43200 6914 43228
rect 12947 43200 12992 43228
rect 4387 43197 4399 43200
rect 4341 43191 4399 43197
rect 12986 43188 12992 43200
rect 13044 43228 13050 43240
rect 13633 43231 13691 43237
rect 13633 43228 13645 43231
rect 13044 43200 13645 43228
rect 13044 43188 13050 43200
rect 13633 43197 13645 43200
rect 13679 43197 13691 43231
rect 13633 43191 13691 43197
rect 50065 43231 50123 43237
rect 50065 43197 50077 43231
rect 50111 43228 50123 43231
rect 60826 43228 60832 43240
rect 50111 43200 60832 43228
rect 50111 43197 50123 43200
rect 50065 43191 50123 43197
rect 60826 43188 60832 43200
rect 60884 43188 60890 43240
rect 3528 43132 4292 43160
rect 1857 43095 1915 43101
rect 1857 43061 1869 43095
rect 1903 43092 1915 43095
rect 3528 43092 3556 43132
rect 3694 43092 3700 43104
rect 1903 43064 3556 43092
rect 3655 43064 3700 43092
rect 1903 43061 1915 43064
rect 1857 43055 1915 43061
rect 3694 43052 3700 43064
rect 3752 43052 3758 43104
rect 4264 43092 4292 43132
rect 6886 43132 16574 43160
rect 6886 43092 6914 43132
rect 4264 43064 6914 43092
rect 13081 43095 13139 43101
rect 13081 43061 13093 43095
rect 13127 43092 13139 43095
rect 13354 43092 13360 43104
rect 13127 43064 13360 43092
rect 13127 43061 13139 43064
rect 13081 43055 13139 43061
rect 13354 43052 13360 43064
rect 13412 43052 13418 43104
rect 16546 43092 16574 43132
rect 33134 43092 33140 43104
rect 16546 43064 33140 43092
rect 33134 43052 33140 43064
rect 33192 43052 33198 43104
rect 1104 43002 68816 43024
rect 1104 42950 9246 43002
rect 9298 42950 9310 43002
rect 9362 42950 9374 43002
rect 9426 42950 9438 43002
rect 9490 42950 19246 43002
rect 19298 42950 19310 43002
rect 19362 42950 19374 43002
rect 19426 42950 19438 43002
rect 19490 42950 29246 43002
rect 29298 42950 29310 43002
rect 29362 42950 29374 43002
rect 29426 42950 29438 43002
rect 29490 42950 39246 43002
rect 39298 42950 39310 43002
rect 39362 42950 39374 43002
rect 39426 42950 39438 43002
rect 39490 42950 49246 43002
rect 49298 42950 49310 43002
rect 49362 42950 49374 43002
rect 49426 42950 49438 43002
rect 49490 42950 59246 43002
rect 59298 42950 59310 43002
rect 59362 42950 59374 43002
rect 59426 42950 59438 43002
rect 59490 42950 68816 43002
rect 1104 42928 68816 42950
rect 13354 42848 13360 42900
rect 13412 42888 13418 42900
rect 27246 42888 27252 42900
rect 13412 42860 27252 42888
rect 13412 42848 13418 42860
rect 27246 42848 27252 42860
rect 27304 42848 27310 42900
rect 49421 42755 49479 42761
rect 49421 42721 49433 42755
rect 49467 42721 49479 42755
rect 49421 42715 49479 42721
rect 48869 42687 48927 42693
rect 48869 42684 48881 42687
rect 45526 42656 48881 42684
rect 37182 42576 37188 42628
rect 37240 42616 37246 42628
rect 45526 42616 45554 42656
rect 48869 42653 48881 42656
rect 48915 42684 48927 42687
rect 49436 42684 49464 42715
rect 66714 42712 66720 42764
rect 66772 42752 66778 42764
rect 67913 42755 67971 42761
rect 67913 42752 67925 42755
rect 66772 42724 67925 42752
rect 66772 42712 66778 42724
rect 67913 42721 67925 42724
rect 67959 42721 67971 42755
rect 68094 42752 68100 42764
rect 68055 42724 68100 42752
rect 67913 42715 67971 42721
rect 68094 42712 68100 42724
rect 68152 42712 68158 42764
rect 50246 42684 50252 42696
rect 48915 42656 49464 42684
rect 50207 42656 50252 42684
rect 48915 42653 48927 42656
rect 48869 42647 48927 42653
rect 50246 42644 50252 42656
rect 50304 42644 50310 42696
rect 60182 42616 60188 42628
rect 37240 42588 45554 42616
rect 48056 42588 60188 42616
rect 37240 42576 37246 42588
rect 7834 42508 7840 42560
rect 7892 42548 7898 42560
rect 11701 42551 11759 42557
rect 11701 42548 11713 42551
rect 7892 42520 11713 42548
rect 7892 42508 7898 42520
rect 11701 42517 11713 42520
rect 11747 42517 11759 42551
rect 12802 42548 12808 42560
rect 12763 42520 12808 42548
rect 11701 42511 11759 42517
rect 12802 42508 12808 42520
rect 12860 42508 12866 42560
rect 20165 42551 20223 42557
rect 20165 42517 20177 42551
rect 20211 42548 20223 42551
rect 48056 42548 48084 42588
rect 60182 42576 60188 42588
rect 60240 42576 60246 42628
rect 20211 42520 48084 42548
rect 20211 42517 20223 42520
rect 20165 42511 20223 42517
rect 1104 42458 68816 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 14246 42458
rect 14298 42406 14310 42458
rect 14362 42406 14374 42458
rect 14426 42406 14438 42458
rect 14490 42406 24246 42458
rect 24298 42406 24310 42458
rect 24362 42406 24374 42458
rect 24426 42406 24438 42458
rect 24490 42406 34246 42458
rect 34298 42406 34310 42458
rect 34362 42406 34374 42458
rect 34426 42406 34438 42458
rect 34490 42406 44246 42458
rect 44298 42406 44310 42458
rect 44362 42406 44374 42458
rect 44426 42406 44438 42458
rect 44490 42406 54246 42458
rect 54298 42406 54310 42458
rect 54362 42406 54374 42458
rect 54426 42406 54438 42458
rect 54490 42406 64246 42458
rect 64298 42406 64310 42458
rect 64362 42406 64374 42458
rect 64426 42406 64438 42458
rect 64490 42406 68816 42458
rect 1104 42384 68816 42406
rect 12802 42304 12808 42356
rect 12860 42344 12866 42356
rect 49970 42344 49976 42356
rect 12860 42316 49976 42344
rect 12860 42304 12866 42316
rect 49970 42304 49976 42316
rect 50028 42304 50034 42356
rect 18322 42236 18328 42288
rect 18380 42276 18386 42288
rect 18693 42279 18751 42285
rect 18693 42276 18705 42279
rect 18380 42248 18705 42276
rect 18380 42236 18386 42248
rect 18693 42245 18705 42248
rect 18739 42276 18751 42279
rect 22922 42276 22928 42288
rect 18739 42248 22928 42276
rect 18739 42245 18751 42248
rect 18693 42239 18751 42245
rect 22922 42236 22928 42248
rect 22980 42236 22986 42288
rect 45526 42180 60734 42208
rect 1578 42140 1584 42152
rect 1539 42112 1584 42140
rect 1578 42100 1584 42112
rect 1636 42140 1642 42152
rect 2041 42143 2099 42149
rect 2041 42140 2053 42143
rect 1636 42112 2053 42140
rect 1636 42100 1642 42112
rect 2041 42109 2053 42112
rect 2087 42109 2099 42143
rect 2041 42103 2099 42109
rect 26605 42143 26663 42149
rect 26605 42109 26617 42143
rect 26651 42140 26663 42143
rect 45526 42140 45554 42180
rect 51350 42140 51356 42152
rect 26651 42112 45554 42140
rect 51311 42112 51356 42140
rect 26651 42109 26663 42112
rect 26605 42103 26663 42109
rect 51350 42100 51356 42112
rect 51408 42100 51414 42152
rect 60706 42140 60734 42180
rect 65518 42140 65524 42152
rect 60706 42112 65524 42140
rect 65518 42100 65524 42112
rect 65576 42100 65582 42152
rect 22922 42032 22928 42084
rect 22980 42072 22986 42084
rect 39114 42072 39120 42084
rect 22980 42044 39120 42072
rect 22980 42032 22986 42044
rect 39114 42032 39120 42044
rect 39172 42032 39178 42084
rect 21358 41964 21364 42016
rect 21416 42004 21422 42016
rect 53466 42004 53472 42016
rect 21416 41976 53472 42004
rect 21416 41964 21422 41976
rect 53466 41964 53472 41976
rect 53524 41964 53530 42016
rect 1104 41914 68816 41936
rect 1104 41862 9246 41914
rect 9298 41862 9310 41914
rect 9362 41862 9374 41914
rect 9426 41862 9438 41914
rect 9490 41862 19246 41914
rect 19298 41862 19310 41914
rect 19362 41862 19374 41914
rect 19426 41862 19438 41914
rect 19490 41862 29246 41914
rect 29298 41862 29310 41914
rect 29362 41862 29374 41914
rect 29426 41862 29438 41914
rect 29490 41862 39246 41914
rect 39298 41862 39310 41914
rect 39362 41862 39374 41914
rect 39426 41862 39438 41914
rect 39490 41862 49246 41914
rect 49298 41862 49310 41914
rect 49362 41862 49374 41914
rect 49426 41862 49438 41914
rect 49490 41862 59246 41914
rect 59298 41862 59310 41914
rect 59362 41862 59374 41914
rect 59426 41862 59438 41914
rect 59490 41862 68816 41914
rect 1104 41840 68816 41862
rect 17673 41803 17731 41809
rect 17673 41769 17685 41803
rect 17719 41800 17731 41803
rect 37826 41800 37832 41812
rect 17719 41772 37832 41800
rect 17719 41769 17731 41772
rect 17673 41763 17731 41769
rect 37826 41760 37832 41772
rect 37884 41760 37890 41812
rect 66898 41760 66904 41812
rect 66956 41800 66962 41812
rect 67269 41803 67327 41809
rect 67269 41800 67281 41803
rect 66956 41772 67281 41800
rect 66956 41760 66962 41772
rect 67269 41769 67281 41772
rect 67315 41769 67327 41803
rect 67269 41763 67327 41769
rect 21358 41732 21364 41744
rect 16040 41704 21364 41732
rect 16040 41673 16068 41704
rect 21358 41692 21364 41704
rect 21416 41692 21422 41744
rect 30742 41732 30748 41744
rect 30703 41704 30748 41732
rect 30742 41692 30748 41704
rect 30800 41692 30806 41744
rect 31297 41735 31355 41741
rect 31297 41701 31309 41735
rect 31343 41732 31355 41735
rect 31386 41732 31392 41744
rect 31343 41704 31392 41732
rect 31343 41701 31355 41704
rect 31297 41695 31355 41701
rect 31386 41692 31392 41704
rect 31444 41692 31450 41744
rect 67284 41732 67312 41763
rect 67913 41735 67971 41741
rect 67913 41732 67925 41735
rect 67284 41704 67925 41732
rect 67913 41701 67925 41704
rect 67959 41701 67971 41735
rect 67913 41695 67971 41701
rect 16025 41667 16083 41673
rect 16025 41633 16037 41667
rect 16071 41633 16083 41667
rect 16025 41627 16083 41633
rect 17678 41624 17684 41676
rect 17736 41664 17742 41676
rect 17860 41667 17918 41673
rect 17860 41664 17872 41667
rect 17736 41636 17872 41664
rect 17736 41624 17742 41636
rect 17860 41633 17872 41636
rect 17906 41633 17918 41667
rect 17860 41627 17918 41633
rect 16669 41463 16727 41469
rect 16669 41429 16681 41463
rect 16715 41460 16727 41463
rect 16942 41460 16948 41472
rect 16715 41432 16948 41460
rect 16715 41429 16727 41432
rect 16669 41423 16727 41429
rect 16942 41420 16948 41432
rect 17000 41420 17006 41472
rect 17880 41460 17908 41627
rect 17954 41624 17960 41676
rect 18012 41664 18018 41676
rect 18138 41673 18144 41676
rect 18095 41667 18144 41673
rect 18012 41636 18057 41664
rect 18012 41624 18018 41636
rect 18095 41633 18107 41667
rect 18141 41633 18144 41667
rect 18095 41627 18144 41633
rect 18138 41624 18144 41627
rect 18196 41624 18202 41676
rect 18233 41667 18291 41673
rect 18233 41633 18245 41667
rect 18279 41664 18291 41667
rect 18598 41664 18604 41676
rect 18279 41636 18604 41664
rect 18279 41633 18291 41636
rect 18233 41627 18291 41633
rect 18598 41624 18604 41636
rect 18656 41624 18662 41676
rect 30760 41596 30788 41692
rect 32677 41667 32735 41673
rect 32677 41633 32689 41667
rect 32723 41664 32735 41667
rect 33505 41667 33563 41673
rect 33505 41664 33517 41667
rect 32723 41636 33517 41664
rect 32723 41633 32735 41636
rect 32677 41627 32735 41633
rect 33505 41633 33517 41636
rect 33551 41664 33563 41667
rect 52086 41664 52092 41676
rect 33551 41636 52092 41664
rect 33551 41633 33563 41636
rect 33505 41627 33563 41633
rect 52086 41624 52092 41636
rect 52144 41624 52150 41676
rect 32953 41599 33011 41605
rect 32953 41596 32965 41599
rect 30760 41568 32965 41596
rect 32953 41565 32965 41568
rect 32999 41596 33011 41599
rect 41598 41596 41604 41608
rect 32999 41568 41604 41596
rect 32999 41565 33011 41568
rect 32953 41559 33011 41565
rect 41598 41556 41604 41568
rect 41656 41556 41662 41608
rect 18785 41531 18843 41537
rect 18785 41497 18797 41531
rect 18831 41528 18843 41531
rect 28258 41528 28264 41540
rect 18831 41500 28264 41528
rect 18831 41497 18843 41500
rect 18785 41491 18843 41497
rect 18800 41460 18828 41491
rect 28258 41488 28264 41500
rect 28316 41528 28322 41540
rect 28442 41528 28448 41540
rect 28316 41500 28448 41528
rect 28316 41488 28322 41500
rect 28442 41488 28448 41500
rect 28500 41488 28506 41540
rect 35897 41531 35955 41537
rect 35897 41497 35909 41531
rect 35943 41528 35955 41531
rect 62298 41528 62304 41540
rect 35943 41500 62304 41528
rect 35943 41497 35955 41500
rect 35897 41491 35955 41497
rect 62298 41488 62304 41500
rect 62356 41488 62362 41540
rect 68094 41528 68100 41540
rect 68055 41500 68100 41528
rect 68094 41488 68100 41500
rect 68152 41488 68158 41540
rect 17880 41432 18828 41460
rect 36722 41420 36728 41472
rect 36780 41460 36786 41472
rect 37182 41460 37188 41472
rect 36780 41432 37188 41460
rect 36780 41420 36786 41432
rect 37182 41420 37188 41432
rect 37240 41420 37246 41472
rect 57698 41460 57704 41472
rect 57659 41432 57704 41460
rect 57698 41420 57704 41432
rect 57756 41420 57762 41472
rect 1104 41370 68816 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 14246 41370
rect 14298 41318 14310 41370
rect 14362 41318 14374 41370
rect 14426 41318 14438 41370
rect 14490 41318 24246 41370
rect 24298 41318 24310 41370
rect 24362 41318 24374 41370
rect 24426 41318 24438 41370
rect 24490 41318 34246 41370
rect 34298 41318 34310 41370
rect 34362 41318 34374 41370
rect 34426 41318 34438 41370
rect 34490 41318 44246 41370
rect 44298 41318 44310 41370
rect 44362 41318 44374 41370
rect 44426 41318 44438 41370
rect 44490 41318 54246 41370
rect 54298 41318 54310 41370
rect 54362 41318 54374 41370
rect 54426 41318 54438 41370
rect 54490 41318 64246 41370
rect 64298 41318 64310 41370
rect 64362 41318 64374 41370
rect 64426 41318 64438 41370
rect 64490 41318 68816 41370
rect 1104 41296 68816 41318
rect 13814 41012 13820 41064
rect 13872 41052 13878 41064
rect 43533 41055 43591 41061
rect 43533 41052 43545 41055
rect 13872 41024 43545 41052
rect 13872 41012 13878 41024
rect 43533 41021 43545 41024
rect 43579 41021 43591 41055
rect 47026 41052 47032 41064
rect 46987 41024 47032 41052
rect 43533 41015 43591 41021
rect 47026 41012 47032 41024
rect 47084 41012 47090 41064
rect 65334 41012 65340 41064
rect 65392 41052 65398 41064
rect 66165 41055 66223 41061
rect 66165 41052 66177 41055
rect 65392 41024 66177 41052
rect 65392 41012 65398 41024
rect 66165 41021 66177 41024
rect 66211 41021 66223 41055
rect 66165 41015 66223 41021
rect 17494 40916 17500 40928
rect 17455 40888 17500 40916
rect 17494 40876 17500 40888
rect 17552 40876 17558 40928
rect 18598 40916 18604 40928
rect 18511 40888 18604 40916
rect 18598 40876 18604 40888
rect 18656 40916 18662 40928
rect 39114 40916 39120 40928
rect 18656 40888 39120 40916
rect 18656 40876 18662 40888
rect 39114 40876 39120 40888
rect 39172 40876 39178 40928
rect 1104 40826 68816 40848
rect 1104 40774 9246 40826
rect 9298 40774 9310 40826
rect 9362 40774 9374 40826
rect 9426 40774 9438 40826
rect 9490 40774 19246 40826
rect 19298 40774 19310 40826
rect 19362 40774 19374 40826
rect 19426 40774 19438 40826
rect 19490 40774 29246 40826
rect 29298 40774 29310 40826
rect 29362 40774 29374 40826
rect 29426 40774 29438 40826
rect 29490 40774 39246 40826
rect 39298 40774 39310 40826
rect 39362 40774 39374 40826
rect 39426 40774 39438 40826
rect 39490 40774 49246 40826
rect 49298 40774 49310 40826
rect 49362 40774 49374 40826
rect 49426 40774 49438 40826
rect 49490 40774 59246 40826
rect 59298 40774 59310 40826
rect 59362 40774 59374 40826
rect 59426 40774 59438 40826
rect 59490 40774 68816 40826
rect 1104 40752 68816 40774
rect 1854 40712 1860 40724
rect 1815 40684 1860 40712
rect 1854 40672 1860 40684
rect 1912 40672 1918 40724
rect 17494 40672 17500 40724
rect 17552 40712 17558 40724
rect 17954 40712 17960 40724
rect 17552 40684 17960 40712
rect 17552 40672 17558 40684
rect 17954 40672 17960 40684
rect 18012 40712 18018 40724
rect 50890 40712 50896 40724
rect 18012 40684 50896 40712
rect 18012 40672 18018 40684
rect 50890 40672 50896 40684
rect 50948 40712 50954 40724
rect 65702 40712 65708 40724
rect 50948 40684 65708 40712
rect 50948 40672 50954 40684
rect 65702 40672 65708 40684
rect 65760 40672 65766 40724
rect 1949 40579 2007 40585
rect 1949 40545 1961 40579
rect 1995 40576 2007 40579
rect 2406 40576 2412 40588
rect 1995 40548 2412 40576
rect 1995 40545 2007 40548
rect 1949 40539 2007 40545
rect 2406 40536 2412 40548
rect 2464 40536 2470 40588
rect 22922 40576 22928 40588
rect 22883 40548 22928 40576
rect 22922 40536 22928 40548
rect 22980 40576 22986 40588
rect 23569 40579 23627 40585
rect 23569 40576 23581 40579
rect 22980 40548 23581 40576
rect 22980 40536 22986 40548
rect 23569 40545 23581 40548
rect 23615 40545 23627 40579
rect 23569 40539 23627 40545
rect 39114 40468 39120 40520
rect 39172 40508 39178 40520
rect 39850 40508 39856 40520
rect 39172 40480 39856 40508
rect 39172 40468 39178 40480
rect 39850 40468 39856 40480
rect 39908 40468 39914 40520
rect 2406 40332 2412 40384
rect 2464 40372 2470 40384
rect 2501 40375 2559 40381
rect 2501 40372 2513 40375
rect 2464 40344 2513 40372
rect 2464 40332 2470 40344
rect 2501 40341 2513 40344
rect 2547 40341 2559 40375
rect 23014 40372 23020 40384
rect 22975 40344 23020 40372
rect 2501 40335 2559 40341
rect 23014 40332 23020 40344
rect 23072 40332 23078 40384
rect 1104 40282 68816 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 14246 40282
rect 14298 40230 14310 40282
rect 14362 40230 14374 40282
rect 14426 40230 14438 40282
rect 14490 40230 24246 40282
rect 24298 40230 24310 40282
rect 24362 40230 24374 40282
rect 24426 40230 24438 40282
rect 24490 40230 34246 40282
rect 34298 40230 34310 40282
rect 34362 40230 34374 40282
rect 34426 40230 34438 40282
rect 34490 40230 44246 40282
rect 44298 40230 44310 40282
rect 44362 40230 44374 40282
rect 44426 40230 44438 40282
rect 44490 40230 54246 40282
rect 54298 40230 54310 40282
rect 54362 40230 54374 40282
rect 54426 40230 54438 40282
rect 54490 40230 64246 40282
rect 64298 40230 64310 40282
rect 64362 40230 64374 40282
rect 64426 40230 64438 40282
rect 64490 40230 68816 40282
rect 1104 40208 68816 40230
rect 67453 39967 67511 39973
rect 67453 39933 67465 39967
rect 67499 39964 67511 39967
rect 68094 39964 68100 39976
rect 67499 39936 68100 39964
rect 67499 39933 67511 39936
rect 67453 39927 67511 39933
rect 68094 39924 68100 39936
rect 68152 39924 68158 39976
rect 1104 39738 68816 39760
rect 1104 39686 9246 39738
rect 9298 39686 9310 39738
rect 9362 39686 9374 39738
rect 9426 39686 9438 39738
rect 9490 39686 19246 39738
rect 19298 39686 19310 39738
rect 19362 39686 19374 39738
rect 19426 39686 19438 39738
rect 19490 39686 29246 39738
rect 29298 39686 29310 39738
rect 29362 39686 29374 39738
rect 29426 39686 29438 39738
rect 29490 39686 39246 39738
rect 39298 39686 39310 39738
rect 39362 39686 39374 39738
rect 39426 39686 39438 39738
rect 39490 39686 49246 39738
rect 49298 39686 49310 39738
rect 49362 39686 49374 39738
rect 49426 39686 49438 39738
rect 49490 39686 59246 39738
rect 59298 39686 59310 39738
rect 59362 39686 59374 39738
rect 59426 39686 59438 39738
rect 59490 39686 68816 39738
rect 1104 39664 68816 39686
rect 2590 39624 2596 39636
rect 2551 39596 2596 39624
rect 2590 39584 2596 39596
rect 2648 39584 2654 39636
rect 1949 39559 2007 39565
rect 1949 39525 1961 39559
rect 1995 39556 2007 39559
rect 2608 39556 2636 39584
rect 1995 39528 2636 39556
rect 1995 39525 2007 39528
rect 1949 39519 2007 39525
rect 1762 39488 1768 39500
rect 1723 39460 1768 39488
rect 1762 39448 1768 39460
rect 1820 39448 1826 39500
rect 9766 39380 9772 39432
rect 9824 39420 9830 39432
rect 64782 39420 64788 39432
rect 9824 39392 64788 39420
rect 9824 39380 9830 39392
rect 64782 39380 64788 39392
rect 64840 39380 64846 39432
rect 2682 39312 2688 39364
rect 2740 39352 2746 39364
rect 66990 39352 66996 39364
rect 2740 39324 66996 39352
rect 2740 39312 2746 39324
rect 66990 39312 66996 39324
rect 67048 39312 67054 39364
rect 28994 39244 29000 39296
rect 29052 39284 29058 39296
rect 29365 39287 29423 39293
rect 29365 39284 29377 39287
rect 29052 39256 29377 39284
rect 29052 39244 29058 39256
rect 29365 39253 29377 39256
rect 29411 39253 29423 39287
rect 29365 39247 29423 39253
rect 33410 39244 33416 39296
rect 33468 39284 33474 39296
rect 33505 39287 33563 39293
rect 33505 39284 33517 39287
rect 33468 39256 33517 39284
rect 33468 39244 33474 39256
rect 33505 39253 33517 39256
rect 33551 39284 33563 39287
rect 33686 39284 33692 39296
rect 33551 39256 33692 39284
rect 33551 39253 33563 39256
rect 33505 39247 33563 39253
rect 33686 39244 33692 39256
rect 33744 39244 33750 39296
rect 1104 39194 68816 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 14246 39194
rect 14298 39142 14310 39194
rect 14362 39142 14374 39194
rect 14426 39142 14438 39194
rect 14490 39142 24246 39194
rect 24298 39142 24310 39194
rect 24362 39142 24374 39194
rect 24426 39142 24438 39194
rect 24490 39142 34246 39194
rect 34298 39142 34310 39194
rect 34362 39142 34374 39194
rect 34426 39142 34438 39194
rect 34490 39142 44246 39194
rect 44298 39142 44310 39194
rect 44362 39142 44374 39194
rect 44426 39142 44438 39194
rect 44490 39142 54246 39194
rect 54298 39142 54310 39194
rect 54362 39142 54374 39194
rect 54426 39142 54438 39194
rect 54490 39142 64246 39194
rect 64298 39142 64310 39194
rect 64362 39142 64374 39194
rect 64426 39142 64438 39194
rect 64490 39142 68816 39194
rect 1104 39120 68816 39142
rect 33134 38972 33140 39024
rect 33192 39012 33198 39024
rect 33594 39012 33600 39024
rect 33192 38984 33600 39012
rect 33192 38972 33198 38984
rect 33594 38972 33600 38984
rect 33652 39012 33658 39024
rect 34241 39015 34299 39021
rect 34241 39012 34253 39015
rect 33652 38984 34253 39012
rect 33652 38972 33658 38984
rect 34241 38981 34253 38984
rect 34287 38981 34299 39015
rect 34241 38975 34299 38981
rect 33686 38904 33692 38956
rect 33744 38944 33750 38956
rect 34333 38947 34391 38953
rect 34333 38944 34345 38947
rect 33744 38916 34345 38944
rect 33744 38904 33750 38916
rect 34333 38913 34345 38916
rect 34379 38913 34391 38947
rect 34333 38907 34391 38913
rect 34112 38879 34170 38885
rect 34112 38845 34124 38879
rect 34158 38876 34170 38879
rect 48961 38879 49019 38885
rect 34158 38848 35296 38876
rect 34158 38845 34170 38848
rect 34112 38839 34170 38845
rect 33965 38811 34023 38817
rect 33965 38808 33977 38811
rect 33428 38780 33977 38808
rect 17034 38700 17040 38752
rect 17092 38740 17098 38752
rect 33428 38749 33456 38780
rect 33965 38777 33977 38780
rect 34011 38777 34023 38811
rect 34698 38808 34704 38820
rect 34659 38780 34704 38808
rect 33965 38771 34023 38777
rect 34698 38768 34704 38780
rect 34756 38768 34762 38820
rect 35268 38749 35296 38848
rect 48961 38845 48973 38879
rect 49007 38876 49019 38879
rect 63310 38876 63316 38888
rect 49007 38848 63316 38876
rect 49007 38845 49019 38848
rect 48961 38839 49019 38845
rect 63310 38836 63316 38848
rect 63368 38836 63374 38888
rect 33413 38743 33471 38749
rect 33413 38740 33425 38743
rect 17092 38712 33425 38740
rect 17092 38700 17098 38712
rect 33413 38709 33425 38712
rect 33459 38709 33471 38743
rect 33413 38703 33471 38709
rect 35253 38743 35311 38749
rect 35253 38709 35265 38743
rect 35299 38740 35311 38743
rect 55674 38740 55680 38752
rect 35299 38712 55680 38740
rect 35299 38709 35311 38712
rect 35253 38703 35311 38709
rect 55674 38700 55680 38712
rect 55732 38700 55738 38752
rect 1104 38650 68816 38672
rect 1104 38598 9246 38650
rect 9298 38598 9310 38650
rect 9362 38598 9374 38650
rect 9426 38598 9438 38650
rect 9490 38598 19246 38650
rect 19298 38598 19310 38650
rect 19362 38598 19374 38650
rect 19426 38598 19438 38650
rect 19490 38598 29246 38650
rect 29298 38598 29310 38650
rect 29362 38598 29374 38650
rect 29426 38598 29438 38650
rect 29490 38598 39246 38650
rect 39298 38598 39310 38650
rect 39362 38598 39374 38650
rect 39426 38598 39438 38650
rect 39490 38598 49246 38650
rect 49298 38598 49310 38650
rect 49362 38598 49374 38650
rect 49426 38598 49438 38650
rect 49490 38598 59246 38650
rect 59298 38598 59310 38650
rect 59362 38598 59374 38650
rect 59426 38598 59438 38650
rect 59490 38598 68816 38650
rect 1104 38576 68816 38598
rect 40770 38496 40776 38548
rect 40828 38536 40834 38548
rect 43714 38536 43720 38548
rect 40828 38508 43720 38536
rect 40828 38496 40834 38508
rect 43714 38496 43720 38508
rect 43772 38496 43778 38548
rect 33594 38196 33600 38208
rect 33555 38168 33600 38196
rect 33594 38156 33600 38168
rect 33652 38156 33658 38208
rect 40954 38196 40960 38208
rect 40915 38168 40960 38196
rect 40954 38156 40960 38168
rect 41012 38156 41018 38208
rect 1104 38106 68816 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 14246 38106
rect 14298 38054 14310 38106
rect 14362 38054 14374 38106
rect 14426 38054 14438 38106
rect 14490 38054 24246 38106
rect 24298 38054 24310 38106
rect 24362 38054 24374 38106
rect 24426 38054 24438 38106
rect 24490 38054 34246 38106
rect 34298 38054 34310 38106
rect 34362 38054 34374 38106
rect 34426 38054 34438 38106
rect 34490 38054 44246 38106
rect 44298 38054 44310 38106
rect 44362 38054 44374 38106
rect 44426 38054 44438 38106
rect 44490 38054 54246 38106
rect 54298 38054 54310 38106
rect 54362 38054 54374 38106
rect 54426 38054 54438 38106
rect 54490 38054 64246 38106
rect 64298 38054 64310 38106
rect 64362 38054 64374 38106
rect 64426 38054 64438 38106
rect 64490 38054 68816 38106
rect 1104 38032 68816 38054
rect 5718 37952 5724 38004
rect 5776 37992 5782 38004
rect 40954 37992 40960 38004
rect 5776 37964 40960 37992
rect 5776 37952 5782 37964
rect 40954 37952 40960 37964
rect 41012 37952 41018 38004
rect 12802 37884 12808 37936
rect 12860 37924 12866 37936
rect 28994 37924 29000 37936
rect 12860 37896 29000 37924
rect 12860 37884 12866 37896
rect 28994 37884 29000 37896
rect 29052 37884 29058 37936
rect 46109 37927 46167 37933
rect 46109 37924 46121 37927
rect 31726 37896 46121 37924
rect 4890 37748 4896 37800
rect 4948 37788 4954 37800
rect 4948 37760 26234 37788
rect 4948 37748 4954 37760
rect 26206 37720 26234 37760
rect 31726 37720 31754 37896
rect 46109 37893 46121 37896
rect 46155 37893 46167 37927
rect 46109 37887 46167 37893
rect 35713 37791 35771 37797
rect 35713 37757 35725 37791
rect 35759 37757 35771 37791
rect 40678 37788 40684 37800
rect 40639 37760 40684 37788
rect 35713 37751 35771 37757
rect 26206 37692 31754 37720
rect 35728 37720 35756 37751
rect 40678 37748 40684 37760
rect 40736 37748 40742 37800
rect 62206 37720 62212 37732
rect 35728 37692 62212 37720
rect 62206 37680 62212 37692
rect 62264 37680 62270 37732
rect 66898 37680 66904 37732
rect 66956 37720 66962 37732
rect 67913 37723 67971 37729
rect 67913 37720 67925 37723
rect 66956 37692 67925 37720
rect 66956 37680 66962 37692
rect 67913 37689 67925 37692
rect 67959 37689 67971 37723
rect 68094 37720 68100 37732
rect 68055 37692 68100 37720
rect 67913 37683 67971 37689
rect 68094 37680 68100 37692
rect 68152 37680 68158 37732
rect 1104 37562 68816 37584
rect 1104 37510 9246 37562
rect 9298 37510 9310 37562
rect 9362 37510 9374 37562
rect 9426 37510 9438 37562
rect 9490 37510 19246 37562
rect 19298 37510 19310 37562
rect 19362 37510 19374 37562
rect 19426 37510 19438 37562
rect 19490 37510 29246 37562
rect 29298 37510 29310 37562
rect 29362 37510 29374 37562
rect 29426 37510 29438 37562
rect 29490 37510 39246 37562
rect 39298 37510 39310 37562
rect 39362 37510 39374 37562
rect 39426 37510 39438 37562
rect 39490 37510 49246 37562
rect 49298 37510 49310 37562
rect 49362 37510 49374 37562
rect 49426 37510 49438 37562
rect 49490 37510 59246 37562
rect 59298 37510 59310 37562
rect 59362 37510 59374 37562
rect 59426 37510 59438 37562
rect 59490 37510 68816 37562
rect 1104 37488 68816 37510
rect 1104 37018 68816 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 14246 37018
rect 14298 36966 14310 37018
rect 14362 36966 14374 37018
rect 14426 36966 14438 37018
rect 14490 36966 24246 37018
rect 24298 36966 24310 37018
rect 24362 36966 24374 37018
rect 24426 36966 24438 37018
rect 24490 36966 34246 37018
rect 34298 36966 34310 37018
rect 34362 36966 34374 37018
rect 34426 36966 34438 37018
rect 34490 36966 44246 37018
rect 44298 36966 44310 37018
rect 44362 36966 44374 37018
rect 44426 36966 44438 37018
rect 44490 36966 54246 37018
rect 54298 36966 54310 37018
rect 54362 36966 54374 37018
rect 54426 36966 54438 37018
rect 54490 36966 64246 37018
rect 64298 36966 64310 37018
rect 64362 36966 64374 37018
rect 64426 36966 64438 37018
rect 64490 36966 68816 37018
rect 1104 36944 68816 36966
rect 1578 36700 1584 36712
rect 1539 36672 1584 36700
rect 1578 36660 1584 36672
rect 1636 36700 1642 36712
rect 2041 36703 2099 36709
rect 2041 36700 2053 36703
rect 1636 36672 2053 36700
rect 1636 36660 1642 36672
rect 2041 36669 2053 36672
rect 2087 36669 2099 36703
rect 2041 36663 2099 36669
rect 1104 36474 68816 36496
rect 1104 36422 9246 36474
rect 9298 36422 9310 36474
rect 9362 36422 9374 36474
rect 9426 36422 9438 36474
rect 9490 36422 19246 36474
rect 19298 36422 19310 36474
rect 19362 36422 19374 36474
rect 19426 36422 19438 36474
rect 19490 36422 29246 36474
rect 29298 36422 29310 36474
rect 29362 36422 29374 36474
rect 29426 36422 29438 36474
rect 29490 36422 39246 36474
rect 39298 36422 39310 36474
rect 39362 36422 39374 36474
rect 39426 36422 39438 36474
rect 39490 36422 49246 36474
rect 49298 36422 49310 36474
rect 49362 36422 49374 36474
rect 49426 36422 49438 36474
rect 49490 36422 59246 36474
rect 59298 36422 59310 36474
rect 59362 36422 59374 36474
rect 59426 36422 59438 36474
rect 59490 36422 68816 36474
rect 1104 36400 68816 36422
rect 5537 36227 5595 36233
rect 5537 36193 5549 36227
rect 5583 36224 5595 36227
rect 59538 36224 59544 36236
rect 5583 36196 59544 36224
rect 5583 36193 5595 36196
rect 5537 36187 5595 36193
rect 59538 36184 59544 36196
rect 59596 36184 59602 36236
rect 66990 36184 66996 36236
rect 67048 36224 67054 36236
rect 67361 36227 67419 36233
rect 67361 36224 67373 36227
rect 67048 36196 67373 36224
rect 67048 36184 67054 36196
rect 67361 36193 67373 36196
rect 67407 36224 67419 36227
rect 67913 36227 67971 36233
rect 67913 36224 67925 36227
rect 67407 36196 67925 36224
rect 67407 36193 67419 36196
rect 67361 36187 67419 36193
rect 67913 36193 67925 36196
rect 67959 36193 67971 36227
rect 68094 36224 68100 36236
rect 68055 36196 68100 36224
rect 67913 36187 67971 36193
rect 68094 36184 68100 36196
rect 68152 36184 68158 36236
rect 41598 36116 41604 36168
rect 41656 36156 41662 36168
rect 41785 36159 41843 36165
rect 41785 36156 41797 36159
rect 41656 36128 41797 36156
rect 41656 36116 41662 36128
rect 41785 36125 41797 36128
rect 41831 36125 41843 36159
rect 42058 36156 42064 36168
rect 42019 36128 42064 36156
rect 41785 36119 41843 36125
rect 42058 36116 42064 36128
rect 42116 36116 42122 36168
rect 2866 36020 2872 36032
rect 2827 35992 2872 36020
rect 2866 35980 2872 35992
rect 2924 35980 2930 36032
rect 38194 35980 38200 36032
rect 38252 36020 38258 36032
rect 41233 36023 41291 36029
rect 41233 36020 41245 36023
rect 38252 35992 41245 36020
rect 38252 35980 38258 35992
rect 41233 35989 41245 35992
rect 41279 36020 41291 36023
rect 42058 36020 42064 36032
rect 41279 35992 42064 36020
rect 41279 35989 41291 35992
rect 41233 35983 41291 35989
rect 42058 35980 42064 35992
rect 42116 35980 42122 36032
rect 43162 36020 43168 36032
rect 43123 35992 43168 36020
rect 43162 35980 43168 35992
rect 43220 35980 43226 36032
rect 51258 35980 51264 36032
rect 51316 36020 51322 36032
rect 51445 36023 51503 36029
rect 51445 36020 51457 36023
rect 51316 35992 51457 36020
rect 51316 35980 51322 35992
rect 51445 35989 51457 35992
rect 51491 35989 51503 36023
rect 51445 35983 51503 35989
rect 1104 35930 68816 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 14246 35930
rect 14298 35878 14310 35930
rect 14362 35878 14374 35930
rect 14426 35878 14438 35930
rect 14490 35878 24246 35930
rect 24298 35878 24310 35930
rect 24362 35878 24374 35930
rect 24426 35878 24438 35930
rect 24490 35878 34246 35930
rect 34298 35878 34310 35930
rect 34362 35878 34374 35930
rect 34426 35878 34438 35930
rect 34490 35878 44246 35930
rect 44298 35878 44310 35930
rect 44362 35878 44374 35930
rect 44426 35878 44438 35930
rect 44490 35878 54246 35930
rect 54298 35878 54310 35930
rect 54362 35878 54374 35930
rect 54426 35878 54438 35930
rect 54490 35878 64246 35930
rect 64298 35878 64310 35930
rect 64362 35878 64374 35930
rect 64426 35878 64438 35930
rect 64490 35878 68816 35930
rect 1104 35856 68816 35878
rect 59998 35776 60004 35828
rect 60056 35816 60062 35828
rect 61562 35816 61568 35828
rect 60056 35788 61568 35816
rect 60056 35776 60062 35788
rect 61562 35776 61568 35788
rect 61620 35776 61626 35828
rect 58710 35708 58716 35760
rect 58768 35748 58774 35760
rect 60918 35748 60924 35760
rect 58768 35720 60924 35748
rect 58768 35708 58774 35720
rect 60918 35708 60924 35720
rect 60976 35708 60982 35760
rect 5350 35640 5356 35692
rect 5408 35680 5414 35692
rect 67910 35680 67916 35692
rect 5408 35652 67916 35680
rect 5408 35640 5414 35652
rect 67910 35640 67916 35652
rect 67968 35640 67974 35692
rect 1762 35612 1768 35624
rect 1723 35584 1768 35612
rect 1762 35572 1768 35584
rect 1820 35572 1826 35624
rect 7190 35612 7196 35624
rect 7151 35584 7196 35612
rect 7190 35572 7196 35584
rect 7248 35572 7254 35624
rect 44453 35615 44511 35621
rect 44453 35581 44465 35615
rect 44499 35612 44511 35615
rect 50154 35612 50160 35624
rect 44499 35584 50160 35612
rect 44499 35581 44511 35584
rect 44453 35575 44511 35581
rect 50154 35572 50160 35584
rect 50212 35572 50218 35624
rect 55861 35615 55919 35621
rect 55861 35581 55873 35615
rect 55907 35612 55919 35615
rect 60366 35612 60372 35624
rect 55907 35584 60372 35612
rect 55907 35581 55919 35584
rect 55861 35575 55919 35581
rect 60366 35572 60372 35584
rect 60424 35572 60430 35624
rect 61289 35615 61347 35621
rect 61289 35612 61301 35615
rect 60844 35584 61301 35612
rect 1949 35547 2007 35553
rect 1949 35513 1961 35547
rect 1995 35513 2007 35547
rect 1949 35507 2007 35513
rect 1964 35476 1992 35507
rect 2593 35479 2651 35485
rect 2593 35476 2605 35479
rect 1964 35448 2605 35476
rect 2593 35445 2605 35448
rect 2639 35476 2651 35479
rect 10318 35476 10324 35488
rect 2639 35448 10324 35476
rect 2639 35445 2651 35448
rect 2593 35439 2651 35445
rect 10318 35436 10324 35448
rect 10376 35436 10382 35488
rect 41509 35479 41567 35485
rect 41509 35445 41521 35479
rect 41555 35476 41567 35479
rect 41598 35476 41604 35488
rect 41555 35448 41604 35476
rect 41555 35445 41567 35448
rect 41509 35439 41567 35445
rect 41598 35436 41604 35448
rect 41656 35476 41662 35488
rect 60737 35479 60795 35485
rect 60737 35476 60749 35479
rect 41656 35448 60749 35476
rect 41656 35436 41662 35448
rect 60737 35445 60749 35448
rect 60783 35476 60795 35479
rect 60844 35476 60872 35584
rect 61289 35581 61301 35584
rect 61335 35581 61347 35615
rect 61562 35612 61568 35624
rect 61523 35584 61568 35612
rect 61289 35575 61347 35581
rect 61562 35572 61568 35584
rect 61620 35572 61626 35624
rect 67453 35615 67511 35621
rect 67453 35581 67465 35615
rect 67499 35612 67511 35615
rect 68097 35615 68155 35621
rect 68097 35612 68109 35615
rect 67499 35584 68109 35612
rect 67499 35581 67511 35584
rect 67453 35575 67511 35581
rect 68097 35581 68109 35584
rect 68143 35612 68155 35615
rect 68925 35615 68983 35621
rect 68925 35612 68937 35615
rect 68143 35584 68937 35612
rect 68143 35581 68155 35584
rect 68097 35575 68155 35581
rect 68925 35581 68937 35584
rect 68971 35581 68983 35615
rect 68925 35575 68983 35581
rect 60783 35448 60872 35476
rect 60783 35445 60795 35448
rect 60737 35439 60795 35445
rect 60918 35436 60924 35488
rect 60976 35476 60982 35488
rect 62669 35479 62727 35485
rect 62669 35476 62681 35479
rect 60976 35448 62681 35476
rect 60976 35436 60982 35448
rect 62669 35445 62681 35448
rect 62715 35445 62727 35479
rect 62669 35439 62727 35445
rect 1104 35386 68816 35408
rect 1104 35334 9246 35386
rect 9298 35334 9310 35386
rect 9362 35334 9374 35386
rect 9426 35334 9438 35386
rect 9490 35334 19246 35386
rect 19298 35334 19310 35386
rect 19362 35334 19374 35386
rect 19426 35334 19438 35386
rect 19490 35334 29246 35386
rect 29298 35334 29310 35386
rect 29362 35334 29374 35386
rect 29426 35334 29438 35386
rect 29490 35334 39246 35386
rect 39298 35334 39310 35386
rect 39362 35334 39374 35386
rect 39426 35334 39438 35386
rect 39490 35334 49246 35386
rect 49298 35334 49310 35386
rect 49362 35334 49374 35386
rect 49426 35334 49438 35386
rect 49490 35334 59246 35386
rect 59298 35334 59310 35386
rect 59362 35334 59374 35386
rect 59426 35334 59438 35386
rect 59490 35334 68816 35386
rect 1104 35312 68816 35334
rect 2498 35164 2504 35216
rect 2556 35204 2562 35216
rect 44082 35204 44088 35216
rect 2556 35176 44088 35204
rect 2556 35164 2562 35176
rect 44082 35164 44088 35176
rect 44140 35164 44146 35216
rect 60366 35164 60372 35216
rect 60424 35204 60430 35216
rect 65886 35204 65892 35216
rect 60424 35176 65892 35204
rect 60424 35164 60430 35176
rect 65886 35164 65892 35176
rect 65944 35164 65950 35216
rect 1302 35096 1308 35148
rect 1360 35136 1366 35148
rect 30929 35139 30987 35145
rect 30929 35136 30941 35139
rect 1360 35108 30941 35136
rect 1360 35096 1366 35108
rect 30929 35105 30941 35108
rect 30975 35136 30987 35139
rect 31481 35139 31539 35145
rect 31481 35136 31493 35139
rect 30975 35108 31493 35136
rect 30975 35105 30987 35108
rect 30929 35099 30987 35105
rect 31481 35105 31493 35108
rect 31527 35105 31539 35139
rect 31481 35099 31539 35105
rect 32950 35096 32956 35148
rect 33008 35136 33014 35148
rect 36446 35136 36452 35148
rect 33008 35108 36452 35136
rect 33008 35096 33014 35108
rect 36446 35096 36452 35108
rect 36504 35096 36510 35148
rect 67910 35136 67916 35148
rect 67871 35108 67916 35136
rect 67910 35096 67916 35108
rect 67968 35096 67974 35148
rect 9030 35028 9036 35080
rect 9088 35068 9094 35080
rect 39942 35068 39948 35080
rect 9088 35040 39948 35068
rect 9088 35028 9094 35040
rect 39942 35028 39948 35040
rect 40000 35028 40006 35080
rect 8386 34960 8392 35012
rect 8444 35000 8450 35012
rect 12986 35000 12992 35012
rect 8444 34972 12992 35000
rect 8444 34960 8450 34972
rect 12986 34960 12992 34972
rect 13044 34960 13050 35012
rect 35066 34960 35072 35012
rect 35124 35000 35130 35012
rect 67818 35000 67824 35012
rect 35124 34972 67824 35000
rect 35124 34960 35130 34972
rect 67818 34960 67824 34972
rect 67876 34960 67882 35012
rect 6086 34892 6092 34944
rect 6144 34932 6150 34944
rect 11606 34932 11612 34944
rect 6144 34904 11612 34932
rect 6144 34892 6150 34904
rect 11606 34892 11612 34904
rect 11664 34892 11670 34944
rect 30558 34892 30564 34944
rect 30616 34932 30622 34944
rect 32769 34935 32827 34941
rect 32769 34932 32781 34935
rect 30616 34904 32781 34932
rect 30616 34892 30622 34904
rect 32769 34901 32781 34904
rect 32815 34901 32827 34935
rect 32769 34895 32827 34901
rect 34790 34892 34796 34944
rect 34848 34932 34854 34944
rect 56042 34932 56048 34944
rect 34848 34904 56048 34932
rect 34848 34892 34854 34904
rect 56042 34892 56048 34904
rect 56100 34892 56106 34944
rect 57882 34892 57888 34944
rect 57940 34932 57946 34944
rect 60829 34935 60887 34941
rect 60829 34932 60841 34935
rect 57940 34904 60841 34932
rect 57940 34892 57946 34904
rect 60829 34901 60841 34904
rect 60875 34901 60887 34935
rect 68922 34932 68928 34944
rect 68883 34904 68928 34932
rect 60829 34895 60887 34901
rect 68922 34892 68928 34904
rect 68980 34892 68986 34944
rect 1104 34842 68816 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 14246 34842
rect 14298 34790 14310 34842
rect 14362 34790 14374 34842
rect 14426 34790 14438 34842
rect 14490 34790 24246 34842
rect 24298 34790 24310 34842
rect 24362 34790 24374 34842
rect 24426 34790 24438 34842
rect 24490 34790 34246 34842
rect 34298 34790 34310 34842
rect 34362 34790 34374 34842
rect 34426 34790 34438 34842
rect 34490 34790 44246 34842
rect 44298 34790 44310 34842
rect 44362 34790 44374 34842
rect 44426 34790 44438 34842
rect 44490 34790 54246 34842
rect 54298 34790 54310 34842
rect 54362 34790 54374 34842
rect 54426 34790 54438 34842
rect 54490 34790 64246 34842
rect 64298 34790 64310 34842
rect 64362 34790 64374 34842
rect 64426 34790 64438 34842
rect 64490 34790 68816 34842
rect 1104 34768 68816 34790
rect 7098 34688 7104 34740
rect 7156 34728 7162 34740
rect 8386 34728 8392 34740
rect 7156 34700 7788 34728
rect 8347 34700 8392 34728
rect 7156 34688 7162 34700
rect 7760 34660 7788 34700
rect 8386 34688 8392 34700
rect 8444 34688 8450 34740
rect 9030 34728 9036 34740
rect 8991 34700 9036 34728
rect 9030 34688 9036 34700
rect 9088 34688 9094 34740
rect 57882 34728 57888 34740
rect 9140 34700 57888 34728
rect 9140 34660 9168 34700
rect 57882 34688 57888 34700
rect 57940 34688 57946 34740
rect 64693 34731 64751 34737
rect 64693 34697 64705 34731
rect 64739 34728 64751 34731
rect 66806 34728 66812 34740
rect 64739 34700 66812 34728
rect 64739 34697 64751 34700
rect 64693 34691 64751 34697
rect 66806 34688 66812 34700
rect 66864 34688 66870 34740
rect 32030 34660 32036 34672
rect 7760 34632 9168 34660
rect 31991 34632 32036 34660
rect 32030 34620 32036 34632
rect 32088 34620 32094 34672
rect 33226 34620 33232 34672
rect 33284 34660 33290 34672
rect 33413 34663 33471 34669
rect 33413 34660 33425 34663
rect 33284 34632 33425 34660
rect 33284 34620 33290 34632
rect 33413 34629 33425 34632
rect 33459 34629 33471 34663
rect 33413 34623 33471 34629
rect 34885 34663 34943 34669
rect 34885 34629 34897 34663
rect 34931 34660 34943 34663
rect 35066 34660 35072 34672
rect 34931 34632 35072 34660
rect 34931 34629 34943 34632
rect 34885 34623 34943 34629
rect 35066 34620 35072 34632
rect 35124 34620 35130 34672
rect 36446 34620 36452 34672
rect 36504 34660 36510 34672
rect 67266 34660 67272 34672
rect 36504 34632 67272 34660
rect 36504 34620 36510 34632
rect 67266 34620 67272 34632
rect 67324 34620 67330 34672
rect 7101 34595 7159 34601
rect 7101 34561 7113 34595
rect 7147 34592 7159 34595
rect 9030 34592 9036 34604
rect 7147 34564 9036 34592
rect 7147 34561 7159 34564
rect 7101 34555 7159 34561
rect 9030 34552 9036 34564
rect 9088 34552 9094 34604
rect 11606 34552 11612 34604
rect 11664 34592 11670 34604
rect 32766 34592 32772 34604
rect 11664 34564 32772 34592
rect 11664 34552 11670 34564
rect 32766 34552 32772 34564
rect 32824 34552 32830 34604
rect 33134 34592 33140 34604
rect 33095 34564 33140 34592
rect 33134 34552 33140 34564
rect 33192 34552 33198 34604
rect 33870 34552 33876 34604
rect 33928 34592 33934 34604
rect 45097 34595 45155 34601
rect 45097 34592 45109 34595
rect 33928 34564 45109 34592
rect 33928 34552 33934 34564
rect 45097 34561 45109 34564
rect 45143 34561 45155 34595
rect 45097 34555 45155 34561
rect 6825 34527 6883 34533
rect 6825 34493 6837 34527
rect 6871 34524 6883 34527
rect 9582 34524 9588 34536
rect 6871 34496 9588 34524
rect 6871 34493 6883 34496
rect 6825 34487 6883 34493
rect 9582 34484 9588 34496
rect 9640 34484 9646 34536
rect 30285 34527 30343 34533
rect 30285 34493 30297 34527
rect 30331 34524 30343 34527
rect 32950 34524 32956 34536
rect 30331 34496 32956 34524
rect 30331 34493 30343 34496
rect 30285 34487 30343 34493
rect 32950 34484 32956 34496
rect 33008 34484 33014 34536
rect 33318 34484 33324 34536
rect 33376 34533 33382 34536
rect 33376 34527 33390 34533
rect 33378 34524 33390 34527
rect 33505 34527 33563 34533
rect 33378 34496 33421 34524
rect 33378 34493 33390 34496
rect 33376 34487 33390 34493
rect 33505 34493 33517 34527
rect 33551 34493 33563 34527
rect 33505 34487 33563 34493
rect 33597 34527 33655 34533
rect 33597 34493 33609 34527
rect 33643 34493 33655 34527
rect 33597 34487 33655 34493
rect 33781 34527 33839 34533
rect 33781 34493 33793 34527
rect 33827 34524 33839 34527
rect 35066 34524 35072 34536
rect 33827 34496 35072 34524
rect 33827 34493 33839 34496
rect 33781 34487 33839 34493
rect 33376 34484 33382 34487
rect 31754 34416 31760 34468
rect 31812 34456 31818 34468
rect 32030 34456 32036 34468
rect 31812 34428 32036 34456
rect 31812 34416 31818 34428
rect 32030 34416 32036 34428
rect 32088 34456 32094 34468
rect 33520 34456 33548 34487
rect 32088 34428 33548 34456
rect 32088 34416 32094 34428
rect 33134 34348 33140 34400
rect 33192 34388 33198 34400
rect 33612 34388 33640 34487
rect 35066 34484 35072 34496
rect 35124 34484 35130 34536
rect 44082 34484 44088 34536
rect 44140 34524 44146 34536
rect 44453 34527 44511 34533
rect 44453 34524 44465 34527
rect 44140 34496 44465 34524
rect 44140 34484 44146 34496
rect 44453 34493 44465 34496
rect 44499 34493 44511 34527
rect 44453 34487 44511 34493
rect 34241 34391 34299 34397
rect 34241 34388 34253 34391
rect 33192 34360 34253 34388
rect 33192 34348 33198 34360
rect 34241 34357 34253 34360
rect 34287 34388 34299 34391
rect 34790 34388 34796 34400
rect 34287 34360 34796 34388
rect 34287 34357 34299 34360
rect 34241 34351 34299 34357
rect 34790 34348 34796 34360
rect 34848 34348 34854 34400
rect 1104 34298 68816 34320
rect 1104 34246 9246 34298
rect 9298 34246 9310 34298
rect 9362 34246 9374 34298
rect 9426 34246 9438 34298
rect 9490 34246 19246 34298
rect 19298 34246 19310 34298
rect 19362 34246 19374 34298
rect 19426 34246 19438 34298
rect 19490 34246 29246 34298
rect 29298 34246 29310 34298
rect 29362 34246 29374 34298
rect 29426 34246 29438 34298
rect 29490 34246 39246 34298
rect 39298 34246 39310 34298
rect 39362 34246 39374 34298
rect 39426 34246 39438 34298
rect 39490 34246 49246 34298
rect 49298 34246 49310 34298
rect 49362 34246 49374 34298
rect 49426 34246 49438 34298
rect 49490 34246 59246 34298
rect 59298 34246 59310 34298
rect 59362 34246 59374 34298
rect 59426 34246 59438 34298
rect 59490 34246 68816 34298
rect 1104 34224 68816 34246
rect 1854 34184 1860 34196
rect 1815 34156 1860 34184
rect 1854 34144 1860 34156
rect 1912 34144 1918 34196
rect 32401 34187 32459 34193
rect 32401 34153 32413 34187
rect 32447 34184 32459 34187
rect 32490 34184 32496 34196
rect 32447 34156 32496 34184
rect 32447 34153 32459 34156
rect 32401 34147 32459 34153
rect 32490 34144 32496 34156
rect 32548 34184 32554 34196
rect 33318 34184 33324 34196
rect 32548 34156 33324 34184
rect 32548 34144 32554 34156
rect 33318 34144 33324 34156
rect 33376 34144 33382 34196
rect 32953 34119 33011 34125
rect 32953 34085 32965 34119
rect 32999 34116 33011 34119
rect 33226 34116 33232 34128
rect 32999 34088 33232 34116
rect 32999 34085 33011 34088
rect 32953 34079 33011 34085
rect 33226 34076 33232 34088
rect 33284 34116 33290 34128
rect 33778 34116 33784 34128
rect 33284 34088 33784 34116
rect 33284 34076 33290 34088
rect 33778 34076 33784 34088
rect 33836 34076 33842 34128
rect 1949 34051 2007 34057
rect 1949 34017 1961 34051
rect 1995 34048 2007 34051
rect 2130 34048 2136 34060
rect 1995 34020 2136 34048
rect 1995 34017 2007 34020
rect 1949 34011 2007 34017
rect 2130 34008 2136 34020
rect 2188 34008 2194 34060
rect 10134 34048 10140 34060
rect 10095 34020 10140 34048
rect 10134 34008 10140 34020
rect 10192 34008 10198 34060
rect 2130 33804 2136 33856
rect 2188 33844 2194 33856
rect 2501 33847 2559 33853
rect 2501 33844 2513 33847
rect 2188 33816 2513 33844
rect 2188 33804 2194 33816
rect 2501 33813 2513 33816
rect 2547 33813 2559 33847
rect 55306 33844 55312 33856
rect 55267 33816 55312 33844
rect 2501 33807 2559 33813
rect 55306 33804 55312 33816
rect 55364 33804 55370 33856
rect 1104 33754 68816 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 14246 33754
rect 14298 33702 14310 33754
rect 14362 33702 14374 33754
rect 14426 33702 14438 33754
rect 14490 33702 24246 33754
rect 24298 33702 24310 33754
rect 24362 33702 24374 33754
rect 24426 33702 24438 33754
rect 24490 33702 34246 33754
rect 34298 33702 34310 33754
rect 34362 33702 34374 33754
rect 34426 33702 34438 33754
rect 34490 33702 44246 33754
rect 44298 33702 44310 33754
rect 44362 33702 44374 33754
rect 44426 33702 44438 33754
rect 44490 33702 54246 33754
rect 54298 33702 54310 33754
rect 54362 33702 54374 33754
rect 54426 33702 54438 33754
rect 54490 33702 64246 33754
rect 64298 33702 64310 33754
rect 64362 33702 64374 33754
rect 64426 33702 64438 33754
rect 64490 33702 68816 33754
rect 1104 33680 68816 33702
rect 36909 33575 36967 33581
rect 36909 33541 36921 33575
rect 36955 33572 36967 33575
rect 36955 33544 41414 33572
rect 36955 33541 36967 33544
rect 36909 33535 36967 33541
rect 41386 33504 41414 33544
rect 67174 33504 67180 33516
rect 31726 33476 39436 33504
rect 41386 33476 67180 33504
rect 25133 33439 25191 33445
rect 25133 33405 25145 33439
rect 25179 33436 25191 33439
rect 31726 33436 31754 33476
rect 25179 33408 31754 33436
rect 39301 33439 39359 33445
rect 25179 33405 25191 33408
rect 25133 33399 25191 33405
rect 39301 33405 39313 33439
rect 39347 33405 39359 33439
rect 39408 33436 39436 33476
rect 67174 33464 67180 33476
rect 67232 33464 67238 33516
rect 57330 33436 57336 33448
rect 39408 33408 57336 33436
rect 39301 33399 39359 33405
rect 39316 33368 39344 33399
rect 57330 33396 57336 33408
rect 57388 33396 57394 33448
rect 62942 33436 62948 33448
rect 62903 33408 62948 33436
rect 62942 33396 62948 33408
rect 63000 33396 63006 33448
rect 62850 33368 62856 33380
rect 39316 33340 62856 33368
rect 62850 33328 62856 33340
rect 62908 33328 62914 33380
rect 1104 33210 68816 33232
rect 1104 33158 9246 33210
rect 9298 33158 9310 33210
rect 9362 33158 9374 33210
rect 9426 33158 9438 33210
rect 9490 33158 19246 33210
rect 19298 33158 19310 33210
rect 19362 33158 19374 33210
rect 19426 33158 19438 33210
rect 19490 33158 29246 33210
rect 29298 33158 29310 33210
rect 29362 33158 29374 33210
rect 29426 33158 29438 33210
rect 29490 33158 39246 33210
rect 39298 33158 39310 33210
rect 39362 33158 39374 33210
rect 39426 33158 39438 33210
rect 39490 33158 49246 33210
rect 49298 33158 49310 33210
rect 49362 33158 49374 33210
rect 49426 33158 49438 33210
rect 49490 33158 59246 33210
rect 59298 33158 59310 33210
rect 59362 33158 59374 33210
rect 59426 33158 59438 33210
rect 59490 33158 68816 33210
rect 1104 33136 68816 33158
rect 64874 32716 64880 32768
rect 64932 32756 64938 32768
rect 64932 32728 64977 32756
rect 64932 32716 64938 32728
rect 1104 32666 68816 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 14246 32666
rect 14298 32614 14310 32666
rect 14362 32614 14374 32666
rect 14426 32614 14438 32666
rect 14490 32614 24246 32666
rect 24298 32614 24310 32666
rect 24362 32614 24374 32666
rect 24426 32614 24438 32666
rect 24490 32614 34246 32666
rect 34298 32614 34310 32666
rect 34362 32614 34374 32666
rect 34426 32614 34438 32666
rect 34490 32614 44246 32666
rect 44298 32614 44310 32666
rect 44362 32614 44374 32666
rect 44426 32614 44438 32666
rect 44490 32614 54246 32666
rect 54298 32614 54310 32666
rect 54362 32614 54374 32666
rect 54426 32614 54438 32666
rect 54490 32614 64246 32666
rect 64298 32614 64310 32666
rect 64362 32614 64374 32666
rect 64426 32614 64438 32666
rect 64490 32614 68816 32666
rect 1104 32592 68816 32614
rect 49878 32444 49884 32496
rect 49936 32484 49942 32496
rect 62390 32484 62396 32496
rect 49936 32456 62396 32484
rect 49936 32444 49942 32456
rect 62390 32444 62396 32456
rect 62448 32444 62454 32496
rect 16758 32376 16764 32428
rect 16816 32416 16822 32428
rect 30466 32416 30472 32428
rect 16816 32388 30472 32416
rect 16816 32376 16822 32388
rect 30466 32376 30472 32388
rect 30524 32376 30530 32428
rect 41230 32376 41236 32428
rect 41288 32416 41294 32428
rect 65150 32416 65156 32428
rect 41288 32388 65156 32416
rect 41288 32376 41294 32388
rect 65150 32376 65156 32388
rect 65208 32376 65214 32428
rect 7009 32351 7067 32357
rect 7009 32317 7021 32351
rect 7055 32348 7067 32351
rect 17678 32348 17684 32360
rect 7055 32320 17684 32348
rect 7055 32317 7067 32320
rect 7009 32311 7067 32317
rect 17678 32308 17684 32320
rect 17736 32308 17742 32360
rect 66346 32240 66352 32292
rect 66404 32280 66410 32292
rect 67913 32283 67971 32289
rect 67913 32280 67925 32283
rect 66404 32252 67925 32280
rect 66404 32240 66410 32252
rect 67913 32249 67925 32252
rect 67959 32249 67971 32283
rect 68094 32280 68100 32292
rect 68055 32252 68100 32280
rect 67913 32243 67971 32249
rect 68094 32240 68100 32252
rect 68152 32240 68158 32292
rect 1104 32122 68816 32144
rect 1104 32070 9246 32122
rect 9298 32070 9310 32122
rect 9362 32070 9374 32122
rect 9426 32070 9438 32122
rect 9490 32070 19246 32122
rect 19298 32070 19310 32122
rect 19362 32070 19374 32122
rect 19426 32070 19438 32122
rect 19490 32070 29246 32122
rect 29298 32070 29310 32122
rect 29362 32070 29374 32122
rect 29426 32070 29438 32122
rect 29490 32070 39246 32122
rect 39298 32070 39310 32122
rect 39362 32070 39374 32122
rect 39426 32070 39438 32122
rect 39490 32070 49246 32122
rect 49298 32070 49310 32122
rect 49362 32070 49374 32122
rect 49426 32070 49438 32122
rect 49490 32070 59246 32122
rect 59298 32070 59310 32122
rect 59362 32070 59374 32122
rect 59426 32070 59438 32122
rect 59490 32070 68816 32122
rect 1104 32048 68816 32070
rect 39574 32008 39580 32020
rect 27540 31980 39580 32008
rect 1578 31872 1584 31884
rect 1539 31844 1584 31872
rect 1578 31832 1584 31844
rect 1636 31872 1642 31884
rect 2041 31875 2099 31881
rect 2041 31872 2053 31875
rect 1636 31844 2053 31872
rect 1636 31832 1642 31844
rect 2041 31841 2053 31844
rect 2087 31841 2099 31875
rect 26878 31872 26884 31884
rect 26839 31844 26884 31872
rect 2041 31835 2099 31841
rect 26878 31832 26884 31844
rect 26936 31832 26942 31884
rect 27540 31881 27568 31980
rect 39574 31968 39580 31980
rect 39632 31968 39638 32020
rect 42426 31968 42432 32020
rect 42484 32008 42490 32020
rect 61838 32008 61844 32020
rect 42484 31980 61844 32008
rect 42484 31968 42490 31980
rect 61838 31968 61844 31980
rect 61896 31968 61902 32020
rect 33778 31900 33784 31952
rect 33836 31940 33842 31952
rect 36630 31940 36636 31952
rect 33836 31912 36636 31940
rect 33836 31900 33842 31912
rect 36630 31900 36636 31912
rect 36688 31940 36694 31952
rect 39942 31940 39948 31952
rect 36688 31912 37412 31940
rect 36688 31900 36694 31912
rect 27525 31875 27583 31881
rect 27525 31841 27537 31875
rect 27571 31841 27583 31875
rect 27525 31835 27583 31841
rect 36998 31832 37004 31884
rect 37056 31872 37062 31884
rect 37185 31875 37243 31881
rect 37185 31872 37197 31875
rect 37056 31844 37197 31872
rect 37056 31832 37062 31844
rect 37185 31841 37197 31844
rect 37231 31841 37243 31875
rect 37185 31835 37243 31841
rect 37384 31804 37412 31912
rect 37476 31912 39948 31940
rect 37476 31881 37504 31912
rect 39942 31900 39948 31912
rect 40000 31900 40006 31952
rect 55401 31943 55459 31949
rect 55401 31940 55413 31943
rect 55186 31912 55413 31940
rect 37461 31875 37519 31881
rect 37461 31841 37473 31875
rect 37507 31841 37519 31875
rect 37461 31835 37519 31841
rect 37737 31875 37795 31881
rect 37737 31841 37749 31875
rect 37783 31841 37795 31875
rect 37737 31835 37795 31841
rect 37921 31875 37979 31881
rect 37921 31841 37933 31875
rect 37967 31872 37979 31875
rect 39025 31875 39083 31881
rect 39025 31872 39037 31875
rect 37967 31844 39037 31872
rect 37967 31841 37979 31844
rect 37921 31835 37979 31841
rect 39025 31841 39037 31844
rect 39071 31872 39083 31875
rect 43806 31872 43812 31884
rect 39071 31844 43812 31872
rect 39071 31841 39083 31844
rect 39025 31835 39083 31841
rect 37553 31807 37611 31813
rect 37553 31804 37565 31807
rect 37384 31776 37565 31804
rect 37553 31773 37565 31776
rect 37599 31773 37611 31807
rect 37752 31804 37780 31835
rect 43806 31832 43812 31844
rect 43864 31832 43870 31884
rect 47486 31832 47492 31884
rect 47544 31872 47550 31884
rect 54849 31875 54907 31881
rect 54849 31872 54861 31875
rect 47544 31844 54861 31872
rect 47544 31832 47550 31844
rect 54849 31841 54861 31844
rect 54895 31872 54907 31875
rect 55186 31872 55214 31912
rect 55401 31909 55413 31912
rect 55447 31909 55459 31943
rect 55401 31903 55459 31909
rect 55674 31900 55680 31952
rect 55732 31940 55738 31952
rect 55769 31943 55827 31949
rect 55769 31940 55781 31943
rect 55732 31912 55781 31940
rect 55732 31900 55738 31912
rect 55769 31909 55781 31912
rect 55815 31909 55827 31943
rect 55769 31903 55827 31909
rect 56413 31943 56471 31949
rect 56413 31909 56425 31943
rect 56459 31940 56471 31943
rect 58710 31940 58716 31952
rect 56459 31912 58716 31940
rect 56459 31909 56471 31912
rect 56413 31903 56471 31909
rect 54895 31844 55214 31872
rect 55585 31875 55643 31881
rect 54895 31841 54907 31844
rect 54849 31835 54907 31841
rect 55585 31841 55597 31875
rect 55631 31872 55643 31875
rect 56226 31872 56232 31884
rect 55631 31844 56232 31872
rect 55631 31841 55643 31844
rect 55585 31835 55643 31841
rect 56226 31832 56232 31844
rect 56284 31872 56290 31884
rect 56428 31872 56456 31903
rect 58710 31900 58716 31912
rect 58768 31900 58774 31952
rect 56284 31844 56456 31872
rect 56284 31832 56290 31844
rect 38473 31807 38531 31813
rect 38473 31804 38485 31807
rect 37752 31776 38485 31804
rect 37553 31767 37611 31773
rect 38473 31773 38485 31776
rect 38519 31804 38531 31807
rect 49878 31804 49884 31816
rect 38519 31776 49884 31804
rect 38519 31773 38531 31776
rect 38473 31767 38531 31773
rect 49878 31764 49884 31776
rect 49936 31764 49942 31816
rect 37642 31736 37648 31748
rect 37603 31708 37648 31736
rect 37642 31696 37648 31708
rect 37700 31696 37706 31748
rect 42426 31736 42432 31748
rect 42387 31708 42432 31736
rect 42426 31696 42432 31708
rect 42484 31696 42490 31748
rect 1104 31578 68816 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 14246 31578
rect 14298 31526 14310 31578
rect 14362 31526 14374 31578
rect 14426 31526 14438 31578
rect 14490 31526 24246 31578
rect 24298 31526 24310 31578
rect 24362 31526 24374 31578
rect 24426 31526 24438 31578
rect 24490 31526 34246 31578
rect 34298 31526 34310 31578
rect 34362 31526 34374 31578
rect 34426 31526 34438 31578
rect 34490 31526 44246 31578
rect 44298 31526 44310 31578
rect 44362 31526 44374 31578
rect 44426 31526 44438 31578
rect 44490 31526 54246 31578
rect 54298 31526 54310 31578
rect 54362 31526 54374 31578
rect 54426 31526 54438 31578
rect 54490 31526 64246 31578
rect 64298 31526 64310 31578
rect 64362 31526 64374 31578
rect 64426 31526 64438 31578
rect 64490 31526 68816 31578
rect 1104 31504 68816 31526
rect 31754 31424 31760 31476
rect 31812 31464 31818 31476
rect 36817 31467 36875 31473
rect 36817 31464 36829 31467
rect 31812 31436 36829 31464
rect 31812 31424 31818 31436
rect 36817 31433 36829 31436
rect 36863 31464 36875 31467
rect 37642 31464 37648 31476
rect 36863 31436 37648 31464
rect 36863 31433 36875 31436
rect 36817 31427 36875 31433
rect 37642 31424 37648 31436
rect 37700 31424 37706 31476
rect 1104 31034 68816 31056
rect 1104 30982 9246 31034
rect 9298 30982 9310 31034
rect 9362 30982 9374 31034
rect 9426 30982 9438 31034
rect 9490 30982 19246 31034
rect 19298 30982 19310 31034
rect 19362 30982 19374 31034
rect 19426 30982 19438 31034
rect 19490 30982 29246 31034
rect 29298 30982 29310 31034
rect 29362 30982 29374 31034
rect 29426 30982 29438 31034
rect 29490 30982 39246 31034
rect 39298 30982 39310 31034
rect 39362 30982 39374 31034
rect 39426 30982 39438 31034
rect 39490 30982 49246 31034
rect 49298 30982 49310 31034
rect 49362 30982 49374 31034
rect 49426 30982 49438 31034
rect 49490 30982 59246 31034
rect 59298 30982 59310 31034
rect 59362 30982 59374 31034
rect 59426 30982 59438 31034
rect 59490 30982 68816 31034
rect 1104 30960 68816 30982
rect 25961 30923 26019 30929
rect 25961 30889 25973 30923
rect 26007 30920 26019 30923
rect 30558 30920 30564 30932
rect 26007 30892 30564 30920
rect 26007 30889 26019 30892
rect 25961 30883 26019 30889
rect 8128 30824 22094 30852
rect 8128 30793 8156 30824
rect 8113 30787 8171 30793
rect 8113 30753 8125 30787
rect 8159 30753 8171 30787
rect 8113 30747 8171 30753
rect 22066 30716 22094 30824
rect 25409 30787 25467 30793
rect 25409 30753 25421 30787
rect 25455 30784 25467 30787
rect 25976 30784 26004 30883
rect 30558 30880 30564 30892
rect 30616 30880 30622 30932
rect 37090 30812 37096 30864
rect 37148 30852 37154 30864
rect 37829 30855 37887 30861
rect 37829 30852 37841 30855
rect 37148 30824 37841 30852
rect 37148 30812 37154 30824
rect 37829 30821 37841 30824
rect 37875 30852 37887 30855
rect 40310 30852 40316 30864
rect 37875 30824 40316 30852
rect 37875 30821 37887 30824
rect 37829 30815 37887 30821
rect 40310 30812 40316 30824
rect 40368 30812 40374 30864
rect 67542 30812 67548 30864
rect 67600 30852 67606 30864
rect 67913 30855 67971 30861
rect 67913 30852 67925 30855
rect 67600 30824 67925 30852
rect 67600 30812 67606 30824
rect 67913 30821 67925 30824
rect 67959 30821 67971 30855
rect 68094 30852 68100 30864
rect 68055 30824 68100 30852
rect 67913 30815 67971 30821
rect 68094 30812 68100 30824
rect 68152 30812 68158 30864
rect 25455 30756 26004 30784
rect 25455 30753 25467 30756
rect 25409 30747 25467 30753
rect 37642 30744 37648 30796
rect 37700 30793 37706 30796
rect 37700 30787 37743 30793
rect 37731 30753 37743 30787
rect 37700 30747 37743 30753
rect 37921 30787 37979 30793
rect 37921 30753 37933 30787
rect 37967 30753 37979 30787
rect 37921 30747 37979 30753
rect 38105 30787 38163 30793
rect 38105 30753 38117 30787
rect 38151 30784 38163 30787
rect 38654 30784 38660 30796
rect 38151 30756 38660 30784
rect 38151 30753 38163 30756
rect 38105 30747 38163 30753
rect 37700 30744 37706 30747
rect 36446 30716 36452 30728
rect 22066 30688 36452 30716
rect 36446 30676 36452 30688
rect 36504 30676 36510 30728
rect 37936 30716 37964 30747
rect 38654 30744 38660 30756
rect 38712 30784 38718 30796
rect 39114 30784 39120 30796
rect 38712 30756 39120 30784
rect 38712 30744 38718 30756
rect 39114 30744 39120 30756
rect 39172 30744 39178 30796
rect 36924 30688 37964 30716
rect 4433 30651 4491 30657
rect 4433 30617 4445 30651
rect 4479 30648 4491 30651
rect 10870 30648 10876 30660
rect 4479 30620 10876 30648
rect 4479 30617 4491 30620
rect 4433 30611 4491 30617
rect 10870 30608 10876 30620
rect 10928 30608 10934 30660
rect 25222 30580 25228 30592
rect 25183 30552 25228 30580
rect 25222 30540 25228 30552
rect 25280 30540 25286 30592
rect 33686 30540 33692 30592
rect 33744 30580 33750 30592
rect 36924 30589 36952 30688
rect 36909 30583 36967 30589
rect 36909 30580 36921 30583
rect 33744 30552 36921 30580
rect 33744 30540 33750 30552
rect 36909 30549 36921 30552
rect 36955 30549 36967 30583
rect 37550 30580 37556 30592
rect 37511 30552 37556 30580
rect 36909 30543 36967 30549
rect 37550 30540 37556 30552
rect 37608 30540 37614 30592
rect 37642 30540 37648 30592
rect 37700 30580 37706 30592
rect 38565 30583 38623 30589
rect 38565 30580 38577 30583
rect 37700 30552 38577 30580
rect 37700 30540 37706 30552
rect 38565 30549 38577 30552
rect 38611 30580 38623 30583
rect 48958 30580 48964 30592
rect 38611 30552 48964 30580
rect 38611 30549 38623 30552
rect 38565 30543 38623 30549
rect 48958 30540 48964 30552
rect 49016 30540 49022 30592
rect 1104 30490 68816 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 14246 30490
rect 14298 30438 14310 30490
rect 14362 30438 14374 30490
rect 14426 30438 14438 30490
rect 14490 30438 24246 30490
rect 24298 30438 24310 30490
rect 24362 30438 24374 30490
rect 24426 30438 24438 30490
rect 24490 30438 34246 30490
rect 34298 30438 34310 30490
rect 34362 30438 34374 30490
rect 34426 30438 34438 30490
rect 34490 30438 44246 30490
rect 44298 30438 44310 30490
rect 44362 30438 44374 30490
rect 44426 30438 44438 30490
rect 44490 30438 54246 30490
rect 54298 30438 54310 30490
rect 54362 30438 54374 30490
rect 54426 30438 54438 30490
rect 54490 30438 64246 30490
rect 64298 30438 64310 30490
rect 64362 30438 64374 30490
rect 64426 30438 64438 30490
rect 64490 30438 68816 30490
rect 1104 30416 68816 30438
rect 12986 30336 12992 30388
rect 13044 30376 13050 30388
rect 15194 30376 15200 30388
rect 13044 30348 15200 30376
rect 13044 30336 13050 30348
rect 15194 30336 15200 30348
rect 15252 30376 15258 30388
rect 15252 30348 36400 30376
rect 15252 30336 15258 30348
rect 1762 30308 1768 30320
rect 1723 30280 1768 30308
rect 1762 30268 1768 30280
rect 1820 30268 1826 30320
rect 2682 30308 2688 30320
rect 2643 30280 2688 30308
rect 2682 30268 2688 30280
rect 2740 30268 2746 30320
rect 36372 30308 36400 30348
rect 36446 30336 36452 30388
rect 36504 30376 36510 30388
rect 42426 30376 42432 30388
rect 36504 30348 42432 30376
rect 36504 30336 36510 30348
rect 42426 30336 42432 30348
rect 42484 30336 42490 30388
rect 37090 30308 37096 30320
rect 36372 30280 37096 30308
rect 37090 30268 37096 30280
rect 37148 30268 37154 30320
rect 48958 30200 48964 30252
rect 49016 30240 49022 30252
rect 49053 30243 49111 30249
rect 49053 30240 49065 30243
rect 49016 30212 49065 30240
rect 49016 30200 49022 30212
rect 49053 30209 49065 30212
rect 49099 30209 49111 30243
rect 49053 30203 49111 30209
rect 12066 30172 12072 30184
rect 12027 30144 12072 30172
rect 12066 30132 12072 30144
rect 12124 30132 12130 30184
rect 27614 30132 27620 30184
rect 27672 30172 27678 30184
rect 27801 30175 27859 30181
rect 27801 30172 27813 30175
rect 27672 30144 27813 30172
rect 27672 30132 27678 30144
rect 27801 30141 27813 30144
rect 27847 30141 27859 30175
rect 38930 30172 38936 30184
rect 38891 30144 38936 30172
rect 27801 30135 27859 30141
rect 38930 30132 38936 30144
rect 38988 30132 38994 30184
rect 48593 30175 48651 30181
rect 48593 30172 48605 30175
rect 45526 30144 48605 30172
rect 1949 30107 2007 30113
rect 1949 30073 1961 30107
rect 1995 30104 2007 30107
rect 2222 30104 2228 30116
rect 1995 30076 2228 30104
rect 1995 30073 2007 30076
rect 1949 30067 2007 30073
rect 2222 30064 2228 30076
rect 2280 30064 2286 30116
rect 17862 30064 17868 30116
rect 17920 30104 17926 30116
rect 32858 30104 32864 30116
rect 17920 30076 32864 30104
rect 17920 30064 17926 30076
rect 32858 30064 32864 30076
rect 32916 30064 32922 30116
rect 45526 30104 45554 30144
rect 48593 30141 48605 30144
rect 48639 30172 48651 30175
rect 49145 30175 49203 30181
rect 49145 30172 49157 30175
rect 48639 30144 49157 30172
rect 48639 30141 48651 30144
rect 48593 30135 48651 30141
rect 49145 30141 49157 30144
rect 49191 30141 49203 30175
rect 49145 30135 49203 30141
rect 41386 30076 45554 30104
rect 32398 29996 32404 30048
rect 32456 30036 32462 30048
rect 41386 30036 41414 30076
rect 32456 30008 41414 30036
rect 32456 29996 32462 30008
rect 1104 29946 68816 29968
rect 1104 29894 9246 29946
rect 9298 29894 9310 29946
rect 9362 29894 9374 29946
rect 9426 29894 9438 29946
rect 9490 29894 19246 29946
rect 19298 29894 19310 29946
rect 19362 29894 19374 29946
rect 19426 29894 19438 29946
rect 19490 29894 29246 29946
rect 29298 29894 29310 29946
rect 29362 29894 29374 29946
rect 29426 29894 29438 29946
rect 29490 29894 39246 29946
rect 39298 29894 39310 29946
rect 39362 29894 39374 29946
rect 39426 29894 39438 29946
rect 39490 29894 49246 29946
rect 49298 29894 49310 29946
rect 49362 29894 49374 29946
rect 49426 29894 49438 29946
rect 49490 29894 59246 29946
rect 59298 29894 59310 29946
rect 59362 29894 59374 29946
rect 59426 29894 59438 29946
rect 59490 29894 68816 29946
rect 1104 29872 68816 29894
rect 27065 29835 27123 29841
rect 27065 29801 27077 29835
rect 27111 29801 27123 29835
rect 27065 29795 27123 29801
rect 27157 29835 27215 29841
rect 27157 29801 27169 29835
rect 27203 29832 27215 29835
rect 28445 29835 28503 29841
rect 28445 29832 28457 29835
rect 27203 29804 28457 29832
rect 27203 29801 27215 29804
rect 27157 29795 27215 29801
rect 28445 29801 28457 29804
rect 28491 29832 28503 29835
rect 28534 29832 28540 29844
rect 28491 29804 28540 29832
rect 28491 29801 28503 29804
rect 28445 29795 28503 29801
rect 27080 29764 27108 29795
rect 28534 29792 28540 29804
rect 28592 29792 28598 29844
rect 27985 29767 28043 29773
rect 27985 29764 27997 29767
rect 27080 29736 27997 29764
rect 27985 29733 27997 29736
rect 28031 29764 28043 29767
rect 29546 29764 29552 29776
rect 28031 29736 29552 29764
rect 28031 29733 28043 29736
rect 27985 29727 28043 29733
rect 29546 29724 29552 29736
rect 29604 29764 29610 29776
rect 50706 29764 50712 29776
rect 29604 29736 50712 29764
rect 29604 29724 29610 29736
rect 50706 29724 50712 29736
rect 50764 29724 50770 29776
rect 2958 29656 2964 29708
rect 3016 29696 3022 29708
rect 26878 29696 26884 29708
rect 3016 29668 26884 29696
rect 3016 29656 3022 29668
rect 26878 29656 26884 29668
rect 26936 29656 26942 29708
rect 27249 29699 27307 29705
rect 27249 29665 27261 29699
rect 27295 29665 27307 29699
rect 27249 29659 27307 29665
rect 35897 29699 35955 29705
rect 35897 29665 35909 29699
rect 35943 29696 35955 29699
rect 54754 29696 54760 29708
rect 35943 29668 54760 29696
rect 35943 29665 35955 29668
rect 35897 29659 35955 29665
rect 27264 29628 27292 29659
rect 54754 29656 54760 29668
rect 54812 29656 54818 29708
rect 67453 29699 67511 29705
rect 67453 29665 67465 29699
rect 67499 29696 67511 29699
rect 68094 29696 68100 29708
rect 67499 29668 68100 29696
rect 67499 29665 67511 29668
rect 67453 29659 67511 29665
rect 68094 29656 68100 29668
rect 68152 29656 68158 29708
rect 26344 29600 27292 29628
rect 26344 29504 26372 29600
rect 28534 29588 28540 29640
rect 28592 29628 28598 29640
rect 50246 29628 50252 29640
rect 28592 29600 50252 29628
rect 28592 29588 28598 29600
rect 50246 29588 50252 29600
rect 50304 29588 50310 29640
rect 27433 29563 27491 29569
rect 27433 29529 27445 29563
rect 27479 29560 27491 29563
rect 53006 29560 53012 29572
rect 27479 29532 53012 29560
rect 27479 29529 27491 29532
rect 27433 29523 27491 29529
rect 53006 29520 53012 29532
rect 53064 29520 53070 29572
rect 2222 29492 2228 29504
rect 2183 29464 2228 29492
rect 2222 29452 2228 29464
rect 2280 29452 2286 29504
rect 7009 29495 7067 29501
rect 7009 29461 7021 29495
rect 7055 29492 7067 29495
rect 7374 29492 7380 29504
rect 7055 29464 7380 29492
rect 7055 29461 7067 29464
rect 7009 29455 7067 29461
rect 7374 29452 7380 29464
rect 7432 29452 7438 29504
rect 20990 29492 20996 29504
rect 20951 29464 20996 29492
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 26326 29492 26332 29504
rect 26287 29464 26332 29492
rect 26326 29452 26332 29464
rect 26384 29452 26390 29504
rect 1104 29402 68816 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 14246 29402
rect 14298 29350 14310 29402
rect 14362 29350 14374 29402
rect 14426 29350 14438 29402
rect 14490 29350 24246 29402
rect 24298 29350 24310 29402
rect 24362 29350 24374 29402
rect 24426 29350 24438 29402
rect 24490 29350 34246 29402
rect 34298 29350 34310 29402
rect 34362 29350 34374 29402
rect 34426 29350 34438 29402
rect 34490 29350 44246 29402
rect 44298 29350 44310 29402
rect 44362 29350 44374 29402
rect 44426 29350 44438 29402
rect 44490 29350 54246 29402
rect 54298 29350 54310 29402
rect 54362 29350 54374 29402
rect 54426 29350 54438 29402
rect 54490 29350 64246 29402
rect 64298 29350 64310 29402
rect 64362 29350 64374 29402
rect 64426 29350 64438 29402
rect 64490 29350 68816 29402
rect 1104 29328 68816 29350
rect 2222 29248 2228 29300
rect 2280 29288 2286 29300
rect 16666 29288 16672 29300
rect 2280 29260 16672 29288
rect 2280 29248 2286 29260
rect 16666 29248 16672 29260
rect 16724 29288 16730 29300
rect 17862 29288 17868 29300
rect 16724 29260 17868 29288
rect 16724 29248 16730 29260
rect 17862 29248 17868 29260
rect 17920 29248 17926 29300
rect 20990 29248 20996 29300
rect 21048 29288 21054 29300
rect 64046 29288 64052 29300
rect 21048 29260 64052 29288
rect 21048 29248 21054 29260
rect 64046 29248 64052 29260
rect 64104 29248 64110 29300
rect 26878 29180 26884 29232
rect 26936 29220 26942 29232
rect 27893 29223 27951 29229
rect 27893 29220 27905 29223
rect 26936 29192 27905 29220
rect 26936 29180 26942 29192
rect 27893 29189 27905 29192
rect 27939 29220 27951 29223
rect 34882 29220 34888 29232
rect 27939 29192 34888 29220
rect 27939 29189 27951 29192
rect 27893 29183 27951 29189
rect 34882 29180 34888 29192
rect 34940 29180 34946 29232
rect 22066 29124 31754 29152
rect 1762 29084 1768 29096
rect 1723 29056 1768 29084
rect 1762 29044 1768 29056
rect 1820 29044 1826 29096
rect 1949 29087 2007 29093
rect 1949 29053 1961 29087
rect 1995 29084 2007 29087
rect 2038 29084 2044 29096
rect 1995 29056 2044 29084
rect 1995 29053 2007 29056
rect 1949 29047 2007 29053
rect 2038 29044 2044 29056
rect 2096 29084 2102 29096
rect 2501 29087 2559 29093
rect 2501 29084 2513 29087
rect 2096 29056 2513 29084
rect 2096 29044 2102 29056
rect 2501 29053 2513 29056
rect 2547 29053 2559 29087
rect 2501 29047 2559 29053
rect 4798 29044 4804 29096
rect 4856 29084 4862 29096
rect 22066 29084 22094 29124
rect 4856 29056 22094 29084
rect 29089 29087 29147 29093
rect 4856 29044 4862 29056
rect 29089 29053 29101 29087
rect 29135 29053 29147 29087
rect 31726 29084 31754 29124
rect 59265 29087 59323 29093
rect 59265 29084 59277 29087
rect 31726 29056 59277 29084
rect 29089 29047 29147 29053
rect 59265 29053 59277 29056
rect 59311 29053 59323 29087
rect 59265 29047 59323 29053
rect 4982 28976 4988 29028
rect 5040 29016 5046 29028
rect 29104 29016 29132 29047
rect 5040 28988 29132 29016
rect 5040 28976 5046 28988
rect 1104 28858 68816 28880
rect 1104 28806 9246 28858
rect 9298 28806 9310 28858
rect 9362 28806 9374 28858
rect 9426 28806 9438 28858
rect 9490 28806 19246 28858
rect 19298 28806 19310 28858
rect 19362 28806 19374 28858
rect 19426 28806 19438 28858
rect 19490 28806 29246 28858
rect 29298 28806 29310 28858
rect 29362 28806 29374 28858
rect 29426 28806 29438 28858
rect 29490 28806 39246 28858
rect 39298 28806 39310 28858
rect 39362 28806 39374 28858
rect 39426 28806 39438 28858
rect 39490 28806 49246 28858
rect 49298 28806 49310 28858
rect 49362 28806 49374 28858
rect 49426 28806 49438 28858
rect 49490 28806 59246 28858
rect 59298 28806 59310 28858
rect 59362 28806 59374 28858
rect 59426 28806 59438 28858
rect 59490 28806 68816 28858
rect 1104 28784 68816 28806
rect 23014 28704 23020 28756
rect 23072 28744 23078 28756
rect 30929 28747 30987 28753
rect 30929 28744 30941 28747
rect 23072 28716 30941 28744
rect 23072 28704 23078 28716
rect 30929 28713 30941 28716
rect 30975 28744 30987 28747
rect 31478 28744 31484 28756
rect 30975 28716 31484 28744
rect 30975 28713 30987 28716
rect 30929 28707 30987 28713
rect 31478 28704 31484 28716
rect 31536 28704 31542 28756
rect 54941 28543 54999 28549
rect 54941 28509 54953 28543
rect 54987 28540 54999 28543
rect 66346 28540 66352 28552
rect 54987 28512 66352 28540
rect 54987 28509 54999 28512
rect 54941 28503 54999 28509
rect 66346 28500 66352 28512
rect 66404 28500 66410 28552
rect 31754 28364 31760 28416
rect 31812 28404 31818 28416
rect 38194 28404 38200 28416
rect 31812 28376 38200 28404
rect 31812 28364 31818 28376
rect 38194 28364 38200 28376
rect 38252 28364 38258 28416
rect 1104 28314 68816 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 14246 28314
rect 14298 28262 14310 28314
rect 14362 28262 14374 28314
rect 14426 28262 14438 28314
rect 14490 28262 24246 28314
rect 24298 28262 24310 28314
rect 24362 28262 24374 28314
rect 24426 28262 24438 28314
rect 24490 28262 34246 28314
rect 34298 28262 34310 28314
rect 34362 28262 34374 28314
rect 34426 28262 34438 28314
rect 34490 28262 44246 28314
rect 44298 28262 44310 28314
rect 44362 28262 44374 28314
rect 44426 28262 44438 28314
rect 44490 28262 54246 28314
rect 54298 28262 54310 28314
rect 54362 28262 54374 28314
rect 54426 28262 54438 28314
rect 54490 28262 64246 28314
rect 64298 28262 64310 28314
rect 64362 28262 64374 28314
rect 64426 28262 64438 28314
rect 64490 28262 68816 28314
rect 1104 28240 68816 28262
rect 13449 28203 13507 28209
rect 13449 28169 13461 28203
rect 13495 28200 13507 28203
rect 13538 28200 13544 28212
rect 13495 28172 13544 28200
rect 13495 28169 13507 28172
rect 13449 28163 13507 28169
rect 13538 28160 13544 28172
rect 13596 28160 13602 28212
rect 31481 28203 31539 28209
rect 31481 28169 31493 28203
rect 31527 28200 31539 28203
rect 31754 28200 31760 28212
rect 31527 28172 31760 28200
rect 31527 28169 31539 28172
rect 31481 28163 31539 28169
rect 31754 28160 31760 28172
rect 31812 28160 31818 28212
rect 32769 28203 32827 28209
rect 32769 28200 32781 28203
rect 31864 28172 32781 28200
rect 18693 28135 18751 28141
rect 18693 28101 18705 28135
rect 18739 28132 18751 28135
rect 31662 28132 31668 28144
rect 18739 28104 31668 28132
rect 18739 28101 18751 28104
rect 18693 28095 18751 28101
rect 31662 28092 31668 28104
rect 31720 28092 31726 28144
rect 2314 28024 2320 28076
rect 2372 28064 2378 28076
rect 17681 28067 17739 28073
rect 17681 28064 17693 28067
rect 2372 28036 17693 28064
rect 2372 28024 2378 28036
rect 17681 28033 17693 28036
rect 17727 28033 17739 28067
rect 17681 28027 17739 28033
rect 30926 28024 30932 28076
rect 30984 28064 30990 28076
rect 31021 28067 31079 28073
rect 31021 28064 31033 28067
rect 30984 28036 31033 28064
rect 30984 28024 30990 28036
rect 31021 28033 31033 28036
rect 31067 28064 31079 28067
rect 31386 28064 31392 28076
rect 31067 28036 31392 28064
rect 31067 28033 31079 28036
rect 31021 28027 31079 28033
rect 31386 28024 31392 28036
rect 31444 28064 31450 28076
rect 31757 28067 31815 28073
rect 31757 28064 31769 28067
rect 31444 28036 31769 28064
rect 31444 28024 31450 28036
rect 31757 28033 31769 28036
rect 31803 28033 31815 28067
rect 31864 28064 31892 28172
rect 32769 28169 32781 28172
rect 32815 28200 32827 28203
rect 33134 28200 33140 28212
rect 32815 28172 33140 28200
rect 32815 28169 32827 28172
rect 32769 28163 32827 28169
rect 33134 28160 33140 28172
rect 33192 28160 33198 28212
rect 32030 28092 32036 28144
rect 32088 28132 32094 28144
rect 46106 28132 46112 28144
rect 32088 28104 46112 28132
rect 32088 28092 32094 28104
rect 46106 28092 46112 28104
rect 46164 28092 46170 28144
rect 31864 28036 31984 28064
rect 31757 28027 31815 28033
rect 31478 27956 31484 28008
rect 31536 27996 31542 28008
rect 31956 28005 31984 28036
rect 31665 27999 31723 28005
rect 31665 27996 31677 27999
rect 31536 27968 31677 27996
rect 31536 27956 31542 27968
rect 31665 27965 31677 27968
rect 31711 27965 31723 27999
rect 31665 27959 31723 27965
rect 31849 27999 31907 28005
rect 31849 27965 31861 27999
rect 31895 27965 31907 27999
rect 31849 27959 31907 27965
rect 31941 27999 31999 28005
rect 31941 27965 31953 27999
rect 31987 27965 31999 27999
rect 31941 27959 31999 27965
rect 8478 27888 8484 27940
rect 8536 27928 8542 27940
rect 8536 27900 22094 27928
rect 8536 27888 8542 27900
rect 22066 27860 22094 27900
rect 31570 27888 31576 27940
rect 31628 27928 31634 27940
rect 31864 27928 31892 27959
rect 32030 27956 32036 28008
rect 32088 27996 32094 28008
rect 32125 27999 32183 28005
rect 32125 27996 32137 27999
rect 32088 27968 32137 27996
rect 32088 27956 32094 27968
rect 32125 27965 32137 27968
rect 32171 27965 32183 27999
rect 32125 27959 32183 27965
rect 35805 27999 35863 28005
rect 35805 27965 35817 27999
rect 35851 27965 35863 27999
rect 60458 27996 60464 28008
rect 60419 27968 60464 27996
rect 35805 27959 35863 27965
rect 35820 27928 35848 27959
rect 60458 27956 60464 27968
rect 60516 27956 60522 28008
rect 31628 27900 31892 27928
rect 32144 27900 35848 27928
rect 31628 27888 31634 27900
rect 32144 27860 32172 27900
rect 22066 27832 32172 27860
rect 32214 27820 32220 27872
rect 32272 27860 32278 27872
rect 33226 27860 33232 27872
rect 32272 27832 33232 27860
rect 32272 27820 32278 27832
rect 33226 27820 33232 27832
rect 33284 27820 33290 27872
rect 1104 27770 68816 27792
rect 1104 27718 9246 27770
rect 9298 27718 9310 27770
rect 9362 27718 9374 27770
rect 9426 27718 9438 27770
rect 9490 27718 19246 27770
rect 19298 27718 19310 27770
rect 19362 27718 19374 27770
rect 19426 27718 19438 27770
rect 19490 27718 29246 27770
rect 29298 27718 29310 27770
rect 29362 27718 29374 27770
rect 29426 27718 29438 27770
rect 29490 27718 39246 27770
rect 39298 27718 39310 27770
rect 39362 27718 39374 27770
rect 39426 27718 39438 27770
rect 39490 27718 49246 27770
rect 49298 27718 49310 27770
rect 49362 27718 49374 27770
rect 49426 27718 49438 27770
rect 49490 27718 59246 27770
rect 59298 27718 59310 27770
rect 59362 27718 59374 27770
rect 59426 27718 59438 27770
rect 59490 27718 68816 27770
rect 1104 27696 68816 27718
rect 30190 27616 30196 27668
rect 30248 27656 30254 27668
rect 33134 27656 33140 27668
rect 30248 27628 33140 27656
rect 30248 27616 30254 27628
rect 33134 27616 33140 27628
rect 33192 27616 33198 27668
rect 43622 27616 43628 27668
rect 43680 27656 43686 27668
rect 66162 27656 66168 27668
rect 43680 27628 66168 27656
rect 43680 27616 43686 27628
rect 66162 27616 66168 27628
rect 66220 27616 66226 27668
rect 47578 27548 47584 27600
rect 47636 27588 47642 27600
rect 48222 27588 48228 27600
rect 47636 27560 48228 27588
rect 47636 27548 47642 27560
rect 48222 27548 48228 27560
rect 48280 27548 48286 27600
rect 17793 27523 17851 27529
rect 17793 27489 17805 27523
rect 17839 27520 17851 27523
rect 18230 27520 18236 27532
rect 17839 27492 18236 27520
rect 17839 27489 17851 27492
rect 17793 27483 17851 27489
rect 18230 27480 18236 27492
rect 18288 27480 18294 27532
rect 18049 27455 18107 27461
rect 18049 27421 18061 27455
rect 18095 27452 18107 27455
rect 18782 27452 18788 27464
rect 18095 27424 18788 27452
rect 18095 27421 18107 27424
rect 18049 27415 18107 27421
rect 18782 27412 18788 27424
rect 18840 27412 18846 27464
rect 16666 27384 16672 27396
rect 16627 27356 16672 27384
rect 16666 27344 16672 27356
rect 16724 27344 16730 27396
rect 7190 27276 7196 27328
rect 7248 27316 7254 27328
rect 7653 27319 7711 27325
rect 7653 27316 7665 27319
rect 7248 27288 7665 27316
rect 7248 27276 7254 27288
rect 7653 27285 7665 27288
rect 7699 27285 7711 27319
rect 18506 27316 18512 27328
rect 18467 27288 18512 27316
rect 7653 27279 7711 27285
rect 18506 27276 18512 27288
rect 18564 27276 18570 27328
rect 31110 27316 31116 27328
rect 31071 27288 31116 27316
rect 31110 27276 31116 27288
rect 31168 27316 31174 27328
rect 31570 27316 31576 27328
rect 31168 27288 31576 27316
rect 31168 27276 31174 27288
rect 31570 27276 31576 27288
rect 31628 27276 31634 27328
rect 60918 27276 60924 27328
rect 60976 27316 60982 27328
rect 64969 27319 65027 27325
rect 64969 27316 64981 27319
rect 60976 27288 64981 27316
rect 60976 27276 60982 27288
rect 64969 27285 64981 27288
rect 65015 27285 65027 27319
rect 64969 27279 65027 27285
rect 1104 27226 68816 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 14246 27226
rect 14298 27174 14310 27226
rect 14362 27174 14374 27226
rect 14426 27174 14438 27226
rect 14490 27174 24246 27226
rect 24298 27174 24310 27226
rect 24362 27174 24374 27226
rect 24426 27174 24438 27226
rect 24490 27174 34246 27226
rect 34298 27174 34310 27226
rect 34362 27174 34374 27226
rect 34426 27174 34438 27226
rect 34490 27174 44246 27226
rect 44298 27174 44310 27226
rect 44362 27174 44374 27226
rect 44426 27174 44438 27226
rect 44490 27174 54246 27226
rect 54298 27174 54310 27226
rect 54362 27174 54374 27226
rect 54426 27174 54438 27226
rect 54490 27174 64246 27226
rect 64298 27174 64310 27226
rect 64362 27174 64374 27226
rect 64426 27174 64438 27226
rect 64490 27174 68816 27226
rect 1104 27152 68816 27174
rect 11054 27072 11060 27124
rect 11112 27112 11118 27124
rect 18782 27112 18788 27124
rect 11112 27084 18788 27112
rect 11112 27072 11118 27084
rect 18782 27072 18788 27084
rect 18840 27112 18846 27124
rect 25222 27112 25228 27124
rect 18840 27084 25228 27112
rect 18840 27072 18846 27084
rect 25222 27072 25228 27084
rect 25280 27112 25286 27124
rect 26142 27112 26148 27124
rect 25280 27084 26148 27112
rect 25280 27072 25286 27084
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 67266 27112 67272 27124
rect 67227 27084 67272 27112
rect 67266 27072 67272 27084
rect 67324 27072 67330 27124
rect 27338 27004 27344 27056
rect 27396 27044 27402 27056
rect 54570 27044 54576 27056
rect 27396 27016 54576 27044
rect 27396 27004 27402 27016
rect 54570 27004 54576 27016
rect 54628 27004 54634 27056
rect 32582 26936 32588 26988
rect 32640 26976 32646 26988
rect 32950 26976 32956 26988
rect 32640 26948 32956 26976
rect 32640 26936 32646 26948
rect 32950 26936 32956 26948
rect 33008 26976 33014 26988
rect 53834 26976 53840 26988
rect 33008 26948 53840 26976
rect 33008 26936 33014 26948
rect 53834 26936 53840 26948
rect 53892 26936 53898 26988
rect 68094 26976 68100 26988
rect 68055 26948 68100 26976
rect 68094 26936 68100 26948
rect 68152 26936 68158 26988
rect 1578 26908 1584 26920
rect 1539 26880 1584 26908
rect 1578 26868 1584 26880
rect 1636 26908 1642 26920
rect 2041 26911 2099 26917
rect 2041 26908 2053 26911
rect 1636 26880 2053 26908
rect 1636 26868 1642 26880
rect 2041 26877 2053 26880
rect 2087 26877 2099 26911
rect 2041 26871 2099 26877
rect 31389 26911 31447 26917
rect 31389 26877 31401 26911
rect 31435 26908 31447 26911
rect 67174 26908 67180 26920
rect 31435 26880 67180 26908
rect 31435 26877 31447 26880
rect 31389 26871 31447 26877
rect 67174 26868 67180 26880
rect 67232 26868 67238 26920
rect 67266 26868 67272 26920
rect 67324 26908 67330 26920
rect 67913 26911 67971 26917
rect 67913 26908 67925 26911
rect 67324 26880 67925 26908
rect 67324 26868 67330 26880
rect 67913 26877 67925 26880
rect 67959 26877 67971 26911
rect 67913 26871 67971 26877
rect 13998 26800 14004 26852
rect 14056 26840 14062 26852
rect 27890 26840 27896 26852
rect 14056 26812 27896 26840
rect 14056 26800 14062 26812
rect 27890 26800 27896 26812
rect 27948 26800 27954 26852
rect 47210 26800 47216 26852
rect 47268 26840 47274 26852
rect 57422 26840 57428 26852
rect 47268 26812 57428 26840
rect 47268 26800 47274 26812
rect 57422 26800 57428 26812
rect 57480 26800 57486 26852
rect 18230 26772 18236 26784
rect 18143 26744 18236 26772
rect 18230 26732 18236 26744
rect 18288 26772 18294 26784
rect 38378 26772 38384 26784
rect 18288 26744 38384 26772
rect 18288 26732 18294 26744
rect 38378 26732 38384 26744
rect 38436 26732 38442 26784
rect 1104 26682 68816 26704
rect 1104 26630 9246 26682
rect 9298 26630 9310 26682
rect 9362 26630 9374 26682
rect 9426 26630 9438 26682
rect 9490 26630 19246 26682
rect 19298 26630 19310 26682
rect 19362 26630 19374 26682
rect 19426 26630 19438 26682
rect 19490 26630 29246 26682
rect 29298 26630 29310 26682
rect 29362 26630 29374 26682
rect 29426 26630 29438 26682
rect 29490 26630 39246 26682
rect 39298 26630 39310 26682
rect 39362 26630 39374 26682
rect 39426 26630 39438 26682
rect 39490 26630 49246 26682
rect 49298 26630 49310 26682
rect 49362 26630 49374 26682
rect 49426 26630 49438 26682
rect 49490 26630 59246 26682
rect 59298 26630 59310 26682
rect 59362 26630 59374 26682
rect 59426 26630 59438 26682
rect 59490 26630 68816 26682
rect 1104 26608 68816 26630
rect 28166 26528 28172 26580
rect 28224 26568 28230 26580
rect 30190 26568 30196 26580
rect 28224 26540 30196 26568
rect 28224 26528 28230 26540
rect 30190 26528 30196 26540
rect 30248 26528 30254 26580
rect 33594 26528 33600 26580
rect 33652 26568 33658 26580
rect 42610 26568 42616 26580
rect 33652 26540 42616 26568
rect 33652 26528 33658 26540
rect 42610 26528 42616 26540
rect 42668 26568 42674 26580
rect 43073 26571 43131 26577
rect 43073 26568 43085 26571
rect 42668 26540 43085 26568
rect 42668 26528 42674 26540
rect 43073 26537 43085 26540
rect 43119 26537 43131 26571
rect 43073 26531 43131 26537
rect 47397 26571 47455 26577
rect 47397 26537 47409 26571
rect 47443 26568 47455 26571
rect 47486 26568 47492 26580
rect 47443 26540 47492 26568
rect 47443 26537 47455 26540
rect 47397 26531 47455 26537
rect 47486 26528 47492 26540
rect 47544 26568 47550 26580
rect 47544 26540 49832 26568
rect 47544 26528 47550 26540
rect 27890 26500 27896 26512
rect 27851 26472 27896 26500
rect 27890 26460 27896 26472
rect 27948 26460 27954 26512
rect 29549 26503 29607 26509
rect 29549 26500 29561 26503
rect 28000 26472 28304 26500
rect 24213 26435 24271 26441
rect 24213 26401 24225 26435
rect 24259 26432 24271 26435
rect 28000 26432 28028 26472
rect 28166 26432 28172 26444
rect 24259 26404 28028 26432
rect 28127 26404 28172 26432
rect 24259 26401 24271 26404
rect 24213 26395 24271 26401
rect 28166 26392 28172 26404
rect 28224 26392 28230 26444
rect 28276 26364 28304 26472
rect 29012 26472 29561 26500
rect 28442 26432 28448 26444
rect 28403 26404 28448 26432
rect 28442 26392 28448 26404
rect 28500 26392 28506 26444
rect 29012 26441 29040 26472
rect 29549 26469 29561 26472
rect 29595 26500 29607 26503
rect 32950 26500 32956 26512
rect 29595 26472 32956 26500
rect 29595 26469 29607 26472
rect 29549 26463 29607 26469
rect 32950 26460 32956 26472
rect 33008 26460 33014 26512
rect 47857 26503 47915 26509
rect 47857 26500 47869 26503
rect 33612 26472 47869 26500
rect 28997 26435 29055 26441
rect 28997 26401 29009 26435
rect 29043 26401 29055 26435
rect 30190 26432 30196 26444
rect 30151 26404 30196 26432
rect 28997 26395 29055 26401
rect 30190 26392 30196 26404
rect 30248 26392 30254 26444
rect 31386 26392 31392 26444
rect 31444 26432 31450 26444
rect 31662 26432 31668 26444
rect 31444 26404 31668 26432
rect 31444 26392 31450 26404
rect 31662 26392 31668 26404
rect 31720 26432 31726 26444
rect 33612 26432 33640 26472
rect 47857 26469 47869 26472
rect 47903 26500 47915 26503
rect 47903 26472 49464 26500
rect 47903 26469 47915 26472
rect 47857 26463 47915 26469
rect 31720 26404 33640 26432
rect 31720 26392 31726 26404
rect 37918 26392 37924 26444
rect 37976 26432 37982 26444
rect 38013 26435 38071 26441
rect 38013 26432 38025 26435
rect 37976 26404 38025 26432
rect 37976 26392 37982 26404
rect 38013 26401 38025 26404
rect 38059 26401 38071 26435
rect 38013 26395 38071 26401
rect 39942 26392 39948 26444
rect 40000 26432 40006 26444
rect 42521 26435 42579 26441
rect 42521 26432 42533 26435
rect 40000 26404 42533 26432
rect 40000 26392 40006 26404
rect 42521 26401 42533 26404
rect 42567 26401 42579 26435
rect 42521 26395 42579 26401
rect 42610 26392 42616 26444
rect 42668 26432 42674 26444
rect 42668 26404 42713 26432
rect 42668 26392 42674 26404
rect 48406 26392 48412 26444
rect 48464 26432 48470 26444
rect 48869 26435 48927 26441
rect 48869 26432 48881 26435
rect 48464 26404 48881 26432
rect 48464 26392 48470 26404
rect 48869 26401 48881 26404
rect 48915 26401 48927 26435
rect 48869 26395 48927 26401
rect 49237 26435 49295 26441
rect 49237 26401 49249 26435
rect 49283 26432 49295 26435
rect 49326 26432 49332 26444
rect 49283 26404 49332 26432
rect 49283 26401 49295 26404
rect 49237 26395 49295 26401
rect 49326 26392 49332 26404
rect 49384 26392 49390 26444
rect 49436 26441 49464 26472
rect 49421 26435 49479 26441
rect 49421 26401 49433 26435
rect 49467 26401 49479 26435
rect 49602 26432 49608 26444
rect 49563 26404 49608 26432
rect 49421 26395 49479 26401
rect 49602 26392 49608 26404
rect 49660 26392 49666 26444
rect 49804 26441 49832 26540
rect 49878 26528 49884 26580
rect 49936 26568 49942 26580
rect 50341 26571 50399 26577
rect 50341 26568 50353 26571
rect 49936 26540 50353 26568
rect 49936 26528 49942 26540
rect 50341 26537 50353 26540
rect 50387 26537 50399 26571
rect 50341 26531 50399 26537
rect 49789 26435 49847 26441
rect 49789 26401 49801 26435
rect 49835 26401 49847 26435
rect 49789 26395 49847 26401
rect 48498 26364 48504 26376
rect 6886 26336 28212 26364
rect 28276 26336 48360 26364
rect 48459 26336 48504 26364
rect 1765 26299 1823 26305
rect 1765 26265 1777 26299
rect 1811 26296 1823 26299
rect 6886 26296 6914 26336
rect 27338 26296 27344 26308
rect 1811 26268 6914 26296
rect 27299 26268 27344 26296
rect 1811 26265 1823 26268
rect 1765 26259 1823 26265
rect 27338 26256 27344 26268
rect 27396 26256 27402 26308
rect 28184 26296 28212 26336
rect 47210 26296 47216 26308
rect 28184 26268 47216 26296
rect 47210 26256 47216 26268
rect 47268 26256 47274 26308
rect 48332 26296 48360 26336
rect 48498 26324 48504 26336
rect 48556 26324 48562 26376
rect 48608 26336 55214 26364
rect 48608 26296 48636 26336
rect 48332 26268 48636 26296
rect 49418 26256 49424 26308
rect 49476 26296 49482 26308
rect 49878 26296 49884 26308
rect 49476 26268 49884 26296
rect 49476 26256 49482 26268
rect 49878 26256 49884 26268
rect 49936 26256 49942 26308
rect 55186 26296 55214 26336
rect 57238 26296 57244 26308
rect 55186 26268 57244 26296
rect 57238 26256 57244 26268
rect 57296 26256 57302 26308
rect 62666 26296 62672 26308
rect 62627 26268 62672 26296
rect 62666 26256 62672 26268
rect 62724 26256 62730 26308
rect 9582 26188 9588 26240
rect 9640 26228 9646 26240
rect 11054 26228 11060 26240
rect 9640 26200 11060 26228
rect 9640 26188 9646 26200
rect 11054 26188 11060 26200
rect 11112 26188 11118 26240
rect 47578 26188 47584 26240
rect 47636 26228 47642 26240
rect 49602 26228 49608 26240
rect 47636 26200 49608 26228
rect 47636 26188 47642 26200
rect 49602 26188 49608 26200
rect 49660 26188 49666 26240
rect 1104 26138 68816 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 14246 26138
rect 14298 26086 14310 26138
rect 14362 26086 14374 26138
rect 14426 26086 14438 26138
rect 14490 26086 24246 26138
rect 24298 26086 24310 26138
rect 24362 26086 24374 26138
rect 24426 26086 24438 26138
rect 24490 26086 34246 26138
rect 34298 26086 34310 26138
rect 34362 26086 34374 26138
rect 34426 26086 34438 26138
rect 34490 26086 44246 26138
rect 44298 26086 44310 26138
rect 44362 26086 44374 26138
rect 44426 26086 44438 26138
rect 44490 26086 54246 26138
rect 54298 26086 54310 26138
rect 54362 26086 54374 26138
rect 54426 26086 54438 26138
rect 54490 26086 64246 26138
rect 64298 26086 64310 26138
rect 64362 26086 64374 26138
rect 64426 26086 64438 26138
rect 64490 26086 68816 26138
rect 1104 26064 68816 26086
rect 27801 26027 27859 26033
rect 27801 25993 27813 26027
rect 27847 26024 27859 26027
rect 28442 26024 28448 26036
rect 27847 25996 28448 26024
rect 27847 25993 27859 25996
rect 27801 25987 27859 25993
rect 28442 25984 28448 25996
rect 28500 25984 28506 26036
rect 67361 26027 67419 26033
rect 67361 25993 67373 26027
rect 67407 26024 67419 26027
rect 67450 26024 67456 26036
rect 67407 25996 67456 26024
rect 67407 25993 67419 25996
rect 67361 25987 67419 25993
rect 67450 25984 67456 25996
rect 67508 25984 67514 26036
rect 2406 25916 2412 25968
rect 2464 25956 2470 25968
rect 55493 25959 55551 25965
rect 55493 25956 55505 25959
rect 2464 25928 55505 25956
rect 2464 25916 2470 25928
rect 55493 25925 55505 25928
rect 55539 25925 55551 25959
rect 55493 25919 55551 25925
rect 15286 25848 15292 25900
rect 15344 25888 15350 25900
rect 36722 25888 36728 25900
rect 15344 25860 36728 25888
rect 15344 25848 15350 25860
rect 36722 25848 36728 25860
rect 36780 25848 36786 25900
rect 13170 25780 13176 25832
rect 13228 25820 13234 25832
rect 58434 25820 58440 25832
rect 13228 25792 58440 25820
rect 13228 25780 13234 25792
rect 58434 25780 58440 25792
rect 58492 25780 58498 25832
rect 67450 25780 67456 25832
rect 67508 25820 67514 25832
rect 67913 25823 67971 25829
rect 67913 25820 67925 25823
rect 67508 25792 67925 25820
rect 67508 25780 67514 25792
rect 67913 25789 67925 25792
rect 67959 25789 67971 25823
rect 67913 25783 67971 25789
rect 17862 25712 17868 25764
rect 17920 25752 17926 25764
rect 42518 25752 42524 25764
rect 17920 25724 42524 25752
rect 17920 25712 17926 25724
rect 42518 25712 42524 25724
rect 42576 25712 42582 25764
rect 55769 25755 55827 25761
rect 55769 25721 55781 25755
rect 55815 25752 55827 25755
rect 56410 25752 56416 25764
rect 55815 25724 56416 25752
rect 55815 25721 55827 25724
rect 55769 25715 55827 25721
rect 56410 25712 56416 25724
rect 56468 25712 56474 25764
rect 68094 25752 68100 25764
rect 68055 25724 68100 25752
rect 68094 25712 68100 25724
rect 68152 25712 68158 25764
rect 47578 25644 47584 25696
rect 47636 25684 47642 25696
rect 47673 25687 47731 25693
rect 47673 25684 47685 25687
rect 47636 25656 47685 25684
rect 47636 25644 47642 25656
rect 47673 25653 47685 25656
rect 47719 25653 47731 25687
rect 48406 25684 48412 25696
rect 48367 25656 48412 25684
rect 47673 25647 47731 25653
rect 48406 25644 48412 25656
rect 48464 25644 48470 25696
rect 1104 25594 68816 25616
rect 1104 25542 9246 25594
rect 9298 25542 9310 25594
rect 9362 25542 9374 25594
rect 9426 25542 9438 25594
rect 9490 25542 19246 25594
rect 19298 25542 19310 25594
rect 19362 25542 19374 25594
rect 19426 25542 19438 25594
rect 19490 25542 29246 25594
rect 29298 25542 29310 25594
rect 29362 25542 29374 25594
rect 29426 25542 29438 25594
rect 29490 25542 39246 25594
rect 39298 25542 39310 25594
rect 39362 25542 39374 25594
rect 39426 25542 39438 25594
rect 39490 25542 49246 25594
rect 49298 25542 49310 25594
rect 49362 25542 49374 25594
rect 49426 25542 49438 25594
rect 49490 25542 59246 25594
rect 59298 25542 59310 25594
rect 59362 25542 59374 25594
rect 59426 25542 59438 25594
rect 59490 25542 68816 25594
rect 1104 25520 68816 25542
rect 11977 25483 12035 25489
rect 11977 25449 11989 25483
rect 12023 25480 12035 25483
rect 13170 25480 13176 25492
rect 12023 25452 13176 25480
rect 12023 25449 12035 25452
rect 11977 25443 12035 25449
rect 1949 25347 2007 25353
rect 1949 25313 1961 25347
rect 1995 25344 2007 25347
rect 11333 25347 11391 25353
rect 1995 25316 2636 25344
rect 1995 25313 2007 25316
rect 1949 25307 2007 25313
rect 1762 25208 1768 25220
rect 1723 25180 1768 25208
rect 1762 25168 1768 25180
rect 1820 25168 1826 25220
rect 2608 25152 2636 25316
rect 11333 25313 11345 25347
rect 11379 25344 11391 25347
rect 11992 25344 12020 25443
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 66165 25483 66223 25489
rect 66165 25449 66177 25483
rect 66211 25480 66223 25483
rect 66898 25480 66904 25492
rect 66211 25452 66904 25480
rect 66211 25449 66223 25452
rect 66165 25443 66223 25449
rect 66898 25440 66904 25452
rect 66956 25440 66962 25492
rect 11379 25316 12020 25344
rect 11379 25313 11391 25316
rect 11333 25307 11391 25313
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25276 11023 25279
rect 15286 25276 15292 25288
rect 11011 25248 15292 25276
rect 11011 25245 11023 25248
rect 10965 25239 11023 25245
rect 15286 25236 15292 25248
rect 15344 25236 15350 25288
rect 2590 25140 2596 25152
rect 2551 25112 2596 25140
rect 2590 25100 2596 25112
rect 2648 25100 2654 25152
rect 7926 25140 7932 25152
rect 7887 25112 7932 25140
rect 7926 25100 7932 25112
rect 7984 25100 7990 25152
rect 1104 25050 68816 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 14246 25050
rect 14298 24998 14310 25050
rect 14362 24998 14374 25050
rect 14426 24998 14438 25050
rect 14490 24998 24246 25050
rect 24298 24998 24310 25050
rect 24362 24998 24374 25050
rect 24426 24998 24438 25050
rect 24490 24998 34246 25050
rect 34298 24998 34310 25050
rect 34362 24998 34374 25050
rect 34426 24998 34438 25050
rect 34490 24998 44246 25050
rect 44298 24998 44310 25050
rect 44362 24998 44374 25050
rect 44426 24998 44438 25050
rect 44490 24998 54246 25050
rect 54298 24998 54310 25050
rect 54362 24998 54374 25050
rect 54426 24998 54438 25050
rect 54490 24998 64246 25050
rect 64298 24998 64310 25050
rect 64362 24998 64374 25050
rect 64426 24998 64438 25050
rect 64490 24998 68816 25050
rect 1104 24976 68816 24998
rect 2590 24896 2596 24948
rect 2648 24936 2654 24948
rect 16574 24936 16580 24948
rect 2648 24908 16580 24936
rect 2648 24896 2654 24908
rect 16574 24896 16580 24908
rect 16632 24936 16638 24948
rect 17862 24936 17868 24948
rect 16632 24908 17868 24936
rect 16632 24896 16638 24908
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 7926 24828 7932 24880
rect 7984 24868 7990 24880
rect 46474 24868 46480 24880
rect 7984 24840 46480 24868
rect 7984 24828 7990 24840
rect 46474 24828 46480 24840
rect 46532 24828 46538 24880
rect 23474 24760 23480 24812
rect 23532 24800 23538 24812
rect 58526 24800 58532 24812
rect 23532 24772 58532 24800
rect 23532 24760 23538 24772
rect 58526 24760 58532 24772
rect 58584 24760 58590 24812
rect 36906 24732 36912 24744
rect 36867 24704 36912 24732
rect 36906 24692 36912 24704
rect 36964 24692 36970 24744
rect 63494 24692 63500 24744
rect 63552 24732 63558 24744
rect 64509 24735 64567 24741
rect 64509 24732 64521 24735
rect 63552 24704 64521 24732
rect 63552 24692 63558 24704
rect 64509 24701 64521 24704
rect 64555 24701 64567 24735
rect 64509 24695 64567 24701
rect 67453 24735 67511 24741
rect 67453 24701 67465 24735
rect 67499 24732 67511 24735
rect 68094 24732 68100 24744
rect 67499 24704 68100 24732
rect 67499 24701 67511 24704
rect 67453 24695 67511 24701
rect 68094 24692 68100 24704
rect 68152 24692 68158 24744
rect 1104 24506 68816 24528
rect 1104 24454 9246 24506
rect 9298 24454 9310 24506
rect 9362 24454 9374 24506
rect 9426 24454 9438 24506
rect 9490 24454 19246 24506
rect 19298 24454 19310 24506
rect 19362 24454 19374 24506
rect 19426 24454 19438 24506
rect 19490 24454 29246 24506
rect 29298 24454 29310 24506
rect 29362 24454 29374 24506
rect 29426 24454 29438 24506
rect 29490 24454 39246 24506
rect 39298 24454 39310 24506
rect 39362 24454 39374 24506
rect 39426 24454 39438 24506
rect 39490 24454 49246 24506
rect 49298 24454 49310 24506
rect 49362 24454 49374 24506
rect 49426 24454 49438 24506
rect 49490 24454 59246 24506
rect 59298 24454 59310 24506
rect 59362 24454 59374 24506
rect 59426 24454 59438 24506
rect 59490 24454 68816 24506
rect 1104 24432 68816 24454
rect 23474 24392 23480 24404
rect 22848 24364 23480 24392
rect 19978 24216 19984 24268
rect 20036 24256 20042 24268
rect 20622 24256 20628 24268
rect 20036 24228 20628 24256
rect 20036 24216 20042 24228
rect 20622 24216 20628 24228
rect 20680 24256 20686 24268
rect 22848 24265 22876 24364
rect 23474 24352 23480 24364
rect 23532 24352 23538 24404
rect 21913 24259 21971 24265
rect 21913 24256 21925 24259
rect 20680 24228 21925 24256
rect 20680 24216 20686 24228
rect 21913 24225 21925 24228
rect 21959 24225 21971 24259
rect 21913 24219 21971 24225
rect 22833 24259 22891 24265
rect 22833 24225 22845 24259
rect 22879 24225 22891 24259
rect 22833 24219 22891 24225
rect 33689 24259 33747 24265
rect 33689 24225 33701 24259
rect 33735 24256 33747 24259
rect 36538 24256 36544 24268
rect 33735 24228 36544 24256
rect 33735 24225 33747 24228
rect 33689 24219 33747 24225
rect 36538 24216 36544 24228
rect 36596 24216 36602 24268
rect 1854 24148 1860 24200
rect 1912 24188 1918 24200
rect 67913 24191 67971 24197
rect 67913 24188 67925 24191
rect 1912 24160 67925 24188
rect 1912 24148 1918 24160
rect 67913 24157 67925 24160
rect 67959 24157 67971 24191
rect 67913 24151 67971 24157
rect 7466 24080 7472 24132
rect 7524 24120 7530 24132
rect 54754 24120 54760 24132
rect 7524 24092 54760 24120
rect 7524 24080 7530 24092
rect 54754 24080 54760 24092
rect 54812 24080 54818 24132
rect 12342 24052 12348 24064
rect 12303 24024 12348 24052
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 29086 24052 29092 24064
rect 29047 24024 29092 24052
rect 29086 24012 29092 24024
rect 29144 24012 29150 24064
rect 54110 24052 54116 24064
rect 54071 24024 54116 24052
rect 54110 24012 54116 24024
rect 54168 24012 54174 24064
rect 1104 23962 68816 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 14246 23962
rect 14298 23910 14310 23962
rect 14362 23910 14374 23962
rect 14426 23910 14438 23962
rect 14490 23910 24246 23962
rect 24298 23910 24310 23962
rect 24362 23910 24374 23962
rect 24426 23910 24438 23962
rect 24490 23910 34246 23962
rect 34298 23910 34310 23962
rect 34362 23910 34374 23962
rect 34426 23910 34438 23962
rect 34490 23910 44246 23962
rect 44298 23910 44310 23962
rect 44362 23910 44374 23962
rect 44426 23910 44438 23962
rect 44490 23910 54246 23962
rect 54298 23910 54310 23962
rect 54362 23910 54374 23962
rect 54426 23910 54438 23962
rect 54490 23910 64246 23962
rect 64298 23910 64310 23962
rect 64362 23910 64374 23962
rect 64426 23910 64438 23962
rect 64490 23910 68816 23962
rect 1104 23888 68816 23910
rect 1854 23848 1860 23860
rect 1815 23820 1860 23848
rect 1854 23808 1860 23820
rect 1912 23808 1918 23860
rect 2593 23851 2651 23857
rect 2593 23817 2605 23851
rect 2639 23848 2651 23851
rect 3142 23848 3148 23860
rect 2639 23820 3148 23848
rect 2639 23817 2651 23820
rect 2593 23811 2651 23817
rect 1949 23647 2007 23653
rect 1949 23613 1961 23647
rect 1995 23644 2007 23647
rect 2608 23644 2636 23811
rect 3142 23808 3148 23820
rect 3200 23808 3206 23860
rect 5442 23808 5448 23860
rect 5500 23848 5506 23860
rect 54110 23848 54116 23860
rect 5500 23820 54116 23848
rect 5500 23808 5506 23820
rect 54110 23808 54116 23820
rect 54168 23808 54174 23860
rect 29086 23740 29092 23792
rect 29144 23780 29150 23792
rect 66714 23780 66720 23792
rect 29144 23752 66720 23780
rect 29144 23740 29150 23752
rect 66714 23740 66720 23752
rect 66772 23740 66778 23792
rect 12342 23672 12348 23724
rect 12400 23712 12406 23724
rect 37734 23712 37740 23724
rect 12400 23684 37740 23712
rect 12400 23672 12406 23684
rect 37734 23672 37740 23684
rect 37792 23672 37798 23724
rect 57333 23715 57391 23721
rect 57333 23712 57345 23715
rect 45526 23684 57345 23712
rect 45526 23644 45554 23684
rect 57333 23681 57345 23684
rect 57379 23681 57391 23715
rect 57333 23675 57391 23681
rect 1995 23616 2636 23644
rect 6886 23616 45554 23644
rect 1995 23613 2007 23616
rect 1949 23607 2007 23613
rect 2314 23536 2320 23588
rect 2372 23576 2378 23588
rect 6886 23576 6914 23616
rect 47578 23604 47584 23656
rect 47636 23644 47642 23656
rect 53009 23647 53067 23653
rect 53009 23644 53021 23647
rect 47636 23616 53021 23644
rect 47636 23604 47642 23616
rect 53009 23613 53021 23616
rect 53055 23644 53067 23647
rect 54297 23647 54355 23653
rect 54297 23644 54309 23647
rect 53055 23616 54309 23644
rect 53055 23613 53067 23616
rect 53009 23607 53067 23613
rect 54297 23613 54309 23616
rect 54343 23613 54355 23647
rect 54297 23607 54355 23613
rect 54386 23604 54392 23656
rect 54444 23644 54450 23656
rect 54573 23647 54631 23653
rect 54444 23616 54489 23644
rect 54444 23604 54450 23616
rect 54573 23613 54585 23647
rect 54619 23613 54631 23647
rect 54573 23607 54631 23613
rect 2372 23548 6914 23576
rect 2372 23536 2378 23548
rect 36630 23536 36636 23588
rect 36688 23576 36694 23588
rect 53834 23576 53840 23588
rect 36688 23548 53144 23576
rect 53795 23548 53840 23576
rect 36688 23536 36694 23548
rect 53116 23508 53144 23548
rect 53834 23536 53840 23548
rect 53892 23576 53898 23588
rect 54588 23576 54616 23607
rect 53892 23548 54616 23576
rect 53892 23536 53898 23548
rect 53926 23508 53932 23520
rect 53116 23480 53932 23508
rect 53926 23468 53932 23480
rect 53984 23508 53990 23520
rect 54386 23508 54392 23520
rect 53984 23480 54392 23508
rect 53984 23468 53990 23480
rect 54386 23468 54392 23480
rect 54444 23468 54450 23520
rect 54754 23508 54760 23520
rect 54715 23480 54760 23508
rect 54754 23468 54760 23480
rect 54812 23468 54818 23520
rect 56413 23511 56471 23517
rect 56413 23477 56425 23511
rect 56459 23508 56471 23511
rect 56502 23508 56508 23520
rect 56459 23480 56508 23508
rect 56459 23477 56471 23480
rect 56413 23471 56471 23477
rect 56502 23468 56508 23480
rect 56560 23468 56566 23520
rect 1104 23418 68816 23440
rect 1104 23366 9246 23418
rect 9298 23366 9310 23418
rect 9362 23366 9374 23418
rect 9426 23366 9438 23418
rect 9490 23366 19246 23418
rect 19298 23366 19310 23418
rect 19362 23366 19374 23418
rect 19426 23366 19438 23418
rect 19490 23366 29246 23418
rect 29298 23366 29310 23418
rect 29362 23366 29374 23418
rect 29426 23366 29438 23418
rect 29490 23366 39246 23418
rect 39298 23366 39310 23418
rect 39362 23366 39374 23418
rect 39426 23366 39438 23418
rect 39490 23366 49246 23418
rect 49298 23366 49310 23418
rect 49362 23366 49374 23418
rect 49426 23366 49438 23418
rect 49490 23366 59246 23418
rect 59298 23366 59310 23418
rect 59362 23366 59374 23418
rect 59426 23366 59438 23418
rect 59490 23366 68816 23418
rect 1104 23344 68816 23366
rect 13170 23264 13176 23316
rect 13228 23304 13234 23316
rect 58434 23304 58440 23316
rect 13228 23276 58296 23304
rect 58395 23276 58440 23304
rect 13228 23264 13234 23276
rect 9214 23196 9220 23248
rect 9272 23236 9278 23248
rect 37550 23236 37556 23248
rect 9272 23208 37556 23236
rect 9272 23196 9278 23208
rect 37550 23196 37556 23208
rect 37608 23196 37614 23248
rect 53926 23236 53932 23248
rect 53887 23208 53932 23236
rect 53926 23196 53932 23208
rect 53984 23196 53990 23248
rect 55769 23239 55827 23245
rect 55769 23236 55781 23239
rect 55186 23208 55781 23236
rect 22922 23128 22928 23180
rect 22980 23168 22986 23180
rect 39666 23168 39672 23180
rect 22980 23140 39672 23168
rect 22980 23128 22986 23140
rect 39666 23128 39672 23140
rect 39724 23128 39730 23180
rect 50062 23128 50068 23180
rect 50120 23168 50126 23180
rect 55186 23168 55214 23208
rect 55769 23205 55781 23208
rect 55815 23236 55827 23239
rect 58268 23236 58296 23276
rect 58434 23264 58440 23276
rect 58492 23264 58498 23316
rect 67358 23304 67364 23316
rect 67319 23276 67364 23304
rect 67358 23264 67364 23276
rect 67416 23304 67422 23316
rect 67416 23276 67956 23304
rect 67416 23264 67422 23276
rect 62390 23236 62396 23248
rect 55815 23208 57454 23236
rect 58268 23208 62396 23236
rect 55815 23205 55827 23208
rect 55769 23199 55827 23205
rect 62390 23196 62396 23208
rect 62448 23196 62454 23248
rect 67928 23245 67956 23276
rect 67913 23239 67971 23245
rect 67913 23205 67925 23239
rect 67959 23205 67971 23239
rect 67913 23199 67971 23205
rect 50120 23140 55214 23168
rect 50120 23128 50126 23140
rect 30098 23060 30104 23112
rect 30156 23100 30162 23112
rect 33686 23100 33692 23112
rect 30156 23072 33692 23100
rect 30156 23060 30162 23072
rect 33686 23060 33692 23072
rect 33744 23060 33750 23112
rect 56502 23060 56508 23112
rect 56560 23100 56566 23112
rect 56689 23103 56747 23109
rect 56689 23100 56701 23103
rect 56560 23072 56701 23100
rect 56560 23060 56566 23072
rect 56689 23069 56701 23072
rect 56735 23069 56747 23103
rect 56962 23100 56968 23112
rect 56923 23072 56968 23100
rect 56689 23063 56747 23069
rect 56962 23060 56968 23072
rect 57020 23060 57026 23112
rect 54110 23032 54116 23044
rect 22066 23004 54116 23032
rect 11701 22967 11759 22973
rect 11701 22933 11713 22967
rect 11747 22964 11759 22967
rect 22066 22964 22094 23004
rect 54110 22992 54116 23004
rect 54168 22992 54174 23044
rect 68094 23032 68100 23044
rect 68055 23004 68100 23032
rect 68094 22992 68100 23004
rect 68152 22992 68158 23044
rect 11747 22936 22094 22964
rect 11747 22933 11759 22936
rect 11701 22927 11759 22933
rect 29914 22924 29920 22976
rect 29972 22964 29978 22976
rect 33594 22964 33600 22976
rect 29972 22936 33600 22964
rect 29972 22924 29978 22936
rect 33594 22924 33600 22936
rect 33652 22924 33658 22976
rect 37918 22964 37924 22976
rect 37879 22936 37924 22964
rect 37918 22924 37924 22936
rect 37976 22924 37982 22976
rect 38194 22924 38200 22976
rect 38252 22964 38258 22976
rect 38654 22964 38660 22976
rect 38252 22936 38660 22964
rect 38252 22924 38258 22936
rect 38654 22924 38660 22936
rect 38712 22924 38718 22976
rect 1104 22874 68816 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 14246 22874
rect 14298 22822 14310 22874
rect 14362 22822 14374 22874
rect 14426 22822 14438 22874
rect 14490 22822 24246 22874
rect 24298 22822 24310 22874
rect 24362 22822 24374 22874
rect 24426 22822 24438 22874
rect 24490 22822 34246 22874
rect 34298 22822 34310 22874
rect 34362 22822 34374 22874
rect 34426 22822 34438 22874
rect 34490 22822 44246 22874
rect 44298 22822 44310 22874
rect 44362 22822 44374 22874
rect 44426 22822 44438 22874
rect 44490 22822 54246 22874
rect 54298 22822 54310 22874
rect 54362 22822 54374 22874
rect 54426 22822 54438 22874
rect 54490 22822 64246 22874
rect 64298 22822 64310 22874
rect 64362 22822 64374 22874
rect 64426 22822 64438 22874
rect 64490 22822 68816 22874
rect 1104 22800 68816 22822
rect 3694 22720 3700 22772
rect 3752 22760 3758 22772
rect 30469 22763 30527 22769
rect 30469 22760 30481 22763
rect 3752 22732 30481 22760
rect 3752 22720 3758 22732
rect 30469 22729 30481 22732
rect 30515 22729 30527 22763
rect 31570 22760 31576 22772
rect 30469 22723 30527 22729
rect 30576 22732 31576 22760
rect 9214 22692 9220 22704
rect 9175 22664 9220 22692
rect 9214 22652 9220 22664
rect 9272 22652 9278 22704
rect 13170 22692 13176 22704
rect 13131 22664 13176 22692
rect 13170 22652 13176 22664
rect 13228 22652 13234 22704
rect 29914 22692 29920 22704
rect 29875 22664 29920 22692
rect 29914 22652 29920 22664
rect 29972 22652 29978 22704
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22624 7343 22627
rect 9232 22624 9260 22652
rect 7331 22596 9260 22624
rect 7331 22593 7343 22596
rect 7285 22587 7343 22593
rect 26142 22584 26148 22636
rect 26200 22624 26206 22636
rect 30576 22624 30604 22732
rect 31570 22720 31576 22732
rect 31628 22720 31634 22772
rect 34974 22720 34980 22772
rect 35032 22760 35038 22772
rect 38562 22760 38568 22772
rect 35032 22732 38568 22760
rect 35032 22720 35038 22732
rect 38562 22720 38568 22732
rect 38620 22720 38626 22772
rect 39666 22760 39672 22772
rect 39627 22732 39672 22760
rect 39666 22720 39672 22732
rect 39724 22720 39730 22772
rect 62025 22763 62083 22769
rect 62025 22729 62037 22763
rect 62071 22760 62083 22763
rect 64598 22760 64604 22772
rect 62071 22732 64604 22760
rect 62071 22729 62083 22732
rect 62025 22723 62083 22729
rect 64598 22720 64604 22732
rect 64656 22720 64662 22772
rect 26200 22596 30604 22624
rect 31036 22664 31708 22692
rect 26200 22584 26206 22596
rect 31036 22565 31064 22664
rect 7009 22559 7067 22565
rect 7009 22525 7021 22559
rect 7055 22556 7067 22559
rect 30648 22559 30706 22565
rect 7055 22528 9812 22556
rect 7055 22525 7067 22528
rect 7009 22519 7067 22525
rect 8570 22420 8576 22432
rect 8531 22392 8576 22420
rect 8570 22380 8576 22392
rect 8628 22380 8634 22432
rect 9784 22429 9812 22528
rect 30648 22525 30660 22559
rect 30694 22556 30706 22559
rect 31021 22559 31079 22565
rect 30694 22528 30972 22556
rect 30694 22525 30706 22528
rect 30648 22519 30706 22525
rect 30098 22448 30104 22500
rect 30156 22488 30162 22500
rect 30745 22491 30803 22497
rect 30745 22488 30757 22491
rect 30156 22460 30757 22488
rect 30156 22448 30162 22460
rect 30745 22457 30757 22460
rect 30791 22457 30803 22491
rect 30745 22451 30803 22457
rect 30837 22491 30895 22497
rect 30837 22457 30849 22491
rect 30883 22457 30895 22491
rect 30944 22488 30972 22528
rect 31021 22525 31033 22559
rect 31067 22525 31079 22559
rect 31680 22556 31708 22664
rect 56502 22624 56508 22636
rect 38304 22596 56508 22624
rect 32033 22559 32091 22565
rect 32033 22556 32045 22559
rect 31680 22528 32045 22556
rect 31021 22519 31079 22525
rect 32033 22525 32045 22528
rect 32079 22556 32091 22559
rect 38194 22556 38200 22568
rect 32079 22528 38200 22556
rect 32079 22525 32091 22528
rect 32033 22519 32091 22525
rect 38194 22516 38200 22528
rect 38252 22516 38258 22568
rect 38304 22565 38332 22596
rect 56502 22584 56508 22596
rect 56560 22584 56566 22636
rect 38289 22559 38347 22565
rect 38289 22525 38301 22559
rect 38335 22525 38347 22559
rect 38565 22559 38623 22565
rect 38565 22556 38577 22559
rect 38289 22519 38347 22525
rect 38396 22528 38577 22556
rect 31481 22491 31539 22497
rect 31481 22488 31493 22491
rect 30944 22460 31493 22488
rect 30837 22451 30895 22457
rect 31481 22457 31493 22460
rect 31527 22457 31539 22491
rect 31481 22451 31539 22457
rect 9769 22423 9827 22429
rect 9769 22389 9781 22423
rect 9815 22420 9827 22423
rect 11054 22420 11060 22432
rect 9815 22392 11060 22420
rect 9815 22389 9827 22392
rect 9769 22383 9827 22389
rect 11054 22380 11060 22392
rect 11112 22420 11118 22432
rect 11882 22420 11888 22432
rect 11112 22392 11888 22420
rect 11112 22380 11118 22392
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 29914 22380 29920 22432
rect 29972 22420 29978 22432
rect 30852 22420 30880 22451
rect 29972 22392 30880 22420
rect 31496 22420 31524 22451
rect 31570 22448 31576 22500
rect 31628 22488 31634 22500
rect 37918 22488 37924 22500
rect 31628 22460 37924 22488
rect 31628 22448 31634 22460
rect 37918 22448 37924 22460
rect 37976 22488 37982 22500
rect 38304 22488 38332 22519
rect 37976 22460 38332 22488
rect 37976 22448 37982 22460
rect 37642 22420 37648 22432
rect 31496 22392 37648 22420
rect 29972 22380 29978 22392
rect 37642 22380 37648 22392
rect 37700 22380 37706 22432
rect 37826 22380 37832 22432
rect 37884 22420 37890 22432
rect 38396 22420 38424 22528
rect 38565 22525 38577 22528
rect 38611 22525 38623 22559
rect 46382 22556 46388 22568
rect 46343 22528 46388 22556
rect 38565 22519 38623 22525
rect 46382 22516 46388 22528
rect 46440 22516 46446 22568
rect 37884 22392 38424 22420
rect 37884 22380 37890 22392
rect 38562 22380 38568 22432
rect 38620 22420 38626 22432
rect 56597 22423 56655 22429
rect 56597 22420 56609 22423
rect 38620 22392 56609 22420
rect 38620 22380 38626 22392
rect 56597 22389 56609 22392
rect 56643 22420 56655 22423
rect 56962 22420 56968 22432
rect 56643 22392 56968 22420
rect 56643 22389 56655 22392
rect 56597 22383 56655 22389
rect 56962 22380 56968 22392
rect 57020 22380 57026 22432
rect 1104 22330 68816 22352
rect 1104 22278 9246 22330
rect 9298 22278 9310 22330
rect 9362 22278 9374 22330
rect 9426 22278 9438 22330
rect 9490 22278 19246 22330
rect 19298 22278 19310 22330
rect 19362 22278 19374 22330
rect 19426 22278 19438 22330
rect 19490 22278 29246 22330
rect 29298 22278 29310 22330
rect 29362 22278 29374 22330
rect 29426 22278 29438 22330
rect 29490 22278 39246 22330
rect 39298 22278 39310 22330
rect 39362 22278 39374 22330
rect 39426 22278 39438 22330
rect 39490 22278 49246 22330
rect 49298 22278 49310 22330
rect 49362 22278 49374 22330
rect 49426 22278 49438 22330
rect 49490 22278 59246 22330
rect 59298 22278 59310 22330
rect 59362 22278 59374 22330
rect 59426 22278 59438 22330
rect 59490 22278 68816 22330
rect 1104 22256 68816 22278
rect 8570 22176 8576 22228
rect 8628 22216 8634 22228
rect 30098 22216 30104 22228
rect 8628 22188 30104 22216
rect 8628 22176 8634 22188
rect 30098 22176 30104 22188
rect 30156 22176 30162 22228
rect 37826 22176 37832 22228
rect 37884 22216 37890 22228
rect 38105 22219 38163 22225
rect 38105 22216 38117 22219
rect 37884 22188 38117 22216
rect 37884 22176 37890 22188
rect 38105 22185 38117 22188
rect 38151 22185 38163 22219
rect 38105 22179 38163 22185
rect 11790 22040 11796 22092
rect 11848 22080 11854 22092
rect 18874 22080 18880 22092
rect 11848 22052 18880 22080
rect 11848 22040 11854 22052
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 15289 21879 15347 21885
rect 15289 21845 15301 21879
rect 15335 21876 15347 21879
rect 22094 21876 22100 21888
rect 15335 21848 22100 21876
rect 15335 21845 15347 21848
rect 15289 21839 15347 21845
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 1104 21786 68816 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 14246 21786
rect 14298 21734 14310 21786
rect 14362 21734 14374 21786
rect 14426 21734 14438 21786
rect 14490 21734 24246 21786
rect 24298 21734 24310 21786
rect 24362 21734 24374 21786
rect 24426 21734 24438 21786
rect 24490 21734 34246 21786
rect 34298 21734 34310 21786
rect 34362 21734 34374 21786
rect 34426 21734 34438 21786
rect 34490 21734 44246 21786
rect 44298 21734 44310 21786
rect 44362 21734 44374 21786
rect 44426 21734 44438 21786
rect 44490 21734 54246 21786
rect 54298 21734 54310 21786
rect 54362 21734 54374 21786
rect 54426 21734 54438 21786
rect 54490 21734 64246 21786
rect 64298 21734 64310 21786
rect 64362 21734 64374 21786
rect 64426 21734 64438 21786
rect 64490 21734 68816 21786
rect 1104 21712 68816 21734
rect 67266 21672 67272 21684
rect 67227 21644 67272 21672
rect 67266 21632 67272 21644
rect 67324 21632 67330 21684
rect 15010 21564 15016 21616
rect 15068 21604 15074 21616
rect 36906 21604 36912 21616
rect 15068 21576 36912 21604
rect 15068 21564 15074 21576
rect 36906 21564 36912 21576
rect 36964 21564 36970 21616
rect 38746 21564 38752 21616
rect 38804 21604 38810 21616
rect 56226 21604 56232 21616
rect 38804 21576 56232 21604
rect 38804 21564 38810 21576
rect 56226 21564 56232 21576
rect 56284 21564 56290 21616
rect 68094 21604 68100 21616
rect 68055 21576 68100 21604
rect 68094 21564 68100 21576
rect 68152 21564 68158 21616
rect 23934 21496 23940 21548
rect 23992 21536 23998 21548
rect 62666 21536 62672 21548
rect 23992 21508 62672 21536
rect 23992 21496 23998 21508
rect 62666 21496 62672 21508
rect 62724 21496 62730 21548
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 2409 21471 2467 21477
rect 2409 21437 2421 21471
rect 2455 21468 2467 21471
rect 11974 21468 11980 21480
rect 2455 21440 11980 21468
rect 2455 21437 2467 21440
rect 2409 21431 2467 21437
rect 11974 21428 11980 21440
rect 12032 21428 12038 21480
rect 13081 21471 13139 21477
rect 13081 21437 13093 21471
rect 13127 21468 13139 21471
rect 25590 21468 25596 21480
rect 13127 21440 25596 21468
rect 13127 21437 13139 21440
rect 13081 21431 13139 21437
rect 25590 21428 25596 21440
rect 25648 21428 25654 21480
rect 31481 21471 31539 21477
rect 31481 21437 31493 21471
rect 31527 21437 31539 21471
rect 31481 21431 31539 21437
rect 33597 21471 33655 21477
rect 33597 21437 33609 21471
rect 33643 21468 33655 21471
rect 36081 21471 36139 21477
rect 33643 21440 35894 21468
rect 33643 21437 33655 21440
rect 33597 21431 33655 21437
rect 31496 21332 31524 21431
rect 35866 21400 35894 21440
rect 36081 21437 36093 21471
rect 36127 21468 36139 21471
rect 39758 21468 39764 21480
rect 36127 21440 39764 21468
rect 36127 21437 36139 21440
rect 36081 21431 36139 21437
rect 39758 21428 39764 21440
rect 39816 21428 39822 21480
rect 67266 21428 67272 21480
rect 67324 21468 67330 21480
rect 67913 21471 67971 21477
rect 67913 21468 67925 21471
rect 67324 21440 67925 21468
rect 67324 21428 67330 21440
rect 67913 21437 67925 21440
rect 67959 21437 67971 21471
rect 67913 21431 67971 21437
rect 39850 21400 39856 21412
rect 35866 21372 39856 21400
rect 39850 21360 39856 21372
rect 39908 21360 39914 21412
rect 55398 21360 55404 21412
rect 55456 21400 55462 21412
rect 67082 21400 67088 21412
rect 55456 21372 67088 21400
rect 55456 21360 55462 21372
rect 67082 21360 67088 21372
rect 67140 21360 67146 21412
rect 47854 21332 47860 21344
rect 31496 21304 47860 21332
rect 47854 21292 47860 21304
rect 47912 21292 47918 21344
rect 1104 21242 68816 21264
rect 1104 21190 9246 21242
rect 9298 21190 9310 21242
rect 9362 21190 9374 21242
rect 9426 21190 9438 21242
rect 9490 21190 19246 21242
rect 19298 21190 19310 21242
rect 19362 21190 19374 21242
rect 19426 21190 19438 21242
rect 19490 21190 29246 21242
rect 29298 21190 29310 21242
rect 29362 21190 29374 21242
rect 29426 21190 29438 21242
rect 29490 21190 39246 21242
rect 39298 21190 39310 21242
rect 39362 21190 39374 21242
rect 39426 21190 39438 21242
rect 39490 21190 49246 21242
rect 49298 21190 49310 21242
rect 49362 21190 49374 21242
rect 49426 21190 49438 21242
rect 49490 21190 59246 21242
rect 59298 21190 59310 21242
rect 59362 21190 59374 21242
rect 59426 21190 59438 21242
rect 59490 21190 68816 21242
rect 1104 21168 68816 21190
rect 1394 21128 1400 21140
rect 1355 21100 1400 21128
rect 1394 21088 1400 21100
rect 1452 21088 1458 21140
rect 57974 20952 57980 21004
rect 58032 20992 58038 21004
rect 60918 20992 60924 21004
rect 58032 20964 60924 20992
rect 58032 20952 58038 20964
rect 60918 20952 60924 20964
rect 60976 20952 60982 21004
rect 33137 20859 33195 20865
rect 33137 20825 33149 20859
rect 33183 20856 33195 20859
rect 52546 20856 52552 20868
rect 33183 20828 52552 20856
rect 33183 20825 33195 20828
rect 33137 20819 33195 20825
rect 52546 20816 52552 20828
rect 52604 20816 52610 20868
rect 37277 20791 37335 20797
rect 37277 20757 37289 20791
rect 37323 20788 37335 20791
rect 38838 20788 38844 20800
rect 37323 20760 38844 20788
rect 37323 20757 37335 20760
rect 37277 20751 37335 20757
rect 38838 20748 38844 20760
rect 38896 20748 38902 20800
rect 1104 20698 68816 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 14246 20698
rect 14298 20646 14310 20698
rect 14362 20646 14374 20698
rect 14426 20646 14438 20698
rect 14490 20646 24246 20698
rect 24298 20646 24310 20698
rect 24362 20646 24374 20698
rect 24426 20646 24438 20698
rect 24490 20646 34246 20698
rect 34298 20646 34310 20698
rect 34362 20646 34374 20698
rect 34426 20646 34438 20698
rect 34490 20646 44246 20698
rect 44298 20646 44310 20698
rect 44362 20646 44374 20698
rect 44426 20646 44438 20698
rect 44490 20646 54246 20698
rect 54298 20646 54310 20698
rect 54362 20646 54374 20698
rect 54426 20646 54438 20698
rect 54490 20646 64246 20698
rect 64298 20646 64310 20698
rect 64362 20646 64374 20698
rect 64426 20646 64438 20698
rect 64490 20646 68816 20698
rect 1104 20624 68816 20646
rect 27798 20584 27804 20596
rect 27759 20556 27804 20584
rect 27798 20544 27804 20556
rect 27856 20544 27862 20596
rect 28445 20587 28503 20593
rect 28445 20553 28457 20587
rect 28491 20584 28503 20587
rect 31110 20584 31116 20596
rect 28491 20556 31116 20584
rect 28491 20553 28503 20556
rect 28445 20547 28503 20553
rect 31110 20544 31116 20556
rect 31168 20544 31174 20596
rect 28994 20340 29000 20392
rect 29052 20380 29058 20392
rect 29273 20383 29331 20389
rect 29273 20380 29285 20383
rect 29052 20352 29285 20380
rect 29052 20340 29058 20352
rect 29273 20349 29285 20352
rect 29319 20349 29331 20383
rect 29273 20343 29331 20349
rect 30285 20383 30343 20389
rect 30285 20349 30297 20383
rect 30331 20380 30343 20383
rect 67082 20380 67088 20392
rect 30331 20352 67088 20380
rect 30331 20349 30343 20352
rect 30285 20343 30343 20349
rect 67082 20340 67088 20352
rect 67140 20340 67146 20392
rect 67453 20383 67511 20389
rect 67453 20349 67465 20383
rect 67499 20380 67511 20383
rect 68094 20380 68100 20392
rect 67499 20352 68100 20380
rect 67499 20349 67511 20352
rect 67453 20343 67511 20349
rect 68094 20340 68100 20352
rect 68152 20340 68158 20392
rect 1104 20154 68816 20176
rect 1104 20102 9246 20154
rect 9298 20102 9310 20154
rect 9362 20102 9374 20154
rect 9426 20102 9438 20154
rect 9490 20102 19246 20154
rect 19298 20102 19310 20154
rect 19362 20102 19374 20154
rect 19426 20102 19438 20154
rect 19490 20102 29246 20154
rect 29298 20102 29310 20154
rect 29362 20102 29374 20154
rect 29426 20102 29438 20154
rect 29490 20102 39246 20154
rect 39298 20102 39310 20154
rect 39362 20102 39374 20154
rect 39426 20102 39438 20154
rect 39490 20102 49246 20154
rect 49298 20102 49310 20154
rect 49362 20102 49374 20154
rect 49426 20102 49438 20154
rect 49490 20102 59246 20154
rect 59298 20102 59310 20154
rect 59362 20102 59374 20154
rect 59426 20102 59438 20154
rect 59490 20102 68816 20154
rect 1104 20080 68816 20102
rect 1854 20040 1860 20052
rect 1815 20012 1860 20040
rect 1854 20000 1860 20012
rect 1912 20000 1918 20052
rect 27246 20040 27252 20052
rect 27207 20012 27252 20040
rect 27246 20000 27252 20012
rect 27304 20000 27310 20052
rect 30009 20043 30067 20049
rect 30009 20009 30021 20043
rect 30055 20040 30067 20043
rect 30098 20040 30104 20052
rect 30055 20012 30104 20040
rect 30055 20009 30067 20012
rect 30009 20003 30067 20009
rect 1949 19907 2007 19913
rect 1949 19873 1961 19907
rect 1995 19904 2007 19907
rect 2593 19907 2651 19913
rect 2593 19904 2605 19907
rect 1995 19876 2605 19904
rect 1995 19873 2007 19876
rect 1949 19867 2007 19873
rect 2593 19873 2605 19876
rect 2639 19904 2651 19907
rect 14826 19904 14832 19916
rect 2639 19876 14832 19904
rect 2639 19873 2651 19876
rect 2593 19867 2651 19873
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 27264 19904 27292 20000
rect 30024 19972 30052 20003
rect 30098 20000 30104 20012
rect 30156 20000 30162 20052
rect 29288 19944 30052 19972
rect 29288 19913 29316 19944
rect 32398 19932 32404 19984
rect 32456 19972 32462 19984
rect 50062 19972 50068 19984
rect 32456 19944 50068 19972
rect 32456 19932 32462 19944
rect 50062 19932 50068 19944
rect 50120 19932 50126 19984
rect 28997 19907 29055 19913
rect 28997 19904 29009 19907
rect 27264 19876 29009 19904
rect 28997 19873 29009 19876
rect 29043 19873 29055 19907
rect 28997 19867 29055 19873
rect 29273 19907 29331 19913
rect 29273 19873 29285 19907
rect 29319 19873 29331 19907
rect 29273 19867 29331 19873
rect 29457 19907 29515 19913
rect 29457 19873 29469 19907
rect 29503 19873 29515 19907
rect 29457 19867 29515 19873
rect 30929 19907 30987 19913
rect 30929 19873 30941 19907
rect 30975 19904 30987 19907
rect 31846 19904 31852 19916
rect 30975 19876 31852 19904
rect 30975 19873 30987 19876
rect 30929 19867 30987 19873
rect 27798 19796 27804 19848
rect 27856 19836 27862 19848
rect 29472 19836 29500 19867
rect 31846 19864 31852 19876
rect 31904 19864 31910 19916
rect 27856 19808 29500 19836
rect 31665 19839 31723 19845
rect 27856 19796 27862 19808
rect 31665 19805 31677 19839
rect 31711 19836 31723 19839
rect 36630 19836 36636 19848
rect 31711 19808 36636 19836
rect 31711 19805 31723 19808
rect 31665 19799 31723 19805
rect 36630 19796 36636 19808
rect 36688 19796 36694 19848
rect 28813 19771 28871 19777
rect 28813 19768 28825 19771
rect 6886 19740 28825 19768
rect 5074 19660 5080 19712
rect 5132 19700 5138 19712
rect 6886 19700 6914 19740
rect 28813 19737 28825 19740
rect 28859 19737 28871 19771
rect 28813 19731 28871 19737
rect 29089 19771 29147 19777
rect 29089 19737 29101 19771
rect 29135 19737 29147 19771
rect 29089 19731 29147 19737
rect 29181 19771 29239 19777
rect 29181 19737 29193 19771
rect 29227 19768 29239 19771
rect 31110 19768 31116 19780
rect 29227 19740 31116 19768
rect 29227 19737 29239 19740
rect 29181 19731 29239 19737
rect 28258 19700 28264 19712
rect 5132 19672 6914 19700
rect 28171 19672 28264 19700
rect 5132 19660 5138 19672
rect 28258 19660 28264 19672
rect 28316 19700 28322 19712
rect 29104 19700 29132 19731
rect 31110 19728 31116 19740
rect 31168 19728 31174 19780
rect 31662 19700 31668 19712
rect 28316 19672 31668 19700
rect 28316 19660 28322 19672
rect 31662 19660 31668 19672
rect 31720 19660 31726 19712
rect 33962 19700 33968 19712
rect 33923 19672 33968 19700
rect 33962 19660 33968 19672
rect 34020 19660 34026 19712
rect 50338 19660 50344 19712
rect 50396 19700 50402 19712
rect 50433 19703 50491 19709
rect 50433 19700 50445 19703
rect 50396 19672 50445 19700
rect 50396 19660 50402 19672
rect 50433 19669 50445 19672
rect 50479 19669 50491 19703
rect 53282 19700 53288 19712
rect 53243 19672 53288 19700
rect 50433 19663 50491 19669
rect 53282 19660 53288 19672
rect 53340 19660 53346 19712
rect 1104 19610 68816 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 14246 19610
rect 14298 19558 14310 19610
rect 14362 19558 14374 19610
rect 14426 19558 14438 19610
rect 14490 19558 24246 19610
rect 24298 19558 24310 19610
rect 24362 19558 24374 19610
rect 24426 19558 24438 19610
rect 24490 19558 34246 19610
rect 34298 19558 34310 19610
rect 34362 19558 34374 19610
rect 34426 19558 34438 19610
rect 34490 19558 44246 19610
rect 44298 19558 44310 19610
rect 44362 19558 44374 19610
rect 44426 19558 44438 19610
rect 44490 19558 54246 19610
rect 54298 19558 54310 19610
rect 54362 19558 54374 19610
rect 54426 19558 54438 19610
rect 54490 19558 64246 19610
rect 64298 19558 64310 19610
rect 64362 19558 64374 19610
rect 64426 19558 64438 19610
rect 64490 19558 68816 19610
rect 1104 19536 68816 19558
rect 18230 19456 18236 19508
rect 18288 19496 18294 19508
rect 28258 19496 28264 19508
rect 18288 19468 28264 19496
rect 18288 19456 18294 19468
rect 28258 19456 28264 19468
rect 28316 19456 28322 19508
rect 49697 19363 49755 19369
rect 49697 19329 49709 19363
rect 49743 19360 49755 19363
rect 61654 19360 61660 19372
rect 49743 19332 61660 19360
rect 49743 19329 49755 19332
rect 49697 19323 49755 19329
rect 61654 19320 61660 19332
rect 61712 19320 61718 19372
rect 67913 19227 67971 19233
rect 67913 19224 67925 19227
rect 67284 19196 67925 19224
rect 41322 19116 41328 19168
rect 41380 19156 41386 19168
rect 67284 19165 67312 19196
rect 67913 19193 67925 19196
rect 67959 19193 67971 19227
rect 68094 19224 68100 19236
rect 68055 19196 68100 19224
rect 67913 19187 67971 19193
rect 68094 19184 68100 19196
rect 68152 19184 68158 19236
rect 67269 19159 67327 19165
rect 67269 19156 67281 19159
rect 41380 19128 67281 19156
rect 41380 19116 41386 19128
rect 67269 19125 67281 19128
rect 67315 19125 67327 19159
rect 67269 19119 67327 19125
rect 1104 19066 18952 19088
rect 1104 19014 9246 19066
rect 9298 19014 9310 19066
rect 9362 19014 9374 19066
rect 9426 19014 9438 19066
rect 9490 19014 18952 19066
rect 1104 18992 18952 19014
rect 37628 19066 68816 19088
rect 37628 19014 39246 19066
rect 39298 19014 39310 19066
rect 39362 19014 39374 19066
rect 39426 19014 39438 19066
rect 39490 19014 49246 19066
rect 49298 19014 49310 19066
rect 49362 19014 49374 19066
rect 49426 19014 49438 19066
rect 49490 19014 59246 19066
rect 59298 19014 59310 19066
rect 59362 19014 59374 19066
rect 59426 19014 59438 19066
rect 59490 19014 68816 19066
rect 37628 18992 68816 19014
rect 2222 18912 2228 18964
rect 2280 18952 2286 18964
rect 2501 18955 2559 18961
rect 2501 18952 2513 18955
rect 2280 18924 2513 18952
rect 2280 18912 2286 18924
rect 2501 18921 2513 18924
rect 2547 18921 2559 18955
rect 2501 18915 2559 18921
rect 15102 18912 15108 18964
rect 15160 18952 15166 18964
rect 26326 18952 26332 18964
rect 15160 18924 26332 18952
rect 15160 18912 15166 18924
rect 26326 18912 26332 18924
rect 26384 18912 26390 18964
rect 33226 18912 33232 18964
rect 33284 18952 33290 18964
rect 50522 18952 50528 18964
rect 33284 18924 50528 18952
rect 33284 18912 33290 18924
rect 50522 18912 50528 18924
rect 50580 18912 50586 18964
rect 1949 18887 2007 18893
rect 1949 18853 1961 18887
rect 1995 18884 2007 18887
rect 2240 18884 2268 18912
rect 1995 18856 2268 18884
rect 1995 18853 2007 18856
rect 1949 18847 2007 18853
rect 16390 18844 16396 18896
rect 16448 18884 16454 18896
rect 33962 18884 33968 18896
rect 16448 18856 33968 18884
rect 16448 18844 16454 18856
rect 33962 18844 33968 18856
rect 34020 18844 34026 18896
rect 13906 18776 13912 18828
rect 13964 18816 13970 18828
rect 38930 18816 38936 18828
rect 13964 18788 38936 18816
rect 13964 18776 13970 18788
rect 38930 18776 38936 18788
rect 38988 18776 38994 18828
rect 50798 18776 50804 18828
rect 50856 18816 50862 18828
rect 51261 18819 51319 18825
rect 51261 18816 51273 18819
rect 50856 18788 51273 18816
rect 50856 18776 50862 18788
rect 51261 18785 51273 18788
rect 51307 18785 51319 18819
rect 51261 18779 51319 18785
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 45002 18748 45008 18760
rect 18380 18720 45008 18748
rect 18380 18708 18386 18720
rect 45002 18708 45008 18720
rect 45060 18708 45066 18760
rect 1762 18680 1768 18692
rect 1723 18652 1768 18680
rect 1762 18640 1768 18652
rect 1820 18640 1826 18692
rect 2866 18640 2872 18692
rect 2924 18680 2930 18692
rect 66070 18680 66076 18692
rect 2924 18652 66076 18680
rect 2924 18640 2930 18652
rect 66070 18640 66076 18652
rect 66128 18640 66134 18692
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 9493 18615 9551 18621
rect 9493 18612 9505 18615
rect 8444 18584 9505 18612
rect 8444 18572 8450 18584
rect 9493 18581 9505 18584
rect 9539 18581 9551 18615
rect 9493 18575 9551 18581
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 48406 18612 48412 18624
rect 15804 18584 48412 18612
rect 15804 18572 15810 18584
rect 48406 18572 48412 18584
rect 48464 18572 48470 18624
rect 1104 18522 18952 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 14246 18522
rect 14298 18470 14310 18522
rect 14362 18470 14374 18522
rect 14426 18470 14438 18522
rect 14490 18470 18952 18522
rect 1104 18448 18952 18470
rect 37628 18522 68816 18544
rect 37628 18470 44246 18522
rect 44298 18470 44310 18522
rect 44362 18470 44374 18522
rect 44426 18470 44438 18522
rect 44490 18470 54246 18522
rect 54298 18470 54310 18522
rect 54362 18470 54374 18522
rect 54426 18470 54438 18522
rect 54490 18470 64246 18522
rect 64298 18470 64310 18522
rect 64362 18470 64374 18522
rect 64426 18470 64438 18522
rect 64490 18470 68816 18522
rect 37628 18448 68816 18470
rect 18230 18408 18236 18420
rect 18191 18380 18236 18408
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 61470 18408 61476 18420
rect 61431 18380 61476 18408
rect 61470 18368 61476 18380
rect 61528 18368 61534 18420
rect 17681 18139 17739 18145
rect 17681 18105 17693 18139
rect 17727 18136 17739 18139
rect 17862 18136 17868 18148
rect 17727 18108 17868 18136
rect 17727 18105 17739 18108
rect 17681 18099 17739 18105
rect 17862 18096 17868 18108
rect 17920 18136 17926 18148
rect 34606 18136 34612 18148
rect 17920 18108 34612 18136
rect 17920 18096 17926 18108
rect 34606 18096 34612 18108
rect 34664 18096 34670 18148
rect 1104 17978 18952 18000
rect 1104 17926 9246 17978
rect 9298 17926 9310 17978
rect 9362 17926 9374 17978
rect 9426 17926 9438 17978
rect 9490 17926 18952 17978
rect 1104 17904 18952 17926
rect 37628 17978 68816 18000
rect 37628 17926 39246 17978
rect 39298 17926 39310 17978
rect 39362 17926 39374 17978
rect 39426 17926 39438 17978
rect 39490 17926 49246 17978
rect 49298 17926 49310 17978
rect 49362 17926 49374 17978
rect 49426 17926 49438 17978
rect 49490 17926 59246 17978
rect 59298 17926 59310 17978
rect 59362 17926 59374 17978
rect 59426 17926 59438 17978
rect 59490 17926 68816 17978
rect 37628 17904 68816 17926
rect 17770 17864 17776 17876
rect 17731 17836 17776 17864
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 66622 17824 66628 17876
rect 66680 17864 66686 17876
rect 67269 17867 67327 17873
rect 67269 17864 67281 17867
rect 66680 17836 67281 17864
rect 66680 17824 66686 17836
rect 67269 17833 67281 17836
rect 67315 17864 67327 17867
rect 67315 17836 67956 17864
rect 67315 17833 67327 17836
rect 67269 17827 67327 17833
rect 18230 17796 18236 17808
rect 17512 17768 18236 17796
rect 17512 17737 17540 17768
rect 18230 17756 18236 17768
rect 18288 17756 18294 17808
rect 67928 17805 67956 17836
rect 67913 17799 67971 17805
rect 67913 17765 67925 17799
rect 67959 17765 67971 17799
rect 67913 17759 67971 17765
rect 17497 17731 17555 17737
rect 17497 17697 17509 17731
rect 17543 17697 17555 17731
rect 17862 17728 17868 17740
rect 17823 17700 17868 17728
rect 17497 17691 17555 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 68094 17728 68100 17740
rect 68055 17700 68100 17728
rect 68094 17688 68100 17700
rect 68152 17688 68158 17740
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 28994 17660 29000 17672
rect 17276 17632 29000 17660
rect 17276 17620 17282 17632
rect 28994 17620 29000 17632
rect 29052 17620 29058 17672
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 48498 17592 48504 17604
rect 11204 17564 48504 17592
rect 11204 17552 11210 17564
rect 48498 17552 48504 17564
rect 48556 17552 48562 17604
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 36998 17524 37004 17536
rect 18196 17496 37004 17524
rect 18196 17484 18202 17496
rect 36998 17484 37004 17496
rect 37056 17484 37062 17536
rect 47673 17527 47731 17533
rect 47673 17493 47685 17527
rect 47719 17524 47731 17527
rect 56042 17524 56048 17536
rect 47719 17496 56048 17524
rect 47719 17493 47731 17496
rect 47673 17487 47731 17493
rect 56042 17484 56048 17496
rect 56100 17484 56106 17536
rect 1104 17434 18952 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 14246 17434
rect 14298 17382 14310 17434
rect 14362 17382 14374 17434
rect 14426 17382 14438 17434
rect 14490 17382 18952 17434
rect 1104 17360 18952 17382
rect 37628 17434 68816 17456
rect 37628 17382 44246 17434
rect 44298 17382 44310 17434
rect 44362 17382 44374 17434
rect 44426 17382 44438 17434
rect 44490 17382 54246 17434
rect 54298 17382 54310 17434
rect 54362 17382 54374 17434
rect 54426 17382 54438 17434
rect 54490 17382 64246 17434
rect 64298 17382 64310 17434
rect 64362 17382 64374 17434
rect 64426 17382 64438 17434
rect 64490 17382 68816 17434
rect 37628 17360 68816 17382
rect 15838 17280 15844 17332
rect 15896 17320 15902 17332
rect 65794 17320 65800 17332
rect 15896 17292 65800 17320
rect 15896 17280 15902 17292
rect 65794 17280 65800 17292
rect 65852 17280 65858 17332
rect 10226 17212 10232 17264
rect 10284 17252 10290 17264
rect 63494 17252 63500 17264
rect 10284 17224 63500 17252
rect 10284 17212 10290 17224
rect 63494 17212 63500 17224
rect 63552 17212 63558 17264
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 18233 17119 18291 17125
rect 10091 17088 16574 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 16546 16980 16574 17088
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18279 17088 26234 17116
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 26206 17048 26234 17088
rect 53926 17076 53932 17128
rect 53984 17116 53990 17128
rect 55769 17119 55827 17125
rect 55769 17116 55781 17119
rect 53984 17088 55781 17116
rect 53984 17076 53990 17088
rect 55769 17085 55781 17088
rect 55815 17085 55827 17119
rect 55769 17079 55827 17085
rect 61565 17119 61623 17125
rect 61565 17085 61577 17119
rect 61611 17085 61623 17119
rect 61565 17079 61623 17085
rect 42518 17048 42524 17060
rect 26206 17020 42524 17048
rect 42518 17008 42524 17020
rect 42576 17008 42582 17060
rect 54938 17008 54944 17060
rect 54996 17048 55002 17060
rect 61580 17048 61608 17079
rect 54996 17020 61608 17048
rect 54996 17008 55002 17020
rect 63862 16980 63868 16992
rect 16546 16952 63868 16980
rect 63862 16940 63868 16952
rect 63920 16940 63926 16992
rect 1104 16890 18952 16912
rect 1104 16838 9246 16890
rect 9298 16838 9310 16890
rect 9362 16838 9374 16890
rect 9426 16838 9438 16890
rect 9490 16838 18952 16890
rect 1104 16816 18952 16838
rect 37628 16890 68816 16912
rect 37628 16838 39246 16890
rect 39298 16838 39310 16890
rect 39362 16838 39374 16890
rect 39426 16838 39438 16890
rect 39490 16838 49246 16890
rect 49298 16838 49310 16890
rect 49362 16838 49374 16890
rect 49426 16838 49438 16890
rect 49490 16838 59246 16890
rect 59298 16838 59310 16890
rect 59362 16838 59374 16890
rect 59426 16838 59438 16890
rect 59490 16838 68816 16890
rect 37628 16816 68816 16838
rect 50706 16668 50712 16720
rect 50764 16708 50770 16720
rect 50764 16680 56732 16708
rect 50764 16668 50770 16680
rect 56134 16600 56140 16652
rect 56192 16640 56198 16652
rect 56704 16649 56732 16680
rect 56505 16643 56563 16649
rect 56505 16640 56517 16643
rect 56192 16612 56517 16640
rect 56192 16600 56198 16612
rect 56505 16609 56517 16612
rect 56551 16609 56563 16643
rect 56505 16603 56563 16609
rect 56689 16643 56747 16649
rect 56689 16609 56701 16643
rect 56735 16640 56747 16643
rect 57149 16643 57207 16649
rect 57149 16640 57161 16643
rect 56735 16612 57161 16640
rect 56735 16609 56747 16612
rect 56689 16603 56747 16609
rect 57149 16609 57161 16612
rect 57195 16609 57207 16643
rect 57149 16603 57207 16609
rect 67453 16643 67511 16649
rect 67453 16609 67465 16643
rect 67499 16640 67511 16643
rect 68094 16640 68100 16652
rect 67499 16612 68100 16640
rect 67499 16609 67511 16612
rect 67453 16603 67511 16609
rect 68094 16600 68100 16612
rect 68152 16600 68158 16652
rect 27614 16572 27620 16584
rect 27575 16544 27620 16572
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 56502 16504 56508 16516
rect 56463 16476 56508 16504
rect 56502 16464 56508 16476
rect 56560 16464 56566 16516
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16436 18291 16439
rect 63494 16436 63500 16448
rect 18279 16408 63500 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 63494 16396 63500 16408
rect 63552 16396 63558 16448
rect 1104 16346 18952 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 14246 16346
rect 14298 16294 14310 16346
rect 14362 16294 14374 16346
rect 14426 16294 14438 16346
rect 14490 16294 18952 16346
rect 1104 16272 18952 16294
rect 37628 16346 68816 16368
rect 37628 16294 44246 16346
rect 44298 16294 44310 16346
rect 44362 16294 44374 16346
rect 44426 16294 44438 16346
rect 44490 16294 54246 16346
rect 54298 16294 54310 16346
rect 54362 16294 54374 16346
rect 54426 16294 54438 16346
rect 54490 16294 64246 16346
rect 64298 16294 64310 16346
rect 64362 16294 64374 16346
rect 64426 16294 64438 16346
rect 64490 16294 68816 16346
rect 37628 16272 68816 16294
rect 18046 16232 18052 16244
rect 18007 16204 18052 16232
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 56134 16232 56140 16244
rect 56095 16204 56140 16232
rect 56134 16192 56140 16204
rect 56192 16192 56198 16244
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 16028 1642 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1636 16000 2053 16028
rect 1636 15988 1642 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 16028 7067 16031
rect 66990 16028 66996 16040
rect 7055 16000 66996 16028
rect 7055 15997 7067 16000
rect 7009 15991 7067 15997
rect 66990 15988 66996 16000
rect 67048 15988 67054 16040
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 27617 15895 27675 15901
rect 27617 15892 27629 15895
rect 17368 15864 27629 15892
rect 17368 15852 17374 15864
rect 27617 15861 27629 15864
rect 27663 15861 27675 15895
rect 27617 15855 27675 15861
rect 32582 15852 32588 15904
rect 32640 15892 32646 15904
rect 47578 15892 47584 15904
rect 32640 15864 47584 15892
rect 32640 15852 32646 15864
rect 47578 15852 47584 15864
rect 47636 15852 47642 15904
rect 50614 15852 50620 15904
rect 50672 15892 50678 15904
rect 56134 15892 56140 15904
rect 50672 15864 56140 15892
rect 50672 15852 50678 15864
rect 56134 15852 56140 15864
rect 56192 15852 56198 15904
rect 1104 15802 18952 15824
rect 1104 15750 9246 15802
rect 9298 15750 9310 15802
rect 9362 15750 9374 15802
rect 9426 15750 9438 15802
rect 9490 15750 18952 15802
rect 1104 15728 18952 15750
rect 37628 15802 68816 15824
rect 37628 15750 39246 15802
rect 39298 15750 39310 15802
rect 39362 15750 39374 15802
rect 39426 15750 39438 15802
rect 39490 15750 49246 15802
rect 49298 15750 49310 15802
rect 49362 15750 49374 15802
rect 49426 15750 49438 15802
rect 49490 15750 59246 15802
rect 59298 15750 59310 15802
rect 59362 15750 59374 15802
rect 59426 15750 59438 15802
rect 59490 15750 68816 15802
rect 37628 15728 68816 15750
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 11296 15660 11345 15688
rect 11296 15648 11302 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 67726 15688 67732 15700
rect 67687 15660 67732 15688
rect 11333 15651 11391 15657
rect 67726 15648 67732 15660
rect 67784 15648 67790 15700
rect 2130 15512 2136 15564
rect 2188 15552 2194 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 2188 15524 5917 15552
rect 2188 15512 2194 15524
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15552 10563 15555
rect 10778 15552 10784 15564
rect 10551 15524 10784 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 10778 15512 10784 15524
rect 10836 15552 10842 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 10836 15524 11437 15552
rect 10836 15512 10842 15524
rect 11425 15521 11437 15524
rect 11471 15552 11483 15555
rect 17402 15552 17408 15564
rect 11471 15524 17408 15552
rect 11471 15521 11483 15524
rect 11425 15515 11483 15521
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 11882 15308 11888 15360
rect 11940 15348 11946 15360
rect 12250 15348 12256 15360
rect 11940 15320 12256 15348
rect 11940 15308 11946 15320
rect 12250 15308 12256 15320
rect 12308 15348 12314 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 12308 15320 17693 15348
rect 12308 15308 12314 15320
rect 17681 15317 17693 15320
rect 17727 15348 17739 15351
rect 18230 15348 18236 15360
rect 17727 15320 18236 15348
rect 17727 15317 17739 15320
rect 17681 15311 17739 15317
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 1104 15258 18952 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 14246 15258
rect 14298 15206 14310 15258
rect 14362 15206 14374 15258
rect 14426 15206 14438 15258
rect 14490 15206 18952 15258
rect 1104 15184 18952 15206
rect 37628 15258 68816 15280
rect 37628 15206 44246 15258
rect 44298 15206 44310 15258
rect 44362 15206 44374 15258
rect 44426 15206 44438 15258
rect 44490 15206 54246 15258
rect 54298 15206 54310 15258
rect 54362 15206 54374 15258
rect 54426 15206 54438 15258
rect 54490 15206 64246 15258
rect 64298 15206 64310 15258
rect 64362 15206 64374 15258
rect 64426 15206 64438 15258
rect 64490 15206 68816 15258
rect 37628 15184 68816 15206
rect 9766 15144 9772 15156
rect 9727 15116 9772 15144
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 68094 15008 68100 15020
rect 68055 14980 68100 15008
rect 68094 14968 68100 14980
rect 68152 14968 68158 15020
rect 53742 14900 53748 14952
rect 53800 14940 53806 14952
rect 66349 14943 66407 14949
rect 66349 14940 66361 14943
rect 53800 14912 66361 14940
rect 53800 14900 53806 14912
rect 66349 14909 66361 14912
rect 66395 14909 66407 14943
rect 67174 14940 67180 14952
rect 67135 14912 67180 14940
rect 66349 14903 66407 14909
rect 67174 14900 67180 14912
rect 67232 14900 67238 14952
rect 67726 14900 67732 14952
rect 67784 14940 67790 14952
rect 67913 14943 67971 14949
rect 67913 14940 67925 14943
rect 67784 14912 67925 14940
rect 67784 14900 67790 14912
rect 67913 14909 67925 14912
rect 67959 14909 67971 14943
rect 67913 14903 67971 14909
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 4706 14872 4712 14884
rect 1995 14844 4712 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 2608 14816 2636 14844
rect 4706 14832 4712 14844
rect 4764 14832 4770 14884
rect 17313 14875 17371 14881
rect 17313 14841 17325 14875
rect 17359 14872 17371 14875
rect 18506 14872 18512 14884
rect 17359 14844 18512 14872
rect 17359 14841 17371 14844
rect 17313 14835 17371 14841
rect 18506 14832 18512 14844
rect 18564 14832 18570 14884
rect 1854 14804 1860 14816
rect 1815 14776 1860 14804
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 2590 14804 2596 14816
rect 2551 14776 2596 14804
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 18233 14807 18291 14813
rect 18233 14773 18245 14807
rect 18279 14804 18291 14807
rect 18782 14804 18788 14816
rect 18279 14776 18788 14804
rect 18279 14773 18291 14776
rect 18233 14767 18291 14773
rect 18782 14764 18788 14776
rect 18840 14764 18846 14816
rect 1104 14714 18952 14736
rect 1104 14662 9246 14714
rect 9298 14662 9310 14714
rect 9362 14662 9374 14714
rect 9426 14662 9438 14714
rect 9490 14662 18952 14714
rect 1104 14640 18952 14662
rect 37628 14714 68816 14736
rect 37628 14662 39246 14714
rect 39298 14662 39310 14714
rect 39362 14662 39374 14714
rect 39426 14662 39438 14714
rect 39490 14662 49246 14714
rect 49298 14662 49310 14714
rect 49362 14662 49374 14714
rect 49426 14662 49438 14714
rect 49490 14662 59246 14714
rect 59298 14662 59310 14714
rect 59362 14662 59374 14714
rect 59426 14662 59438 14714
rect 59490 14662 68816 14714
rect 37628 14640 68816 14662
rect 15197 14603 15255 14609
rect 15197 14569 15209 14603
rect 15243 14600 15255 14603
rect 16022 14600 16028 14612
rect 15243 14572 16028 14600
rect 15243 14569 15255 14572
rect 15197 14563 15255 14569
rect 16022 14560 16028 14572
rect 16080 14600 16086 14612
rect 17126 14600 17132 14612
rect 16080 14572 17132 14600
rect 16080 14560 16086 14572
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 17310 14600 17316 14612
rect 17271 14572 17316 14600
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 18046 14532 18052 14544
rect 5684 14504 18052 14532
rect 5684 14492 5690 14504
rect 18046 14492 18052 14504
rect 18104 14492 18110 14544
rect 38102 14492 38108 14544
rect 38160 14532 38166 14544
rect 48590 14532 48596 14544
rect 38160 14504 48596 14532
rect 38160 14492 38166 14504
rect 48590 14492 48596 14504
rect 48648 14492 48654 14544
rect 6730 14424 6736 14476
rect 6788 14464 6794 14476
rect 12066 14464 12072 14476
rect 6788 14436 12072 14464
rect 6788 14424 6794 14436
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 18690 14464 18696 14476
rect 17184 14436 18696 14464
rect 17184 14424 17190 14436
rect 18690 14424 18696 14436
rect 18748 14464 18754 14476
rect 48774 14464 48780 14476
rect 18748 14436 48780 14464
rect 18748 14424 18754 14436
rect 48774 14424 48780 14436
rect 48832 14424 48838 14476
rect 55950 14424 55956 14476
rect 56008 14464 56014 14476
rect 67266 14464 67272 14476
rect 56008 14436 67272 14464
rect 56008 14424 56014 14436
rect 67266 14424 67272 14436
rect 67324 14424 67330 14476
rect 48682 14396 48688 14408
rect 16546 14368 48688 14396
rect 16546 14272 16574 14368
rect 48682 14356 48688 14368
rect 48740 14356 48746 14408
rect 16761 14331 16819 14337
rect 16761 14297 16773 14331
rect 16807 14328 16819 14331
rect 17402 14328 17408 14340
rect 16807 14300 17408 14328
rect 16807 14297 16819 14300
rect 16761 14291 16819 14297
rect 17402 14288 17408 14300
rect 17460 14328 17466 14340
rect 35710 14328 35716 14340
rect 17460 14300 35716 14328
rect 17460 14288 17466 14300
rect 35710 14288 35716 14300
rect 35768 14288 35774 14340
rect 16209 14263 16267 14269
rect 16209 14229 16221 14263
rect 16255 14260 16267 14263
rect 16482 14260 16488 14272
rect 16255 14232 16488 14260
rect 16255 14229 16267 14232
rect 16209 14223 16267 14229
rect 16482 14220 16488 14232
rect 16540 14232 16574 14272
rect 16540 14220 16546 14232
rect 17678 14220 17684 14272
rect 17736 14260 17742 14272
rect 17865 14263 17923 14269
rect 17865 14260 17877 14263
rect 17736 14232 17877 14260
rect 17736 14220 17742 14232
rect 17865 14229 17877 14232
rect 17911 14260 17923 14263
rect 17954 14260 17960 14272
rect 17911 14232 17960 14260
rect 17911 14229 17923 14232
rect 17865 14223 17923 14229
rect 17954 14220 17960 14232
rect 18012 14220 18018 14272
rect 38194 14260 38200 14272
rect 38107 14232 38200 14260
rect 38194 14220 38200 14232
rect 38252 14260 38258 14272
rect 38378 14260 38384 14272
rect 38252 14232 38384 14260
rect 38252 14220 38258 14232
rect 38378 14220 38384 14232
rect 38436 14220 38442 14272
rect 51810 14220 51816 14272
rect 51868 14260 51874 14272
rect 55858 14260 55864 14272
rect 51868 14232 55864 14260
rect 51868 14220 51874 14232
rect 55858 14220 55864 14232
rect 55916 14220 55922 14272
rect 58434 14220 58440 14272
rect 58492 14260 58498 14272
rect 65334 14260 65340 14272
rect 58492 14232 65340 14260
rect 58492 14220 58498 14232
rect 65334 14220 65340 14232
rect 65392 14220 65398 14272
rect 67634 14220 67640 14272
rect 67692 14260 67698 14272
rect 67729 14263 67787 14269
rect 67729 14260 67741 14263
rect 67692 14232 67741 14260
rect 67692 14220 67698 14232
rect 67729 14229 67741 14232
rect 67775 14229 67787 14263
rect 67729 14223 67787 14229
rect 1104 14170 18952 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 14246 14170
rect 14298 14118 14310 14170
rect 14362 14118 14374 14170
rect 14426 14118 14438 14170
rect 14490 14118 18952 14170
rect 1104 14096 18952 14118
rect 37628 14170 68816 14192
rect 37628 14118 44246 14170
rect 44298 14118 44310 14170
rect 44362 14118 44374 14170
rect 44426 14118 44438 14170
rect 44490 14118 54246 14170
rect 54298 14118 54310 14170
rect 54362 14118 54374 14170
rect 54426 14118 54438 14170
rect 54490 14118 64246 14170
rect 64298 14118 64310 14170
rect 64362 14118 64374 14170
rect 64426 14118 64438 14170
rect 64490 14118 68816 14170
rect 37628 14096 68816 14118
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 17586 14056 17592 14068
rect 13136 14028 17592 14056
rect 13136 14016 13142 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 18046 14056 18052 14068
rect 18007 14028 18052 14056
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 55122 14056 55128 14068
rect 26206 14028 55128 14056
rect 14642 13988 14648 14000
rect 14603 13960 14648 13988
rect 14642 13948 14648 13960
rect 14700 13948 14706 14000
rect 26206 13988 26234 14028
rect 55122 14016 55128 14028
rect 55180 14016 55186 14068
rect 66438 14016 66444 14068
rect 66496 14056 66502 14068
rect 67269 14059 67327 14065
rect 67269 14056 67281 14059
rect 66496 14028 67281 14056
rect 66496 14016 66502 14028
rect 67269 14025 67281 14028
rect 67315 14025 67327 14059
rect 67269 14019 67327 14025
rect 38102 13988 38108 14000
rect 16316 13960 26234 13988
rect 38063 13960 38108 13988
rect 16316 13864 16344 13960
rect 38102 13948 38108 13960
rect 38160 13948 38166 14000
rect 38562 13948 38568 14000
rect 38620 13988 38626 14000
rect 39117 13991 39175 13997
rect 39117 13988 39129 13991
rect 38620 13960 39129 13988
rect 38620 13948 38626 13960
rect 39117 13957 39129 13960
rect 39163 13957 39175 13991
rect 39117 13951 39175 13957
rect 39758 13948 39764 14000
rect 39816 13988 39822 14000
rect 46198 13988 46204 14000
rect 39816 13960 46204 13988
rect 39816 13948 39822 13960
rect 46198 13948 46204 13960
rect 46256 13948 46262 14000
rect 47394 13920 47400 13932
rect 16408 13892 47400 13920
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14090 13852 14096 13864
rect 14047 13824 14096 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13852 15255 13855
rect 15654 13852 15660 13864
rect 15243 13824 15660 13852
rect 15243 13821 15255 13824
rect 15197 13815 15255 13821
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15838 13852 15844 13864
rect 15799 13824 15844 13852
rect 15838 13812 15844 13824
rect 15896 13852 15902 13864
rect 16298 13852 16304 13864
rect 15896 13824 16160 13852
rect 16259 13824 16304 13852
rect 15896 13812 15902 13824
rect 16132 13784 16160 13824
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 16408 13784 16436 13892
rect 47394 13880 47400 13892
rect 47452 13880 47458 13932
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13852 17095 13855
rect 17126 13852 17132 13864
rect 17083 13824 17132 13852
rect 17083 13821 17095 13824
rect 17037 13815 17095 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 17586 13852 17592 13864
rect 17499 13824 17592 13852
rect 17586 13812 17592 13824
rect 17644 13852 17650 13864
rect 18598 13852 18604 13864
rect 17644 13824 18604 13852
rect 17644 13812 17650 13824
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 37642 13812 37648 13864
rect 37700 13852 37706 13864
rect 37918 13852 37924 13864
rect 37700 13824 37924 13852
rect 37700 13812 37706 13824
rect 37918 13812 37924 13824
rect 37976 13852 37982 13864
rect 38657 13855 38715 13861
rect 38657 13852 38669 13855
rect 37976 13824 38669 13852
rect 37976 13812 37982 13824
rect 38657 13821 38669 13824
rect 38703 13821 38715 13855
rect 39758 13852 39764 13864
rect 39719 13824 39764 13852
rect 38657 13815 38715 13821
rect 39758 13812 39764 13824
rect 39816 13812 39822 13864
rect 67284 13852 67312 14019
rect 67913 13855 67971 13861
rect 67913 13852 67925 13855
rect 67284 13824 67925 13852
rect 67913 13821 67925 13824
rect 67959 13821 67971 13855
rect 68094 13852 68100 13864
rect 68055 13824 68100 13852
rect 67913 13815 67971 13821
rect 68094 13812 68100 13824
rect 68152 13812 68158 13864
rect 53834 13784 53840 13796
rect 16132 13756 16436 13784
rect 16546 13756 53840 13784
rect 14090 13676 14096 13728
rect 14148 13716 14154 13728
rect 16546 13716 16574 13756
rect 53834 13744 53840 13756
rect 53892 13744 53898 13796
rect 14148 13688 16574 13716
rect 14148 13676 14154 13688
rect 1104 13626 18952 13648
rect 1104 13574 9246 13626
rect 9298 13574 9310 13626
rect 9362 13574 9374 13626
rect 9426 13574 9438 13626
rect 9490 13574 18952 13626
rect 1104 13552 18952 13574
rect 37628 13626 68816 13648
rect 37628 13574 39246 13626
rect 39298 13574 39310 13626
rect 39362 13574 39374 13626
rect 39426 13574 39438 13626
rect 39490 13574 49246 13626
rect 49298 13574 49310 13626
rect 49362 13574 49374 13626
rect 49426 13574 49438 13626
rect 49490 13574 59246 13626
rect 59298 13574 59310 13626
rect 59362 13574 59374 13626
rect 59426 13574 59438 13626
rect 59490 13574 68816 13626
rect 37628 13552 68816 13574
rect 1854 13512 1860 13524
rect 1815 13484 1860 13512
rect 1854 13472 1860 13484
rect 1912 13472 1918 13524
rect 12250 13512 12256 13524
rect 12211 13484 12256 13512
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 21361 13515 21419 13521
rect 21361 13481 21373 13515
rect 21407 13512 21419 13515
rect 62942 13512 62948 13524
rect 21407 13484 62948 13512
rect 21407 13481 21419 13484
rect 21361 13475 21419 13481
rect 62942 13472 62948 13484
rect 63000 13472 63006 13524
rect 1949 13447 2007 13453
rect 1949 13413 1961 13447
rect 1995 13444 2007 13447
rect 2314 13444 2320 13456
rect 1995 13416 2320 13444
rect 1995 13413 2007 13416
rect 1949 13407 2007 13413
rect 2314 13404 2320 13416
rect 2372 13404 2378 13456
rect 2406 13404 2412 13456
rect 2464 13444 2470 13456
rect 2464 13416 26234 13444
rect 2464 13404 2470 13416
rect 13354 13336 13360 13388
rect 13412 13376 13418 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 13412 13348 21373 13376
rect 13412 13336 13418 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 26206 13376 26234 13416
rect 40034 13404 40040 13456
rect 40092 13444 40098 13456
rect 40678 13444 40684 13456
rect 40092 13416 40684 13444
rect 40092 13404 40098 13416
rect 40678 13404 40684 13416
rect 40736 13404 40742 13456
rect 41138 13404 41144 13456
rect 41196 13444 41202 13456
rect 41196 13416 45554 13444
rect 41196 13404 41202 13416
rect 45526 13376 45554 13416
rect 55306 13376 55312 13388
rect 26206 13348 41552 13376
rect 45526 13348 55312 13376
rect 21361 13339 21419 13345
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 37369 13311 37427 13317
rect 37369 13308 37381 13311
rect 14967 13280 37381 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 37369 13277 37381 13280
rect 37415 13277 37427 13311
rect 37369 13271 37427 13277
rect 37458 13268 37464 13320
rect 37516 13308 37522 13320
rect 38657 13311 38715 13317
rect 38657 13308 38669 13311
rect 37516 13280 38669 13308
rect 37516 13268 37522 13280
rect 38657 13277 38669 13280
rect 38703 13308 38715 13311
rect 40034 13308 40040 13320
rect 38703 13280 40040 13308
rect 38703 13277 38715 13280
rect 38657 13271 38715 13277
rect 40034 13268 40040 13280
rect 40092 13268 40098 13320
rect 40126 13268 40132 13320
rect 40184 13308 40190 13320
rect 40957 13311 41015 13317
rect 40957 13308 40969 13311
rect 40184 13280 40969 13308
rect 40184 13268 40190 13280
rect 40957 13277 40969 13280
rect 41003 13277 41015 13311
rect 41524 13308 41552 13348
rect 55306 13336 55312 13348
rect 55364 13336 55370 13388
rect 43162 13308 43168 13320
rect 41524 13280 43168 13308
rect 40957 13271 41015 13277
rect 43162 13268 43168 13280
rect 43220 13308 43226 13320
rect 51902 13308 51908 13320
rect 43220 13280 51908 13308
rect 43220 13268 43226 13280
rect 51902 13268 51908 13280
rect 51960 13268 51966 13320
rect 2685 13243 2743 13249
rect 2685 13209 2697 13243
rect 2731 13240 2743 13243
rect 15562 13240 15568 13252
rect 2731 13212 15568 13240
rect 2731 13209 2743 13212
rect 2685 13203 2743 13209
rect 15562 13200 15568 13212
rect 15620 13200 15626 13252
rect 15657 13243 15715 13249
rect 15657 13209 15669 13243
rect 15703 13240 15715 13243
rect 16298 13240 16304 13252
rect 15703 13212 16304 13240
rect 15703 13209 15715 13212
rect 15657 13203 15715 13209
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 18233 13243 18291 13249
rect 18233 13209 18245 13243
rect 18279 13240 18291 13243
rect 55674 13240 55680 13252
rect 18279 13212 55680 13240
rect 18279 13209 18291 13212
rect 18233 13203 18291 13209
rect 55674 13200 55680 13212
rect 55732 13200 55738 13252
rect 13538 13172 13544 13184
rect 13499 13144 13544 13172
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 16117 13175 16175 13181
rect 16117 13172 16129 13175
rect 15988 13144 16129 13172
rect 15988 13132 15994 13144
rect 16117 13141 16129 13144
rect 16163 13172 16175 13175
rect 16390 13172 16396 13184
rect 16163 13144 16396 13172
rect 16163 13141 16175 13144
rect 16117 13135 16175 13141
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 16758 13172 16764 13184
rect 16719 13144 16764 13172
rect 16758 13132 16764 13144
rect 16816 13132 16822 13184
rect 17589 13175 17647 13181
rect 17589 13141 17601 13175
rect 17635 13172 17647 13175
rect 18414 13172 18420 13184
rect 17635 13144 18420 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 37734 13132 37740 13184
rect 37792 13172 37798 13184
rect 37921 13175 37979 13181
rect 37921 13172 37933 13175
rect 37792 13144 37933 13172
rect 37792 13132 37798 13144
rect 37921 13141 37933 13144
rect 37967 13141 37979 13175
rect 39206 13172 39212 13184
rect 39167 13144 39212 13172
rect 37921 13135 37979 13141
rect 39206 13132 39212 13144
rect 39264 13132 39270 13184
rect 39666 13132 39672 13184
rect 39724 13172 39730 13184
rect 39761 13175 39819 13181
rect 39761 13172 39773 13175
rect 39724 13144 39773 13172
rect 39724 13132 39730 13144
rect 39761 13141 39773 13144
rect 39807 13141 39819 13175
rect 39761 13135 39819 13141
rect 40310 13132 40316 13184
rect 40368 13172 40374 13184
rect 40405 13175 40463 13181
rect 40405 13172 40417 13175
rect 40368 13144 40417 13172
rect 40368 13132 40374 13144
rect 40405 13141 40417 13144
rect 40451 13172 40463 13175
rect 41138 13172 41144 13184
rect 40451 13144 41144 13172
rect 40451 13141 40463 13144
rect 40405 13135 40463 13141
rect 41138 13132 41144 13144
rect 41196 13132 41202 13184
rect 41601 13175 41659 13181
rect 41601 13141 41613 13175
rect 41647 13172 41659 13175
rect 41966 13172 41972 13184
rect 41647 13144 41972 13172
rect 41647 13141 41659 13144
rect 41601 13135 41659 13141
rect 41966 13132 41972 13144
rect 42024 13132 42030 13184
rect 1104 13082 18952 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 14246 13082
rect 14298 13030 14310 13082
rect 14362 13030 14374 13082
rect 14426 13030 14438 13082
rect 14490 13030 18952 13082
rect 1104 13008 18952 13030
rect 37628 13082 68816 13104
rect 37628 13030 44246 13082
rect 44298 13030 44310 13082
rect 44362 13030 44374 13082
rect 44426 13030 44438 13082
rect 44490 13030 54246 13082
rect 54298 13030 54310 13082
rect 54362 13030 54374 13082
rect 54426 13030 54438 13082
rect 54490 13030 64246 13082
rect 64298 13030 64310 13082
rect 64362 13030 64374 13082
rect 64426 13030 64438 13082
rect 64490 13030 68816 13082
rect 37628 13008 68816 13030
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2314 12968 2320 12980
rect 2271 12940 2320 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 15470 12968 15476 12980
rect 14783 12940 15476 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 17221 12971 17279 12977
rect 17221 12937 17233 12971
rect 17267 12968 17279 12971
rect 18138 12968 18144 12980
rect 17267 12940 18144 12968
rect 17267 12937 17279 12940
rect 17221 12931 17279 12937
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 38286 12928 38292 12980
rect 38344 12968 38350 12980
rect 38746 12968 38752 12980
rect 38344 12940 38752 12968
rect 38344 12928 38350 12940
rect 38746 12928 38752 12940
rect 38804 12968 38810 12980
rect 39025 12971 39083 12977
rect 39025 12968 39037 12971
rect 38804 12940 39037 12968
rect 38804 12928 38810 12940
rect 39025 12937 39037 12940
rect 39071 12937 39083 12971
rect 39025 12931 39083 12937
rect 39942 12928 39948 12980
rect 40000 12968 40006 12980
rect 40129 12971 40187 12977
rect 40129 12968 40141 12971
rect 40000 12940 40141 12968
rect 40000 12928 40006 12940
rect 40129 12937 40141 12940
rect 40175 12937 40187 12971
rect 53834 12968 53840 12980
rect 53795 12940 53840 12968
rect 40129 12931 40187 12937
rect 53834 12928 53840 12940
rect 53892 12928 53898 12980
rect 15746 12900 15752 12912
rect 15707 12872 15752 12900
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 37369 12903 37427 12909
rect 37369 12869 37381 12903
rect 37415 12900 37427 12903
rect 40954 12900 40960 12912
rect 37415 12872 40960 12900
rect 37415 12869 37427 12872
rect 37369 12863 37427 12869
rect 40954 12860 40960 12872
rect 41012 12860 41018 12912
rect 42610 12900 42616 12912
rect 41432 12872 42616 12900
rect 16298 12792 16304 12844
rect 16356 12832 16362 12844
rect 23290 12832 23296 12844
rect 16356 12804 23296 12832
rect 16356 12792 16362 12804
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 37550 12792 37556 12844
rect 37608 12832 37614 12844
rect 40310 12832 40316 12844
rect 37608 12804 40316 12832
rect 37608 12792 37614 12804
rect 40310 12792 40316 12804
rect 40368 12792 40374 12844
rect 16209 12767 16267 12773
rect 16209 12764 16221 12767
rect 15396 12736 16221 12764
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 14093 12699 14151 12705
rect 14093 12696 14105 12699
rect 10560 12668 14105 12696
rect 10560 12656 10566 12668
rect 14093 12665 14105 12668
rect 14139 12696 14151 12699
rect 15197 12699 15255 12705
rect 15197 12696 15209 12699
rect 14139 12668 15209 12696
rect 14139 12665 14151 12668
rect 14093 12659 14151 12665
rect 15197 12665 15209 12668
rect 15243 12665 15255 12699
rect 15197 12659 15255 12665
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 12216 12600 12265 12628
rect 12216 12588 12222 12600
rect 12253 12597 12265 12600
rect 12299 12597 12311 12631
rect 12253 12591 12311 12597
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12768 12600 12817 12628
rect 12768 12588 12774 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 13354 12628 13360 12640
rect 13315 12600 13360 12628
rect 12805 12591 12863 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 15396 12637 15424 12736
rect 16209 12733 16221 12736
rect 16255 12764 16267 12767
rect 19978 12764 19984 12776
rect 16255 12736 19984 12764
rect 16255 12733 16267 12736
rect 16209 12727 16267 12733
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 40586 12724 40592 12776
rect 40644 12764 40650 12776
rect 41432 12773 41460 12872
rect 42610 12860 42616 12872
rect 42668 12860 42674 12912
rect 53282 12832 53288 12844
rect 41984 12804 53288 12832
rect 41417 12767 41475 12773
rect 41417 12764 41429 12767
rect 40644 12736 41429 12764
rect 40644 12724 40650 12736
rect 41417 12733 41429 12736
rect 41463 12733 41475 12767
rect 41417 12727 41475 12733
rect 15565 12699 15623 12705
rect 15565 12665 15577 12699
rect 15611 12696 15623 12699
rect 16114 12696 16120 12708
rect 15611 12668 16120 12696
rect 15611 12665 15623 12668
rect 15565 12659 15623 12665
rect 16114 12656 16120 12668
rect 16172 12656 16178 12708
rect 37182 12656 37188 12708
rect 37240 12696 37246 12708
rect 38473 12699 38531 12705
rect 38473 12696 38485 12699
rect 37240 12668 38485 12696
rect 37240 12656 37246 12668
rect 38473 12665 38485 12668
rect 38519 12665 38531 12699
rect 38473 12659 38531 12665
rect 40678 12656 40684 12708
rect 40736 12696 40742 12708
rect 41984 12705 42012 12804
rect 53282 12792 53288 12804
rect 53340 12792 53346 12844
rect 65242 12764 65248 12776
rect 42352 12736 47992 12764
rect 41969 12699 42027 12705
rect 41969 12696 41981 12699
rect 40736 12668 41981 12696
rect 40736 12656 40742 12668
rect 41969 12665 41981 12668
rect 42015 12665 42027 12699
rect 41969 12659 42027 12665
rect 15381 12631 15439 12637
rect 15381 12597 15393 12631
rect 15427 12597 15439 12631
rect 15381 12591 15439 12597
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 15528 12600 15573 12628
rect 15528 12588 15534 12600
rect 17586 12588 17592 12640
rect 17644 12628 17650 12640
rect 17681 12631 17739 12637
rect 17681 12628 17693 12631
rect 17644 12600 17693 12628
rect 17644 12588 17650 12600
rect 17681 12597 17693 12600
rect 17727 12597 17739 12631
rect 17681 12591 17739 12597
rect 37826 12588 37832 12640
rect 37884 12628 37890 12640
rect 37921 12631 37979 12637
rect 37921 12628 37933 12631
rect 37884 12600 37933 12628
rect 37884 12588 37890 12600
rect 37921 12597 37933 12600
rect 37967 12597 37979 12631
rect 37921 12591 37979 12597
rect 39114 12588 39120 12640
rect 39172 12628 39178 12640
rect 39574 12628 39580 12640
rect 39172 12600 39580 12628
rect 39172 12588 39178 12600
rect 39574 12588 39580 12600
rect 39632 12588 39638 12640
rect 40862 12628 40868 12640
rect 40823 12600 40868 12628
rect 40862 12588 40868 12600
rect 40920 12628 40926 12640
rect 42352 12628 42380 12736
rect 42610 12656 42616 12708
rect 42668 12696 42674 12708
rect 47964 12696 47992 12736
rect 55186 12736 65248 12764
rect 55186 12696 55214 12736
rect 65242 12724 65248 12736
rect 65300 12724 65306 12776
rect 42668 12668 45554 12696
rect 47964 12668 55214 12696
rect 42668 12656 42674 12668
rect 40920 12600 42380 12628
rect 45526 12628 45554 12668
rect 53926 12628 53932 12640
rect 45526 12600 53932 12628
rect 40920 12588 40926 12600
rect 53926 12588 53932 12600
rect 53984 12588 53990 12640
rect 1104 12538 18952 12560
rect 1104 12486 9246 12538
rect 9298 12486 9310 12538
rect 9362 12486 9374 12538
rect 9426 12486 9438 12538
rect 9490 12486 18952 12538
rect 1104 12464 18952 12486
rect 37628 12538 68816 12560
rect 37628 12486 39246 12538
rect 39298 12486 39310 12538
rect 39362 12486 39374 12538
rect 39426 12486 39438 12538
rect 39490 12486 49246 12538
rect 49298 12486 49310 12538
rect 49362 12486 49374 12538
rect 49426 12486 49438 12538
rect 49490 12486 59246 12538
rect 59298 12486 59310 12538
rect 59362 12486 59374 12538
rect 59426 12486 59438 12538
rect 59490 12486 68816 12538
rect 37628 12464 68816 12486
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 23934 12424 23940 12436
rect 9732 12396 23940 12424
rect 9732 12384 9738 12396
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 12618 12356 12624 12368
rect 12579 12328 12624 12356
rect 12618 12316 12624 12328
rect 12676 12316 12682 12368
rect 16574 12356 16580 12368
rect 16535 12328 16580 12356
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 16942 12288 16948 12300
rect 12406 12260 16948 12288
rect 11149 12087 11207 12093
rect 11149 12053 11161 12087
rect 11195 12084 11207 12087
rect 11422 12084 11428 12096
rect 11195 12056 11428 12084
rect 11195 12053 11207 12056
rect 11149 12047 11207 12053
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11848 12056 12081 12084
rect 11848 12044 11854 12056
rect 12069 12053 12081 12056
rect 12115 12084 12127 12087
rect 12406 12084 12434 12260
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 18230 12288 18236 12300
rect 18191 12260 18236 12288
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 67453 12291 67511 12297
rect 67453 12257 67465 12291
rect 67499 12288 67511 12291
rect 68094 12288 68100 12300
rect 67499 12260 68100 12288
rect 67499 12257 67511 12260
rect 67453 12251 67511 12257
rect 68094 12248 68100 12260
rect 68152 12248 68158 12300
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 13814 12220 13820 12232
rect 13311 12192 13820 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18046 12220 18052 12232
rect 18003 12192 18052 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 39758 12180 39764 12232
rect 39816 12220 39822 12232
rect 41509 12223 41567 12229
rect 41509 12220 41521 12223
rect 39816 12192 41521 12220
rect 39816 12180 39822 12192
rect 41509 12189 41521 12192
rect 41555 12189 41567 12223
rect 41509 12183 41567 12189
rect 39850 12112 39856 12164
rect 39908 12152 39914 12164
rect 42061 12155 42119 12161
rect 42061 12152 42073 12155
rect 39908 12124 42073 12152
rect 39908 12112 39914 12124
rect 42061 12121 42073 12124
rect 42107 12121 42119 12155
rect 42061 12115 42119 12121
rect 12115 12056 12434 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13504 12056 13829 12084
rect 13504 12044 13510 12056
rect 13817 12053 13829 12056
rect 13863 12053 13875 12087
rect 13817 12047 13875 12053
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 14734 12084 14740 12096
rect 14691 12056 14740 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15194 12084 15200 12096
rect 15068 12056 15200 12084
rect 15068 12044 15074 12056
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 38102 12084 38108 12096
rect 38063 12056 38108 12084
rect 38102 12044 38108 12056
rect 38160 12044 38166 12096
rect 38194 12044 38200 12096
rect 38252 12084 38258 12096
rect 38657 12087 38715 12093
rect 38657 12084 38669 12087
rect 38252 12056 38669 12084
rect 38252 12044 38258 12056
rect 38657 12053 38669 12056
rect 38703 12053 38715 12087
rect 39114 12084 39120 12096
rect 39075 12056 39120 12084
rect 38657 12047 38715 12053
rect 39114 12044 39120 12056
rect 39172 12044 39178 12096
rect 39758 12084 39764 12096
rect 39719 12056 39764 12084
rect 39758 12044 39764 12056
rect 39816 12044 39822 12096
rect 40310 12044 40316 12096
rect 40368 12084 40374 12096
rect 40405 12087 40463 12093
rect 40405 12084 40417 12087
rect 40368 12056 40417 12084
rect 40368 12044 40374 12056
rect 40405 12053 40417 12056
rect 40451 12053 40463 12087
rect 40954 12084 40960 12096
rect 40915 12056 40960 12084
rect 40405 12047 40463 12053
rect 40954 12044 40960 12056
rect 41012 12044 41018 12096
rect 42702 12084 42708 12096
rect 42663 12056 42708 12084
rect 42702 12044 42708 12056
rect 42760 12044 42766 12096
rect 43254 12084 43260 12096
rect 43215 12056 43260 12084
rect 43254 12044 43260 12056
rect 43312 12044 43318 12096
rect 48041 12087 48099 12093
rect 48041 12053 48053 12087
rect 48087 12084 48099 12087
rect 48682 12084 48688 12096
rect 48087 12056 48688 12084
rect 48087 12053 48099 12056
rect 48041 12047 48099 12053
rect 48682 12044 48688 12056
rect 48740 12044 48746 12096
rect 1104 11994 18952 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 14246 11994
rect 14298 11942 14310 11994
rect 14362 11942 14374 11994
rect 14426 11942 14438 11994
rect 14490 11942 18952 11994
rect 1104 11920 18952 11942
rect 37628 11994 68816 12016
rect 37628 11942 44246 11994
rect 44298 11942 44310 11994
rect 44362 11942 44374 11994
rect 44426 11942 44438 11994
rect 44490 11942 54246 11994
rect 54298 11942 54310 11994
rect 54362 11942 54374 11994
rect 54426 11942 54438 11994
rect 54490 11942 64246 11994
rect 64298 11942 64310 11994
rect 64362 11942 64374 11994
rect 64426 11942 64438 11994
rect 64490 11942 68816 11994
rect 37628 11920 68816 11942
rect 38010 11880 38016 11892
rect 37971 11852 38016 11880
rect 38010 11840 38016 11852
rect 38068 11840 38074 11892
rect 41969 11883 42027 11889
rect 41969 11849 41981 11883
rect 42015 11880 42027 11883
rect 42150 11880 42156 11892
rect 42015 11852 42156 11880
rect 42015 11849 42027 11852
rect 41969 11843 42027 11849
rect 42150 11840 42156 11852
rect 42208 11880 42214 11892
rect 45646 11880 45652 11892
rect 42208 11852 45652 11880
rect 42208 11840 42214 11852
rect 45646 11840 45652 11852
rect 45704 11840 45710 11892
rect 38102 11772 38108 11824
rect 38160 11812 38166 11824
rect 53006 11812 53012 11824
rect 38160 11784 53012 11812
rect 38160 11772 38166 11784
rect 53006 11772 53012 11784
rect 53064 11772 53070 11824
rect 62114 11772 62120 11824
rect 62172 11812 62178 11824
rect 65058 11812 65064 11824
rect 62172 11784 65064 11812
rect 62172 11772 62178 11784
rect 65058 11772 65064 11784
rect 65116 11772 65122 11824
rect 45554 11704 45560 11756
rect 45612 11744 45618 11756
rect 53190 11744 53196 11756
rect 45612 11716 53196 11744
rect 45612 11704 45618 11716
rect 53190 11704 53196 11716
rect 53248 11704 53254 11756
rect 38105 11679 38163 11685
rect 38105 11645 38117 11679
rect 38151 11676 38163 11679
rect 38286 11676 38292 11688
rect 38151 11648 38292 11676
rect 38151 11645 38163 11648
rect 38105 11639 38163 11645
rect 38286 11636 38292 11648
rect 38344 11636 38350 11688
rect 38654 11636 38660 11688
rect 38712 11676 38718 11688
rect 39117 11679 39175 11685
rect 39117 11676 39129 11679
rect 38712 11648 39129 11676
rect 38712 11636 38718 11648
rect 39117 11645 39129 11648
rect 39163 11645 39175 11679
rect 67174 11676 67180 11688
rect 39117 11639 39175 11645
rect 44100 11648 67180 11676
rect 9950 11568 9956 11620
rect 10008 11608 10014 11620
rect 10689 11611 10747 11617
rect 10689 11608 10701 11611
rect 10008 11580 10701 11608
rect 10008 11568 10014 11580
rect 10689 11577 10701 11580
rect 10735 11577 10747 11611
rect 10689 11571 10747 11577
rect 42242 11568 42248 11620
rect 42300 11608 42306 11620
rect 42426 11608 42432 11620
rect 42300 11580 42432 11608
rect 42300 11568 42306 11580
rect 42426 11568 42432 11580
rect 42484 11608 42490 11620
rect 43533 11611 43591 11617
rect 43533 11608 43545 11611
rect 42484 11580 43545 11608
rect 42484 11568 42490 11580
rect 43533 11577 43545 11580
rect 43579 11577 43591 11611
rect 43533 11571 43591 11577
rect 10134 11540 10140 11552
rect 10095 11512 10140 11540
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 12032 11512 12173 11540
rect 12032 11500 12038 11512
rect 12161 11509 12173 11512
rect 12207 11540 12219 11543
rect 12342 11540 12348 11552
rect 12207 11512 12348 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12676 11512 12817 11540
rect 12676 11500 12682 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 13044 11512 13369 11540
rect 13044 11500 13050 11512
rect 13357 11509 13369 11512
rect 13403 11509 13415 11543
rect 13357 11503 13415 11509
rect 14461 11543 14519 11549
rect 14461 11509 14473 11543
rect 14507 11540 14519 11543
rect 14826 11540 14832 11552
rect 14507 11512 14832 11540
rect 14507 11509 14519 11512
rect 14461 11503 14519 11509
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 15565 11543 15623 11549
rect 14976 11512 15021 11540
rect 14976 11500 14982 11512
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 15654 11540 15660 11552
rect 15611 11512 15660 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 16482 11540 16488 11552
rect 16255 11512 16488 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 16942 11540 16948 11552
rect 16903 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17678 11540 17684 11552
rect 17639 11512 17684 11540
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18141 11543 18199 11549
rect 18141 11540 18153 11543
rect 18104 11512 18153 11540
rect 18104 11500 18110 11512
rect 18141 11509 18153 11512
rect 18187 11509 18199 11543
rect 18141 11503 18199 11509
rect 38470 11500 38476 11552
rect 38528 11540 38534 11552
rect 38657 11543 38715 11549
rect 38657 11540 38669 11543
rect 38528 11512 38669 11540
rect 38528 11500 38534 11512
rect 38657 11509 38669 11512
rect 38703 11509 38715 11543
rect 38657 11503 38715 11509
rect 39761 11543 39819 11549
rect 39761 11509 39773 11543
rect 39807 11540 39819 11543
rect 40126 11540 40132 11552
rect 39807 11512 40132 11540
rect 39807 11509 39819 11512
rect 39761 11503 39819 11509
rect 40126 11500 40132 11512
rect 40184 11500 40190 11552
rect 40405 11543 40463 11549
rect 40405 11509 40417 11543
rect 40451 11540 40463 11543
rect 40494 11540 40500 11552
rect 40451 11512 40500 11540
rect 40451 11509 40463 11512
rect 40405 11503 40463 11509
rect 40494 11500 40500 11512
rect 40552 11500 40558 11552
rect 41046 11540 41052 11552
rect 41007 11512 41052 11540
rect 41046 11500 41052 11512
rect 41104 11500 41110 11552
rect 42886 11500 42892 11552
rect 42944 11540 42950 11552
rect 42981 11543 43039 11549
rect 42981 11540 42993 11543
rect 42944 11512 42993 11540
rect 42944 11500 42950 11512
rect 42981 11509 42993 11512
rect 43027 11540 43039 11543
rect 44100 11540 44128 11648
rect 67174 11636 67180 11648
rect 67232 11636 67238 11688
rect 44177 11611 44235 11617
rect 44177 11577 44189 11611
rect 44223 11608 44235 11611
rect 45554 11608 45560 11620
rect 44223 11580 45560 11608
rect 44223 11577 44235 11580
rect 44177 11571 44235 11577
rect 45554 11568 45560 11580
rect 45612 11568 45618 11620
rect 45646 11568 45652 11620
rect 45704 11608 45710 11620
rect 57698 11608 57704 11620
rect 45704 11580 57704 11608
rect 45704 11568 45710 11580
rect 57698 11568 57704 11580
rect 57756 11568 57762 11620
rect 44634 11540 44640 11552
rect 43027 11512 44128 11540
rect 44595 11512 44640 11540
rect 43027 11509 43039 11512
rect 42981 11503 43039 11509
rect 44634 11500 44640 11512
rect 44692 11500 44698 11552
rect 65978 11500 65984 11552
rect 66036 11540 66042 11552
rect 66073 11543 66131 11549
rect 66073 11540 66085 11543
rect 66036 11512 66085 11540
rect 66036 11500 66042 11512
rect 66073 11509 66085 11512
rect 66119 11540 66131 11543
rect 66346 11540 66352 11552
rect 66119 11512 66352 11540
rect 66119 11509 66131 11512
rect 66073 11503 66131 11509
rect 66346 11500 66352 11512
rect 66404 11500 66410 11552
rect 66622 11540 66628 11552
rect 66583 11512 66628 11540
rect 66622 11500 66628 11512
rect 66680 11500 66686 11552
rect 67082 11500 67088 11552
rect 67140 11540 67146 11552
rect 67177 11543 67235 11549
rect 67177 11540 67189 11543
rect 67140 11512 67189 11540
rect 67140 11500 67146 11512
rect 67177 11509 67189 11512
rect 67223 11540 67235 11543
rect 67358 11540 67364 11552
rect 67223 11512 67364 11540
rect 67223 11509 67235 11512
rect 67177 11503 67235 11509
rect 67358 11500 67364 11512
rect 67416 11500 67422 11552
rect 67634 11540 67640 11552
rect 67595 11512 67640 11540
rect 67634 11500 67640 11512
rect 67692 11500 67698 11552
rect 1104 11450 18952 11472
rect 1104 11398 9246 11450
rect 9298 11398 9310 11450
rect 9362 11398 9374 11450
rect 9426 11398 9438 11450
rect 9490 11398 18952 11450
rect 1104 11376 18952 11398
rect 37628 11450 68816 11472
rect 37628 11398 39246 11450
rect 39298 11398 39310 11450
rect 39362 11398 39374 11450
rect 39426 11398 39438 11450
rect 39490 11398 49246 11450
rect 49298 11398 49310 11450
rect 49362 11398 49374 11450
rect 49426 11398 49438 11450
rect 49490 11398 59246 11450
rect 59298 11398 59310 11450
rect 59362 11398 59374 11450
rect 59426 11398 59438 11450
rect 59490 11398 68816 11450
rect 37628 11376 68816 11398
rect 67266 11336 67272 11348
rect 48332 11308 60734 11336
rect 67227 11308 67272 11336
rect 13354 11268 13360 11280
rect 10980 11240 13360 11268
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1578 11160 1584 11172
rect 1636 11200 1642 11212
rect 2041 11203 2099 11209
rect 2041 11200 2053 11203
rect 1636 11172 2053 11200
rect 1636 11160 1642 11172
rect 2041 11169 2053 11172
rect 2087 11169 2099 11203
rect 2041 11163 2099 11169
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11200 9551 11203
rect 9674 11200 9680 11212
rect 9539 11172 9680 11200
rect 9539 11169 9551 11172
rect 9493 11163 9551 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10980 11144 11008 11240
rect 13354 11228 13360 11240
rect 13412 11228 13418 11280
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11200 11575 11203
rect 15102 11200 15108 11212
rect 11563 11172 15108 11200
rect 11563 11169 11575 11172
rect 11517 11163 11575 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 37918 11200 37924 11212
rect 37879 11172 37924 11200
rect 37918 11160 37924 11172
rect 37976 11160 37982 11212
rect 39758 11160 39764 11212
rect 39816 11200 39822 11212
rect 48332 11209 48360 11308
rect 48317 11203 48375 11209
rect 39816 11172 39896 11200
rect 39816 11160 39822 11172
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 10962 11132 10968 11144
rect 10091 11104 10968 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 10870 11064 10876 11076
rect 10652 11036 10876 11064
rect 10652 11024 10658 11036
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 11698 11024 11704 11076
rect 11756 11064 11762 11076
rect 11977 11067 12035 11073
rect 11977 11064 11989 11067
rect 11756 11036 11989 11064
rect 11756 11024 11762 11036
rect 11977 11033 11989 11036
rect 12023 11033 12035 11067
rect 11977 11027 12035 11033
rect 12621 11067 12679 11073
rect 12621 11033 12633 11067
rect 12667 11064 12679 11067
rect 12710 11064 12716 11076
rect 12667 11036 12716 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 13262 11024 13268 11076
rect 13320 11064 13326 11076
rect 13357 11067 13415 11073
rect 13357 11064 13369 11067
rect 13320 11036 13369 11064
rect 13320 11024 13326 11036
rect 13357 11033 13369 11036
rect 13403 11033 13415 11067
rect 13357 11027 13415 11033
rect 13906 11024 13912 11076
rect 13964 11064 13970 11076
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 13964 11036 14381 11064
rect 13964 11024 13970 11036
rect 14369 11033 14381 11036
rect 14415 11033 14427 11067
rect 14369 11027 14427 11033
rect 15289 11067 15347 11073
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 15378 11064 15384 11076
rect 15335 11036 15384 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 15470 11024 15476 11076
rect 15528 11064 15534 11076
rect 15841 11067 15899 11073
rect 15841 11064 15853 11067
rect 15528 11036 15853 11064
rect 15528 11024 15534 11036
rect 15841 11033 15853 11036
rect 15887 11033 15899 11067
rect 15841 11027 15899 11033
rect 16577 11067 16635 11073
rect 16577 11033 16589 11067
rect 16623 11064 16635 11067
rect 16666 11064 16672 11076
rect 16623 11036 16672 11064
rect 16623 11033 16635 11036
rect 16577 11027 16635 11033
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 17126 11064 17132 11076
rect 17087 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 17770 11064 17776 11076
rect 17731 11036 17776 11064
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 38102 11024 38108 11076
rect 38160 11064 38166 11076
rect 38657 11067 38715 11073
rect 38657 11064 38669 11067
rect 38160 11036 38669 11064
rect 38160 11024 38166 11036
rect 38657 11033 38669 11036
rect 38703 11033 38715 11067
rect 38657 11027 38715 11033
rect 38746 11024 38752 11076
rect 38804 11064 38810 11076
rect 39117 11067 39175 11073
rect 39117 11064 39129 11067
rect 38804 11036 39129 11064
rect 38804 11024 38810 11036
rect 39117 11033 39129 11036
rect 39163 11033 39175 11067
rect 39758 11064 39764 11076
rect 39719 11036 39764 11064
rect 39117 11027 39175 11033
rect 39758 11024 39764 11036
rect 39816 11024 39822 11076
rect 39666 10956 39672 11008
rect 39724 10996 39730 11008
rect 39868 10996 39896 11172
rect 48317 11169 48329 11203
rect 48363 11169 48375 11203
rect 60706 11200 60734 11308
rect 67266 11296 67272 11308
rect 67324 11296 67330 11348
rect 67284 11268 67312 11296
rect 67913 11271 67971 11277
rect 67913 11268 67925 11271
rect 67284 11240 67925 11268
rect 67913 11237 67925 11240
rect 67959 11237 67971 11271
rect 67913 11231 67971 11237
rect 67634 11200 67640 11212
rect 60706 11172 67640 11200
rect 48317 11163 48375 11169
rect 67634 11160 67640 11172
rect 67692 11160 67698 11212
rect 42426 11092 42432 11144
rect 42484 11132 42490 11144
rect 44269 11135 44327 11141
rect 44269 11132 44281 11135
rect 42484 11104 44281 11132
rect 42484 11092 42490 11104
rect 44269 11101 44281 11104
rect 44315 11101 44327 11135
rect 51258 11132 51264 11144
rect 44269 11095 44327 11101
rect 44836 11104 51264 11132
rect 40034 11024 40040 11076
rect 40092 11064 40098 11076
rect 40405 11067 40463 11073
rect 40405 11064 40417 11067
rect 40092 11036 40417 11064
rect 40092 11024 40098 11036
rect 40405 11033 40417 11036
rect 40451 11033 40463 11067
rect 40405 11027 40463 11033
rect 40862 11024 40868 11076
rect 40920 11064 40926 11076
rect 40957 11067 41015 11073
rect 40957 11064 40969 11067
rect 40920 11036 40969 11064
rect 40920 11024 40926 11036
rect 40957 11033 40969 11036
rect 41003 11033 41015 11067
rect 40957 11027 41015 11033
rect 41414 11024 41420 11076
rect 41472 11064 41478 11076
rect 41509 11067 41567 11073
rect 41509 11064 41521 11067
rect 41472 11036 41521 11064
rect 41472 11024 41478 11036
rect 41509 11033 41521 11036
rect 41555 11033 41567 11067
rect 42058 11064 42064 11076
rect 42019 11036 42064 11064
rect 41509 11027 41567 11033
rect 42058 11024 42064 11036
rect 42116 11024 42122 11076
rect 42150 11024 42156 11076
rect 42208 11064 42214 11076
rect 42610 11064 42616 11076
rect 42208 11036 42380 11064
rect 42571 11036 42616 11064
rect 42208 11024 42214 11036
rect 42352 11008 42380 11036
rect 42610 11024 42616 11036
rect 42668 11024 42674 11076
rect 42702 11024 42708 11076
rect 42760 11064 42766 11076
rect 43165 11067 43223 11073
rect 43165 11064 43177 11067
rect 42760 11036 43177 11064
rect 42760 11024 42766 11036
rect 43165 11033 43177 11036
rect 43211 11033 43223 11067
rect 43806 11064 43812 11076
rect 43767 11036 43812 11064
rect 43165 11027 43223 11033
rect 43806 11024 43812 11036
rect 43864 11024 43870 11076
rect 44542 11024 44548 11076
rect 44600 11064 44606 11076
rect 44836 11073 44864 11104
rect 51258 11092 51264 11104
rect 51316 11092 51322 11144
rect 65426 11092 65432 11144
rect 65484 11132 65490 11144
rect 65521 11135 65579 11141
rect 65521 11132 65533 11135
rect 65484 11104 65533 11132
rect 65484 11092 65490 11104
rect 65521 11101 65533 11104
rect 65567 11132 65579 11135
rect 66530 11132 66536 11144
rect 65567 11104 66536 11132
rect 65567 11101 65579 11104
rect 65521 11095 65579 11101
rect 66530 11092 66536 11104
rect 66588 11092 66594 11144
rect 44821 11067 44879 11073
rect 44821 11064 44833 11067
rect 44600 11036 44833 11064
rect 44600 11024 44606 11036
rect 44821 11033 44833 11036
rect 44867 11033 44879 11067
rect 44821 11027 44879 11033
rect 45094 11024 45100 11076
rect 45152 11064 45158 11076
rect 45462 11064 45468 11076
rect 45152 11036 45468 11064
rect 45152 11024 45158 11036
rect 45462 11024 45468 11036
rect 45520 11064 45526 11076
rect 45649 11067 45707 11073
rect 45649 11064 45661 11067
rect 45520 11036 45661 11064
rect 45520 11024 45526 11036
rect 45649 11033 45661 11036
rect 45695 11033 45707 11067
rect 45649 11027 45707 11033
rect 65886 11024 65892 11076
rect 65944 11064 65950 11076
rect 66070 11064 66076 11076
rect 65944 11036 66076 11064
rect 65944 11024 65950 11036
rect 66070 11024 66076 11036
rect 66128 11024 66134 11076
rect 66806 11064 66812 11076
rect 66767 11036 66812 11064
rect 66806 11024 66812 11036
rect 66864 11024 66870 11076
rect 68094 11064 68100 11076
rect 68055 11036 68100 11064
rect 68094 11024 68100 11036
rect 68152 11024 68158 11076
rect 39724 10968 39896 10996
rect 39724 10956 39730 10968
rect 42334 10956 42340 11008
rect 42392 10956 42398 11008
rect 1104 10906 18952 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 14246 10906
rect 14298 10854 14310 10906
rect 14362 10854 14374 10906
rect 14426 10854 14438 10906
rect 14490 10854 18952 10906
rect 1104 10832 18952 10854
rect 37628 10906 68816 10928
rect 37628 10854 44246 10906
rect 44298 10854 44310 10906
rect 44362 10854 44374 10906
rect 44426 10854 44438 10906
rect 44490 10854 54246 10906
rect 54298 10854 54310 10906
rect 54362 10854 54374 10906
rect 54426 10854 54438 10906
rect 54490 10854 64246 10906
rect 64298 10854 64310 10906
rect 64362 10854 64374 10906
rect 64426 10854 64438 10906
rect 64490 10854 68816 10906
rect 37628 10832 68816 10854
rect 17494 10792 17500 10804
rect 17455 10764 17500 10792
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 18230 10792 18236 10804
rect 18191 10764 18236 10792
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 10045 10727 10103 10733
rect 10045 10693 10057 10727
rect 10091 10724 10103 10727
rect 14458 10724 14464 10736
rect 10091 10696 14464 10724
rect 10091 10693 10103 10696
rect 10045 10687 10103 10693
rect 14458 10684 14464 10696
rect 14516 10684 14522 10736
rect 51350 10724 51356 10736
rect 51046 10696 51356 10724
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4798 10656 4804 10668
rect 4387 10628 4804 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4798 10616 4804 10628
rect 4856 10656 4862 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4856 10628 4905 10656
rect 4856 10616 4862 10628
rect 4893 10625 4905 10628
rect 4939 10656 4951 10659
rect 12250 10656 12256 10668
rect 4939 10628 12256 10656
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 43990 10616 43996 10668
rect 44048 10656 44054 10668
rect 45741 10659 45799 10665
rect 45741 10656 45753 10659
rect 44048 10628 45753 10656
rect 44048 10616 44054 10628
rect 45741 10625 45753 10628
rect 45787 10656 45799 10659
rect 51046 10656 51074 10696
rect 51350 10684 51356 10696
rect 51408 10684 51414 10736
rect 45787 10628 51074 10656
rect 45787 10625 45799 10628
rect 45741 10619 45799 10625
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10588 10655 10591
rect 17218 10588 17224 10600
rect 10643 10560 17224 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 37366 10548 37372 10600
rect 37424 10588 37430 10600
rect 37734 10588 37740 10600
rect 37424 10560 37740 10588
rect 37424 10548 37430 10560
rect 37734 10548 37740 10560
rect 37792 10588 37798 10600
rect 37921 10591 37979 10597
rect 37921 10588 37933 10591
rect 37792 10560 37933 10588
rect 37792 10548 37798 10560
rect 37921 10557 37933 10560
rect 37967 10557 37979 10591
rect 37921 10551 37979 10557
rect 38010 10548 38016 10600
rect 38068 10588 38074 10600
rect 38562 10588 38568 10600
rect 38068 10560 38568 10588
rect 38068 10548 38074 10560
rect 38562 10548 38568 10560
rect 38620 10548 38626 10600
rect 42518 10548 42524 10600
rect 42576 10588 42582 10600
rect 45189 10591 45247 10597
rect 45189 10588 45201 10591
rect 42576 10560 45201 10588
rect 42576 10548 42582 10560
rect 45189 10557 45201 10560
rect 45235 10557 45247 10591
rect 45189 10551 45247 10557
rect 66993 10591 67051 10597
rect 66993 10557 67005 10591
rect 67039 10588 67051 10591
rect 67450 10588 67456 10600
rect 67039 10560 67456 10588
rect 67039 10557 67051 10560
rect 66993 10551 67051 10557
rect 67450 10548 67456 10560
rect 67508 10548 67514 10600
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 9401 10523 9459 10529
rect 9401 10520 9413 10523
rect 8536 10492 9413 10520
rect 8536 10480 8542 10492
rect 9401 10489 9413 10492
rect 9447 10520 9459 10523
rect 10686 10520 10692 10532
rect 9447 10492 10692 10520
rect 9447 10489 9459 10492
rect 9401 10483 9459 10489
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 12253 10523 12311 10529
rect 12253 10520 12265 10523
rect 11388 10492 12265 10520
rect 11388 10480 11394 10492
rect 12253 10489 12265 10492
rect 12299 10489 12311 10523
rect 12253 10483 12311 10489
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 15194 10520 15200 10532
rect 13136 10492 15200 10520
rect 13136 10480 13142 10492
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 39117 10523 39175 10529
rect 39117 10520 39129 10523
rect 37936 10492 39129 10520
rect 37936 10464 37964 10492
rect 39117 10489 39129 10492
rect 39163 10489 39175 10523
rect 39117 10483 39175 10489
rect 44818 10480 44824 10532
rect 44876 10520 44882 10532
rect 45002 10520 45008 10532
rect 44876 10492 45008 10520
rect 44876 10480 44882 10492
rect 45002 10480 45008 10492
rect 45060 10520 45066 10532
rect 46293 10523 46351 10529
rect 46293 10520 46305 10523
rect 45060 10492 46305 10520
rect 45060 10480 45066 10492
rect 46293 10489 46305 10492
rect 46339 10489 46351 10523
rect 64138 10520 64144 10532
rect 46293 10483 46351 10489
rect 51046 10492 64144 10520
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 8846 10452 8852 10464
rect 8720 10424 8852 10452
rect 8720 10412 8726 10424
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 11146 10452 11152 10464
rect 11107 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11296 10424 11713 10452
rect 11296 10412 11302 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 13173 10455 13231 10461
rect 13173 10452 13185 10455
rect 12952 10424 13185 10452
rect 12952 10412 12958 10424
rect 13173 10421 13185 10424
rect 13219 10421 13231 10455
rect 13173 10415 13231 10421
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 13872 10424 13921 10452
rect 13872 10412 13878 10424
rect 13909 10421 13921 10424
rect 13955 10421 13967 10455
rect 14550 10452 14556 10464
rect 14511 10424 14556 10452
rect 13909 10415 13967 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15838 10452 15844 10464
rect 15335 10424 15844 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16114 10452 16120 10464
rect 16075 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 37918 10412 37924 10464
rect 37976 10412 37982 10464
rect 38562 10412 38568 10464
rect 38620 10452 38626 10464
rect 38657 10455 38715 10461
rect 38657 10452 38669 10455
rect 38620 10424 38669 10452
rect 38620 10412 38626 10424
rect 38657 10421 38669 10424
rect 38703 10421 38715 10455
rect 38657 10415 38715 10421
rect 39022 10412 39028 10464
rect 39080 10452 39086 10464
rect 39669 10455 39727 10461
rect 39669 10452 39681 10455
rect 39080 10424 39681 10452
rect 39080 10412 39086 10424
rect 39669 10421 39681 10424
rect 39715 10421 39727 10455
rect 39669 10415 39727 10421
rect 40126 10412 40132 10464
rect 40184 10452 40190 10464
rect 40221 10455 40279 10461
rect 40221 10452 40233 10455
rect 40184 10424 40233 10452
rect 40184 10412 40190 10424
rect 40221 10421 40233 10424
rect 40267 10421 40279 10455
rect 40770 10452 40776 10464
rect 40731 10424 40776 10452
rect 40221 10415 40279 10421
rect 40770 10412 40776 10424
rect 40828 10412 40834 10464
rect 41417 10455 41475 10461
rect 41417 10421 41429 10455
rect 41463 10452 41475 10455
rect 41506 10452 41512 10464
rect 41463 10424 41512 10452
rect 41463 10421 41475 10424
rect 41417 10415 41475 10421
rect 41506 10412 41512 10424
rect 41564 10412 41570 10464
rect 41874 10452 41880 10464
rect 41835 10424 41880 10452
rect 41874 10412 41880 10424
rect 41932 10412 41938 10464
rect 42978 10452 42984 10464
rect 42939 10424 42984 10452
rect 42978 10412 42984 10424
rect 43036 10412 43042 10464
rect 43530 10452 43536 10464
rect 43491 10424 43536 10452
rect 43530 10412 43536 10424
rect 43588 10412 43594 10464
rect 44174 10452 44180 10464
rect 44135 10424 44180 10452
rect 44174 10412 44180 10424
rect 44232 10412 44238 10464
rect 44729 10455 44787 10461
rect 44729 10421 44741 10455
rect 44775 10452 44787 10455
rect 45094 10452 45100 10464
rect 44775 10424 45100 10452
rect 44775 10421 44787 10424
rect 44729 10415 44787 10421
rect 45094 10412 45100 10424
rect 45152 10412 45158 10464
rect 46474 10412 46480 10464
rect 46532 10452 46538 10464
rect 46937 10455 46995 10461
rect 46937 10452 46949 10455
rect 46532 10424 46949 10452
rect 46532 10412 46538 10424
rect 46937 10421 46949 10424
rect 46983 10421 46995 10455
rect 46937 10415 46995 10421
rect 47489 10455 47547 10461
rect 47489 10421 47501 10455
rect 47535 10452 47547 10455
rect 47670 10452 47676 10464
rect 47535 10424 47676 10452
rect 47535 10421 47547 10424
rect 47489 10415 47547 10421
rect 47670 10412 47676 10424
rect 47728 10452 47734 10464
rect 51046 10452 51074 10492
rect 64138 10480 64144 10492
rect 64196 10480 64202 10532
rect 66162 10520 66168 10532
rect 66075 10492 66168 10520
rect 66162 10480 66168 10492
rect 66220 10520 66226 10532
rect 67542 10520 67548 10532
rect 66220 10492 67548 10520
rect 66220 10480 66226 10492
rect 67542 10480 67548 10492
rect 67600 10480 67606 10532
rect 47728 10424 51074 10452
rect 47728 10412 47734 10424
rect 64690 10412 64696 10464
rect 64748 10452 64754 10464
rect 64785 10455 64843 10461
rect 64785 10452 64797 10455
rect 64748 10424 64797 10452
rect 64748 10412 64754 10424
rect 64785 10421 64797 10424
rect 64831 10452 64843 10455
rect 64874 10452 64880 10464
rect 64831 10424 64880 10452
rect 64831 10421 64843 10424
rect 64785 10415 64843 10421
rect 64874 10412 64880 10424
rect 64932 10412 64938 10464
rect 65518 10412 65524 10464
rect 65576 10452 65582 10464
rect 65613 10455 65671 10461
rect 65613 10452 65625 10455
rect 65576 10424 65625 10452
rect 65576 10412 65582 10424
rect 65613 10421 65625 10424
rect 65659 10452 65671 10455
rect 65702 10452 65708 10464
rect 65659 10424 65708 10452
rect 65659 10421 65671 10424
rect 65613 10415 65671 10421
rect 65702 10412 65708 10424
rect 65760 10412 65766 10464
rect 67174 10412 67180 10464
rect 67232 10452 67238 10464
rect 67453 10455 67511 10461
rect 67453 10452 67465 10455
rect 67232 10424 67465 10452
rect 67232 10412 67238 10424
rect 67453 10421 67465 10424
rect 67499 10421 67511 10455
rect 68002 10452 68008 10464
rect 67963 10424 68008 10452
rect 67453 10415 67511 10421
rect 68002 10412 68008 10424
rect 68060 10412 68066 10464
rect 1104 10362 18952 10384
rect 1104 10310 9246 10362
rect 9298 10310 9310 10362
rect 9362 10310 9374 10362
rect 9426 10310 9438 10362
rect 9490 10310 18952 10362
rect 1104 10288 18952 10310
rect 37628 10362 68816 10384
rect 37628 10310 39246 10362
rect 39298 10310 39310 10362
rect 39362 10310 39374 10362
rect 39426 10310 39438 10362
rect 39490 10310 49246 10362
rect 49298 10310 49310 10362
rect 49362 10310 49374 10362
rect 49426 10310 49438 10362
rect 49490 10310 59246 10362
rect 59298 10310 59310 10362
rect 59362 10310 59374 10362
rect 59426 10310 59438 10362
rect 59490 10310 68816 10362
rect 37628 10288 68816 10310
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 2406 10248 2412 10260
rect 2271 10220 2412 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 9217 10251 9275 10257
rect 9217 10217 9229 10251
rect 9263 10248 9275 10251
rect 14090 10248 14096 10260
rect 9263 10220 14096 10248
rect 9263 10217 9275 10220
rect 9217 10211 9275 10217
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 15286 10248 15292 10260
rect 14660 10220 15292 10248
rect 13817 10183 13875 10189
rect 13817 10149 13829 10183
rect 13863 10180 13875 10183
rect 14660 10180 14688 10220
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 45741 10251 45799 10257
rect 45741 10248 45753 10251
rect 41386 10220 45753 10248
rect 13863 10152 14688 10180
rect 14737 10183 14795 10189
rect 13863 10149 13875 10152
rect 13817 10143 13875 10149
rect 14737 10149 14749 10183
rect 14783 10180 14795 10183
rect 16206 10180 16212 10192
rect 14783 10152 16212 10180
rect 14783 10149 14795 10152
rect 14737 10143 14795 10149
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 39390 10140 39396 10192
rect 39448 10180 39454 10192
rect 39666 10180 39672 10192
rect 39448 10152 39672 10180
rect 39448 10140 39454 10152
rect 39666 10140 39672 10152
rect 39724 10140 39730 10192
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 14458 10112 14464 10124
rect 12584 10084 14464 10112
rect 12584 10072 12590 10084
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 15194 10112 15200 10124
rect 15155 10084 15200 10112
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10112 18291 10115
rect 18322 10112 18328 10124
rect 18279 10084 18328 10112
rect 18279 10081 18291 10084
rect 18233 10075 18291 10081
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 32674 10072 32680 10124
rect 32732 10112 32738 10124
rect 37826 10112 37832 10124
rect 32732 10084 37832 10112
rect 32732 10072 32738 10084
rect 37826 10072 37832 10084
rect 37884 10112 37890 10124
rect 37921 10115 37979 10121
rect 37921 10112 37933 10115
rect 37884 10084 37933 10112
rect 37884 10072 37890 10084
rect 37921 10081 37933 10084
rect 37967 10081 37979 10115
rect 37921 10075 37979 10081
rect 38565 10115 38623 10121
rect 38565 10081 38577 10115
rect 38611 10081 38623 10115
rect 38565 10075 38623 10081
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 11606 10044 11612 10056
rect 8067 10016 11612 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 36078 10004 36084 10056
rect 36136 10044 36142 10056
rect 37182 10044 37188 10056
rect 36136 10016 37188 10044
rect 36136 10004 36142 10016
rect 37182 10004 37188 10016
rect 37240 10044 37246 10056
rect 38580 10044 38608 10075
rect 41386 10044 41414 10220
rect 45741 10217 45753 10220
rect 45787 10248 45799 10251
rect 47026 10248 47032 10260
rect 45787 10220 47032 10248
rect 45787 10217 45799 10220
rect 45741 10211 45799 10217
rect 47026 10208 47032 10220
rect 47084 10208 47090 10260
rect 45094 10140 45100 10192
rect 45152 10180 45158 10192
rect 64966 10180 64972 10192
rect 45152 10152 64972 10180
rect 45152 10140 45158 10152
rect 64966 10140 64972 10152
rect 65024 10140 65030 10192
rect 67634 10140 67640 10192
rect 67692 10180 67698 10192
rect 67913 10183 67971 10189
rect 67913 10180 67925 10183
rect 67692 10152 67925 10180
rect 67692 10140 67698 10152
rect 67913 10149 67925 10152
rect 67959 10149 67971 10183
rect 67913 10143 67971 10149
rect 44082 10112 44088 10124
rect 44043 10084 44088 10112
rect 44082 10072 44088 10084
rect 44140 10072 44146 10124
rect 63770 10072 63776 10124
rect 63828 10112 63834 10124
rect 63954 10112 63960 10124
rect 63828 10084 63960 10112
rect 63828 10072 63834 10084
rect 63954 10072 63960 10084
rect 64012 10072 64018 10124
rect 37240 10016 38608 10044
rect 38672 10016 41414 10044
rect 37240 10004 37246 10016
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 12989 9979 13047 9985
rect 12989 9976 13001 9979
rect 12584 9948 13001 9976
rect 12584 9936 12590 9948
rect 12989 9945 13001 9948
rect 13035 9945 13047 9979
rect 12989 9939 13047 9945
rect 17037 9979 17095 9985
rect 17037 9945 17049 9979
rect 17083 9976 17095 9979
rect 18322 9976 18328 9988
rect 17083 9948 18328 9976
rect 17083 9945 17095 9948
rect 17037 9939 17095 9945
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 38286 9936 38292 9988
rect 38344 9976 38350 9988
rect 38672 9976 38700 10016
rect 41690 10004 41696 10056
rect 41748 10044 41754 10056
rect 42518 10044 42524 10056
rect 41748 10016 42524 10044
rect 41748 10004 41754 10016
rect 42518 10004 42524 10016
rect 42576 10004 42582 10056
rect 44910 10004 44916 10056
rect 44968 10004 44974 10056
rect 41230 9976 41236 9988
rect 38344 9948 38700 9976
rect 39224 9948 41236 9976
rect 38344 9936 38350 9948
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2832 9880 2877 9908
rect 2832 9868 2838 9880
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 3878 9908 3884 9920
rect 3752 9880 3884 9908
rect 3752 9868 3758 9880
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 5353 9911 5411 9917
rect 5353 9908 5365 9911
rect 5224 9880 5365 9908
rect 5224 9868 5230 9880
rect 5353 9877 5365 9880
rect 5399 9908 5411 9911
rect 5442 9908 5448 9920
rect 5399 9880 5448 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 6549 9911 6607 9917
rect 6549 9908 6561 9911
rect 6420 9880 6561 9908
rect 6420 9868 6426 9880
rect 6549 9877 6561 9880
rect 6595 9908 6607 9911
rect 6730 9908 6736 9920
rect 6595 9880 6736 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 7190 9908 7196 9920
rect 7151 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 8570 9908 8576 9920
rect 8531 9880 8576 9908
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 9766 9908 9772 9920
rect 9727 9880 9772 9908
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10226 9868 10232 9920
rect 10284 9908 10290 9920
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10284 9880 10333 9908
rect 10284 9868 10290 9880
rect 10321 9877 10333 9880
rect 10367 9877 10379 9911
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 10321 9871 10379 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 11885 9911 11943 9917
rect 11885 9908 11897 9911
rect 11664 9880 11897 9908
rect 11664 9868 11670 9880
rect 11885 9877 11897 9880
rect 11931 9877 11943 9911
rect 11885 9871 11943 9877
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12492 9880 12537 9908
rect 12492 9868 12498 9880
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 15841 9911 15899 9917
rect 15841 9908 15853 9911
rect 15620 9880 15853 9908
rect 15620 9868 15626 9880
rect 15841 9877 15853 9880
rect 15887 9877 15899 9911
rect 15841 9871 15899 9877
rect 16485 9911 16543 9917
rect 16485 9877 16497 9911
rect 16531 9908 16543 9911
rect 16574 9908 16580 9920
rect 16531 9880 16580 9908
rect 16531 9877 16543 9880
rect 16485 9871 16543 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 17589 9911 17647 9917
rect 17589 9877 17601 9911
rect 17635 9908 17647 9911
rect 18138 9908 18144 9920
rect 17635 9880 18144 9908
rect 17635 9877 17647 9880
rect 17589 9871 17647 9877
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 32582 9868 32588 9920
rect 32640 9908 32646 9920
rect 39224 9917 39252 9948
rect 41230 9936 41236 9948
rect 41288 9936 41294 9988
rect 44928 9976 44956 10004
rect 45278 9976 45284 9988
rect 44928 9948 45284 9976
rect 45278 9936 45284 9948
rect 45336 9976 45342 9988
rect 47305 9979 47363 9985
rect 47305 9976 47317 9979
rect 45336 9948 47317 9976
rect 45336 9936 45342 9948
rect 47305 9945 47317 9948
rect 47351 9945 47363 9979
rect 47305 9939 47363 9945
rect 65794 9936 65800 9988
rect 65852 9976 65858 9988
rect 66073 9979 66131 9985
rect 66073 9976 66085 9979
rect 65852 9948 66085 9976
rect 65852 9936 65858 9948
rect 66073 9945 66085 9948
rect 66119 9976 66131 9979
rect 66898 9976 66904 9988
rect 66119 9948 66904 9976
rect 66119 9945 66131 9948
rect 66073 9939 66131 9945
rect 66898 9936 66904 9948
rect 66956 9936 66962 9988
rect 68094 9976 68100 9988
rect 68055 9948 68100 9976
rect 68094 9936 68100 9948
rect 68152 9936 68158 9988
rect 39209 9911 39267 9917
rect 39209 9908 39221 9911
rect 32640 9880 39221 9908
rect 32640 9868 32646 9880
rect 39209 9877 39221 9880
rect 39255 9877 39267 9911
rect 39209 9871 39267 9877
rect 39482 9868 39488 9920
rect 39540 9908 39546 9920
rect 39761 9911 39819 9917
rect 39761 9908 39773 9911
rect 39540 9880 39773 9908
rect 39540 9868 39546 9880
rect 39761 9877 39773 9880
rect 39807 9877 39819 9911
rect 39761 9871 39819 9877
rect 40589 9911 40647 9917
rect 40589 9877 40601 9911
rect 40635 9908 40647 9911
rect 40862 9908 40868 9920
rect 40635 9880 40868 9908
rect 40635 9877 40647 9880
rect 40589 9871 40647 9877
rect 40862 9868 40868 9880
rect 40920 9868 40926 9920
rect 41138 9908 41144 9920
rect 41099 9880 41144 9908
rect 41138 9868 41144 9880
rect 41196 9868 41202 9920
rect 41690 9908 41696 9920
rect 41651 9880 41696 9908
rect 41690 9868 41696 9880
rect 41748 9868 41754 9920
rect 42150 9868 42156 9920
rect 42208 9908 42214 9920
rect 42245 9911 42303 9917
rect 42245 9908 42257 9911
rect 42208 9880 42257 9908
rect 42208 9868 42214 9880
rect 42245 9877 42257 9880
rect 42291 9877 42303 9911
rect 42794 9908 42800 9920
rect 42755 9880 42800 9908
rect 42245 9871 42303 9877
rect 42794 9868 42800 9880
rect 42852 9868 42858 9920
rect 43346 9908 43352 9920
rect 43307 9880 43352 9908
rect 43346 9868 43352 9880
rect 43404 9868 43410 9920
rect 44821 9911 44879 9917
rect 44821 9877 44833 9911
rect 44867 9908 44879 9911
rect 44910 9908 44916 9920
rect 44867 9880 44916 9908
rect 44867 9877 44879 9880
rect 44821 9871 44879 9877
rect 44910 9868 44916 9880
rect 44968 9868 44974 9920
rect 46290 9908 46296 9920
rect 46251 9880 46296 9908
rect 46290 9868 46296 9880
rect 46348 9868 46354 9920
rect 46750 9908 46756 9920
rect 46711 9880 46756 9908
rect 46750 9868 46756 9880
rect 46808 9868 46814 9920
rect 47762 9868 47768 9920
rect 47820 9908 47826 9920
rect 47857 9911 47915 9917
rect 47857 9908 47869 9911
rect 47820 9880 47869 9908
rect 47820 9868 47826 9880
rect 47857 9877 47869 9880
rect 47903 9877 47915 9911
rect 63954 9908 63960 9920
rect 63915 9880 63960 9908
rect 47857 9871 47915 9877
rect 63954 9868 63960 9880
rect 64012 9868 64018 9920
rect 64877 9911 64935 9917
rect 64877 9877 64889 9911
rect 64923 9908 64935 9911
rect 64966 9908 64972 9920
rect 64923 9880 64972 9908
rect 64923 9877 64935 9880
rect 64877 9871 64935 9877
rect 64966 9868 64972 9880
rect 65024 9868 65030 9920
rect 65429 9911 65487 9917
rect 65429 9877 65441 9911
rect 65475 9908 65487 9911
rect 65886 9908 65892 9920
rect 65475 9880 65892 9908
rect 65475 9877 65487 9880
rect 65429 9871 65487 9877
rect 65886 9868 65892 9880
rect 65944 9868 65950 9920
rect 66990 9908 66996 9920
rect 66951 9880 66996 9908
rect 66990 9868 66996 9880
rect 67048 9868 67054 9920
rect 1104 9818 18952 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 14246 9818
rect 14298 9766 14310 9818
rect 14362 9766 14374 9818
rect 14426 9766 14438 9818
rect 14490 9766 18952 9818
rect 1104 9744 18952 9766
rect 37628 9818 68816 9840
rect 37628 9766 44246 9818
rect 44298 9766 44310 9818
rect 44362 9766 44374 9818
rect 44426 9766 44438 9818
rect 44490 9766 54246 9818
rect 54298 9766 54310 9818
rect 54362 9766 54374 9818
rect 54426 9766 54438 9818
rect 54490 9766 64246 9818
rect 64298 9766 64310 9818
rect 64362 9766 64374 9818
rect 64426 9766 64438 9818
rect 64490 9766 68816 9818
rect 37628 9744 68816 9766
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 13078 9704 13084 9716
rect 6604 9676 13084 9704
rect 6604 9664 6610 9676
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 14826 9664 14832 9716
rect 14884 9704 14890 9716
rect 15194 9704 15200 9716
rect 14884 9676 15200 9704
rect 14884 9664 14890 9676
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 39758 9664 39764 9716
rect 39816 9704 39822 9716
rect 41322 9704 41328 9716
rect 39816 9676 41328 9704
rect 39816 9664 39822 9676
rect 41322 9664 41328 9676
rect 41380 9664 41386 9716
rect 1762 9636 1768 9648
rect 1723 9608 1768 9636
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 2590 9636 2596 9648
rect 2551 9608 2596 9636
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 5074 9636 5080 9648
rect 4571 9608 5080 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 4540 9568 4568 9599
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 18049 9639 18107 9645
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 18874 9636 18880 9648
rect 18095 9608 18880 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 18874 9596 18880 9608
rect 18932 9596 18938 9648
rect 37734 9596 37740 9648
rect 37792 9636 37798 9648
rect 38010 9636 38016 9648
rect 37792 9608 38016 9636
rect 37792 9596 37798 9608
rect 38010 9596 38016 9608
rect 38068 9596 38074 9648
rect 3896 9540 4568 9568
rect 10597 9571 10655 9577
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2406 9500 2412 9512
rect 1995 9472 2412 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 3717 9503 3775 9509
rect 3717 9469 3729 9503
rect 3763 9500 3775 9503
rect 3896 9500 3924 9540
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 23934 9568 23940 9580
rect 10643 9540 23940 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 23934 9528 23940 9540
rect 23992 9528 23998 9580
rect 34057 9571 34115 9577
rect 34057 9537 34069 9571
rect 34103 9568 34115 9571
rect 34103 9540 39252 9568
rect 34103 9537 34115 9540
rect 34057 9531 34115 9537
rect 3763 9472 3924 9500
rect 3973 9503 4031 9509
rect 3763 9469 3775 9472
rect 3717 9463 3775 9469
rect 3973 9469 3985 9503
rect 4019 9500 4031 9503
rect 4154 9500 4160 9512
rect 4019 9472 4160 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 4154 9460 4160 9472
rect 4212 9500 4218 9512
rect 4798 9500 4804 9512
rect 4212 9472 4804 9500
rect 4212 9460 4218 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5626 9500 5632 9512
rect 5539 9472 5632 9500
rect 5626 9460 5632 9472
rect 5684 9500 5690 9512
rect 5810 9500 5816 9512
rect 5684 9472 5816 9500
rect 5684 9460 5690 9472
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 6880 9472 8953 9500
rect 6880 9460 6886 9472
rect 8941 9469 8953 9472
rect 8987 9500 8999 9503
rect 9674 9500 9680 9512
rect 8987 9472 9680 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11974 9500 11980 9512
rect 11195 9472 11980 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13872 9472 14013 9500
rect 13872 9460 13878 9472
rect 14001 9469 14013 9472
rect 14047 9500 14059 9503
rect 14918 9500 14924 9512
rect 14047 9472 14924 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 15470 9500 15476 9512
rect 15252 9472 15476 9500
rect 15252 9460 15258 9472
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9500 16451 9503
rect 17494 9500 17500 9512
rect 16439 9472 17500 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9469 17647 9503
rect 17589 9463 17647 9469
rect 7377 9435 7435 9441
rect 7377 9401 7389 9435
rect 7423 9432 7435 9435
rect 13630 9432 13636 9444
rect 7423 9404 13636 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 13630 9392 13636 9404
rect 13688 9392 13694 9444
rect 15289 9435 15347 9441
rect 15289 9401 15301 9435
rect 15335 9432 15347 9435
rect 17604 9432 17632 9463
rect 37274 9460 37280 9512
rect 37332 9500 37338 9512
rect 37921 9503 37979 9509
rect 37921 9500 37933 9503
rect 37332 9472 37933 9500
rect 37332 9460 37338 9472
rect 37921 9469 37933 9472
rect 37967 9469 37979 9503
rect 37921 9463 37979 9469
rect 38749 9503 38807 9509
rect 38749 9469 38761 9503
rect 38795 9500 38807 9503
rect 39114 9500 39120 9512
rect 38795 9472 39120 9500
rect 38795 9469 38807 9472
rect 38749 9463 38807 9469
rect 23842 9432 23848 9444
rect 15335 9404 17540 9432
rect 17604 9404 23848 9432
rect 15335 9401 15347 9404
rect 15289 9395 15347 9401
rect 4982 9324 4988 9376
rect 5040 9364 5046 9376
rect 5077 9367 5135 9373
rect 5077 9364 5089 9367
rect 5040 9336 5089 9364
rect 5040 9324 5046 9336
rect 5077 9333 5089 9336
rect 5123 9364 5135 9367
rect 5258 9364 5264 9376
rect 5123 9336 5264 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 5684 9336 6469 9364
rect 5684 9324 5690 9336
rect 6457 9333 6469 9336
rect 6503 9364 6515 9367
rect 6638 9364 6644 9376
rect 6503 9336 6644 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7834 9364 7840 9376
rect 7795 9336 7840 9364
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 8444 9336 8493 9364
rect 8444 9324 8450 9336
rect 8481 9333 8493 9336
rect 8527 9364 8539 9367
rect 8754 9364 8760 9376
rect 8527 9336 8760 9364
rect 8527 9333 8539 9336
rect 8481 9327 8539 9333
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 12066 9364 12072 9376
rect 12027 9336 12072 9364
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13170 9364 13176 9376
rect 12851 9336 13176 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13354 9364 13360 9376
rect 13315 9336 13360 9364
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 14737 9367 14795 9373
rect 14737 9333 14749 9367
rect 14783 9364 14795 9367
rect 15470 9364 15476 9376
rect 14783 9336 15476 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 16206 9364 16212 9376
rect 15887 9336 16212 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 17512 9364 17540 9404
rect 23842 9392 23848 9404
rect 23900 9392 23906 9444
rect 31481 9435 31539 9441
rect 31481 9401 31493 9435
rect 31527 9432 31539 9435
rect 38764 9432 38792 9463
rect 39114 9460 39120 9472
rect 39172 9460 39178 9512
rect 39224 9500 39252 9540
rect 43898 9528 43904 9580
rect 43956 9568 43962 9580
rect 44082 9568 44088 9580
rect 43956 9540 44088 9568
rect 43956 9528 43962 9540
rect 44082 9528 44088 9540
rect 44140 9568 44146 9580
rect 47581 9571 47639 9577
rect 47581 9568 47593 9571
rect 44140 9540 47593 9568
rect 44140 9528 44146 9540
rect 47581 9537 47593 9540
rect 47627 9537 47639 9571
rect 47581 9531 47639 9537
rect 39390 9500 39396 9512
rect 39224 9472 39396 9500
rect 39390 9460 39396 9472
rect 39448 9460 39454 9512
rect 40037 9503 40095 9509
rect 40037 9469 40049 9503
rect 40083 9500 40095 9503
rect 40310 9500 40316 9512
rect 40083 9472 40316 9500
rect 40083 9469 40095 9472
rect 40037 9463 40095 9469
rect 31527 9404 38792 9432
rect 31527 9401 31539 9404
rect 31481 9395 31539 9401
rect 18230 9364 18236 9376
rect 17512 9336 18236 9364
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 38010 9324 38016 9376
rect 38068 9364 38074 9376
rect 40052 9364 40080 9463
rect 40310 9460 40316 9472
rect 40368 9460 40374 9512
rect 40957 9503 41015 9509
rect 40957 9469 40969 9503
rect 41003 9500 41015 9503
rect 41230 9500 41236 9512
rect 41003 9472 41236 9500
rect 41003 9469 41015 9472
rect 40957 9463 41015 9469
rect 41230 9460 41236 9472
rect 41288 9500 41294 9512
rect 42058 9500 42064 9512
rect 41288 9472 42064 9500
rect 41288 9460 41294 9472
rect 42058 9460 42064 9472
rect 42116 9460 42122 9512
rect 43073 9503 43131 9509
rect 43073 9469 43085 9503
rect 43119 9500 43131 9503
rect 43162 9500 43168 9512
rect 43119 9472 43168 9500
rect 43119 9469 43131 9472
rect 43073 9463 43131 9469
rect 43162 9460 43168 9472
rect 43220 9460 43226 9512
rect 45370 9460 45376 9512
rect 45428 9500 45434 9512
rect 45428 9472 63632 9500
rect 45428 9460 45434 9472
rect 44177 9435 44235 9441
rect 44177 9401 44189 9435
rect 44223 9432 44235 9435
rect 44818 9432 44824 9444
rect 44223 9404 44824 9432
rect 44223 9401 44235 9404
rect 44177 9395 44235 9401
rect 44818 9392 44824 9404
rect 44876 9392 44882 9444
rect 46014 9392 46020 9444
rect 46072 9432 46078 9444
rect 46382 9432 46388 9444
rect 46072 9404 46388 9432
rect 46072 9392 46078 9404
rect 46382 9392 46388 9404
rect 46440 9432 46446 9444
rect 47029 9435 47087 9441
rect 47029 9432 47041 9435
rect 46440 9404 47041 9432
rect 46440 9392 46446 9404
rect 47029 9401 47041 9404
rect 47075 9401 47087 9435
rect 47029 9395 47087 9401
rect 48590 9392 48596 9444
rect 48648 9432 48654 9444
rect 48685 9435 48743 9441
rect 48685 9432 48697 9435
rect 48648 9404 48697 9432
rect 48648 9392 48654 9404
rect 48685 9401 48697 9404
rect 48731 9432 48743 9435
rect 48866 9432 48872 9444
rect 48731 9404 48872 9432
rect 48731 9401 48743 9404
rect 48685 9395 48743 9401
rect 48866 9392 48872 9404
rect 48924 9392 48930 9444
rect 60458 9432 60464 9444
rect 49712 9404 60464 9432
rect 38068 9336 40080 9364
rect 38068 9324 38074 9336
rect 40310 9324 40316 9376
rect 40368 9364 40374 9376
rect 40494 9364 40500 9376
rect 40368 9336 40500 9364
rect 40368 9324 40374 9336
rect 40494 9324 40500 9336
rect 40552 9324 40558 9376
rect 41509 9367 41567 9373
rect 41509 9333 41521 9367
rect 41555 9364 41567 9367
rect 41598 9364 41604 9376
rect 41555 9336 41604 9364
rect 41555 9333 41567 9336
rect 41509 9327 41567 9333
rect 41598 9324 41604 9336
rect 41656 9324 41662 9376
rect 42058 9364 42064 9376
rect 42019 9336 42064 9364
rect 42058 9324 42064 9336
rect 42116 9324 42122 9376
rect 43070 9324 43076 9376
rect 43128 9364 43134 9376
rect 43533 9367 43591 9373
rect 43533 9364 43545 9367
rect 43128 9336 43545 9364
rect 43128 9324 43134 9336
rect 43533 9333 43545 9336
rect 43579 9333 43591 9367
rect 44726 9364 44732 9376
rect 44687 9336 44732 9364
rect 43533 9327 43591 9333
rect 44726 9324 44732 9336
rect 44784 9324 44790 9376
rect 45186 9364 45192 9376
rect 45147 9336 45192 9364
rect 45186 9324 45192 9336
rect 45244 9324 45250 9376
rect 45830 9364 45836 9376
rect 45791 9336 45836 9364
rect 45830 9324 45836 9336
rect 45888 9324 45894 9376
rect 46566 9364 46572 9376
rect 46527 9336 46572 9364
rect 46566 9324 46572 9336
rect 46624 9324 46630 9376
rect 48774 9324 48780 9376
rect 48832 9364 48838 9376
rect 49142 9364 49148 9376
rect 48832 9336 49148 9364
rect 48832 9324 48838 9336
rect 49142 9324 49148 9336
rect 49200 9324 49206 9376
rect 49602 9324 49608 9376
rect 49660 9364 49666 9376
rect 49712 9373 49740 9404
rect 60458 9392 60464 9404
rect 60516 9392 60522 9444
rect 63604 9376 63632 9472
rect 65705 9435 65763 9441
rect 65705 9401 65717 9435
rect 65751 9432 65763 9435
rect 68094 9432 68100 9444
rect 65751 9404 68100 9432
rect 65751 9401 65763 9404
rect 65705 9395 65763 9401
rect 68094 9392 68100 9404
rect 68152 9392 68158 9444
rect 49697 9367 49755 9373
rect 49697 9364 49709 9367
rect 49660 9336 49709 9364
rect 49660 9324 49666 9336
rect 49697 9333 49709 9336
rect 49743 9333 49755 9367
rect 50246 9364 50252 9376
rect 50207 9336 50252 9364
rect 49697 9327 49755 9333
rect 50246 9324 50252 9336
rect 50304 9324 50310 9376
rect 62666 9324 62672 9376
rect 62724 9364 62730 9376
rect 63310 9364 63316 9376
rect 62724 9336 63316 9364
rect 62724 9324 62730 9336
rect 63310 9324 63316 9336
rect 63368 9324 63374 9376
rect 63586 9324 63592 9376
rect 63644 9364 63650 9376
rect 63957 9367 64015 9373
rect 63957 9364 63969 9367
rect 63644 9336 63969 9364
rect 63644 9324 63650 9336
rect 63957 9333 63969 9336
rect 64003 9333 64015 9367
rect 63957 9327 64015 9333
rect 64230 9324 64236 9376
rect 64288 9364 64294 9376
rect 64509 9367 64567 9373
rect 64509 9364 64521 9367
rect 64288 9336 64521 9364
rect 64288 9324 64294 9336
rect 64509 9333 64521 9336
rect 64555 9333 64567 9367
rect 64509 9327 64567 9333
rect 65153 9367 65211 9373
rect 65153 9333 65165 9367
rect 65199 9364 65211 9367
rect 65242 9364 65248 9376
rect 65199 9336 65248 9364
rect 65199 9333 65211 9336
rect 65153 9327 65211 9333
rect 65242 9324 65248 9336
rect 65300 9324 65306 9376
rect 65978 9324 65984 9376
rect 66036 9364 66042 9376
rect 66257 9367 66315 9373
rect 66257 9364 66269 9367
rect 66036 9336 66269 9364
rect 66036 9324 66042 9336
rect 66257 9333 66269 9336
rect 66303 9333 66315 9367
rect 66714 9364 66720 9376
rect 66675 9336 66720 9364
rect 66257 9327 66315 9333
rect 66714 9324 66720 9336
rect 66772 9324 66778 9376
rect 67266 9324 67272 9376
rect 67324 9364 67330 9376
rect 67637 9367 67695 9373
rect 67637 9364 67649 9367
rect 67324 9336 67649 9364
rect 67324 9324 67330 9336
rect 67637 9333 67649 9336
rect 67683 9333 67695 9367
rect 67637 9327 67695 9333
rect 1104 9274 18952 9296
rect 1104 9222 9246 9274
rect 9298 9222 9310 9274
rect 9362 9222 9374 9274
rect 9426 9222 9438 9274
rect 9490 9222 18952 9274
rect 1104 9200 18952 9222
rect 37628 9274 68816 9296
rect 37628 9222 39246 9274
rect 39298 9222 39310 9274
rect 39362 9222 39374 9274
rect 39426 9222 39438 9274
rect 39490 9222 49246 9274
rect 49298 9222 49310 9274
rect 49362 9222 49374 9274
rect 49426 9222 49438 9274
rect 49490 9222 59246 9274
rect 59298 9222 59310 9274
rect 59362 9222 59374 9274
rect 59426 9222 59438 9274
rect 59490 9222 68816 9274
rect 37628 9200 68816 9222
rect 7466 9160 7472 9172
rect 7427 9132 7472 9160
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 8754 9120 8760 9172
rect 8812 9160 8818 9172
rect 17862 9160 17868 9172
rect 8812 9132 17868 9160
rect 8812 9120 8818 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 63678 9120 63684 9172
rect 63736 9160 63742 9172
rect 64509 9163 64567 9169
rect 64509 9160 64521 9163
rect 63736 9132 64521 9160
rect 63736 9120 63742 9132
rect 64509 9129 64521 9132
rect 64555 9160 64567 9163
rect 67818 9160 67824 9172
rect 64555 9132 67824 9160
rect 64555 9129 64567 9132
rect 64509 9123 64567 9129
rect 67818 9120 67824 9132
rect 67876 9120 67882 9172
rect 50890 9092 50896 9104
rect 32324 9064 39160 9092
rect 50803 9064 50896 9092
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13504 8996 13645 9024
rect 13504 8984 13510 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 14734 9024 14740 9036
rect 14695 8996 14740 9024
rect 13633 8987 13691 8993
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 9024 15439 9027
rect 15654 9024 15660 9036
rect 15427 8996 15660 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 17586 9024 17592 9036
rect 17499 8996 17592 9024
rect 17586 8984 17592 8996
rect 17644 9024 17650 9036
rect 24946 9024 24952 9036
rect 17644 8996 24952 9024
rect 17644 8984 17650 8996
rect 24946 8984 24952 8996
rect 25004 8984 25010 9036
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 14090 8956 14096 8968
rect 12483 8928 14096 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 17218 8956 17224 8968
rect 14384 8928 17224 8956
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 4433 8891 4491 8897
rect 4433 8888 4445 8891
rect 2464 8860 4445 8888
rect 2464 8848 2470 8860
rect 4433 8857 4445 8860
rect 4479 8888 4491 8891
rect 6270 8888 6276 8900
rect 4479 8860 6276 8888
rect 4479 8857 4491 8860
rect 4433 8851 4491 8857
rect 6270 8848 6276 8860
rect 6328 8888 6334 8900
rect 7282 8888 7288 8900
rect 6328 8860 7288 8888
rect 6328 8848 6334 8860
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 11885 8891 11943 8897
rect 11885 8857 11897 8891
rect 11931 8888 11943 8891
rect 14384 8888 14412 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 32324 8900 32352 9064
rect 32766 8984 32772 9036
rect 32824 9024 32830 9036
rect 38105 9027 38163 9033
rect 38105 9024 38117 9027
rect 32824 8996 38117 9024
rect 32824 8984 32830 8996
rect 38105 8993 38117 8996
rect 38151 9024 38163 9027
rect 38194 9024 38200 9036
rect 38151 8996 38200 9024
rect 38151 8993 38163 8996
rect 38105 8987 38163 8993
rect 38194 8984 38200 8996
rect 38252 8984 38258 9036
rect 38933 9027 38991 9033
rect 38933 8993 38945 9027
rect 38979 9024 38991 9027
rect 39022 9024 39028 9036
rect 38979 8996 39028 9024
rect 38979 8993 38991 8996
rect 38933 8987 38991 8993
rect 39022 8984 39028 8996
rect 39080 8984 39086 9036
rect 39132 9024 39160 9064
rect 50890 9052 50896 9064
rect 50948 9092 50954 9104
rect 51350 9092 51356 9104
rect 50948 9064 51356 9092
rect 50948 9052 50954 9064
rect 51350 9052 51356 9064
rect 51408 9052 51414 9104
rect 39577 9027 39635 9033
rect 39577 9024 39589 9027
rect 39132 8996 39589 9024
rect 39577 8993 39589 8996
rect 39623 9024 39635 9027
rect 40494 9024 40500 9036
rect 39623 8996 40500 9024
rect 39623 8993 39635 8996
rect 39577 8987 39635 8993
rect 40494 8984 40500 8996
rect 40552 8984 40558 9036
rect 41141 9027 41199 9033
rect 41141 8993 41153 9027
rect 41187 8993 41199 9027
rect 41141 8987 41199 8993
rect 34882 8916 34888 8968
rect 34940 8956 34946 8968
rect 41046 8956 41052 8968
rect 34940 8928 41052 8956
rect 34940 8916 34946 8928
rect 41046 8916 41052 8928
rect 41104 8956 41110 8968
rect 41156 8956 41184 8987
rect 48406 8984 48412 9036
rect 48464 9024 48470 9036
rect 50338 9024 50344 9036
rect 48464 8996 50344 9024
rect 48464 8984 48470 8996
rect 50338 8984 50344 8996
rect 50396 8984 50402 9036
rect 68094 9024 68100 9036
rect 68007 8996 68100 9024
rect 68094 8984 68100 8996
rect 68152 9024 68158 9036
rect 68830 9024 68836 9036
rect 68152 8996 68836 9024
rect 68152 8984 68158 8996
rect 68830 8984 68836 8996
rect 68888 8984 68894 9036
rect 41104 8928 41184 8956
rect 41104 8916 41110 8928
rect 46842 8916 46848 8968
rect 46900 8956 46906 8968
rect 48961 8959 49019 8965
rect 48961 8956 48973 8959
rect 46900 8928 48973 8956
rect 46900 8916 46906 8928
rect 48961 8925 48973 8928
rect 49007 8925 49019 8959
rect 48961 8919 49019 8925
rect 11931 8860 14412 8888
rect 16945 8891 17003 8897
rect 11931 8857 11943 8860
rect 11885 8851 11943 8857
rect 16945 8857 16957 8891
rect 16991 8888 17003 8891
rect 19334 8888 19340 8900
rect 16991 8860 19340 8888
rect 16991 8857 17003 8860
rect 16945 8851 17003 8857
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 32306 8848 32312 8900
rect 32364 8848 32370 8900
rect 37734 8848 37740 8900
rect 37792 8888 37798 8900
rect 61378 8888 61384 8900
rect 37792 8860 61384 8888
rect 37792 8848 37798 8860
rect 61378 8848 61384 8860
rect 61436 8848 61442 8900
rect 62298 8848 62304 8900
rect 62356 8888 62362 8900
rect 62393 8891 62451 8897
rect 62393 8888 62405 8891
rect 62356 8860 62405 8888
rect 62356 8848 62362 8860
rect 62393 8857 62405 8860
rect 62439 8888 62451 8891
rect 65518 8888 65524 8900
rect 62439 8860 65524 8888
rect 62439 8857 62451 8860
rect 62393 8851 62451 8857
rect 65518 8848 65524 8860
rect 65576 8848 65582 8900
rect 66901 8891 66959 8897
rect 66901 8857 66913 8891
rect 66947 8888 66959 8891
rect 67726 8888 67732 8900
rect 66947 8860 67732 8888
rect 66947 8857 66959 8860
rect 66901 8851 66959 8857
rect 67726 8848 67732 8860
rect 67784 8848 67790 8900
rect 1394 8820 1400 8832
rect 1355 8792 1400 8820
rect 1394 8780 1400 8792
rect 1452 8780 1458 8832
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 1949 8823 2007 8829
rect 1949 8820 1961 8823
rect 1728 8792 1961 8820
rect 1728 8780 1734 8792
rect 1949 8789 1961 8792
rect 1995 8789 2007 8823
rect 2498 8820 2504 8832
rect 2459 8792 2504 8820
rect 1949 8783 2007 8789
rect 2498 8780 2504 8792
rect 2556 8780 2562 8832
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3016 8792 3249 8820
rect 3016 8780 3022 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3970 8820 3976 8832
rect 3931 8792 3976 8820
rect 3237 8783 3295 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 5350 8820 5356 8832
rect 5311 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 6086 8820 6092 8832
rect 5960 8792 6092 8820
rect 5960 8780 5966 8792
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 7009 8823 7067 8829
rect 7009 8789 7021 8823
rect 7055 8820 7067 8823
rect 7098 8820 7104 8832
rect 7055 8792 7104 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 8294 8820 8300 8832
rect 8255 8792 8300 8820
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8904 8792 9137 8820
rect 8904 8780 8910 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 9125 8783 9183 8789
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 11149 8823 11207 8829
rect 11149 8820 11161 8823
rect 11112 8792 11161 8820
rect 11112 8780 11118 8792
rect 11149 8789 11161 8792
rect 11195 8789 11207 8823
rect 11149 8783 11207 8789
rect 12989 8823 13047 8829
rect 12989 8789 13001 8823
rect 13035 8820 13047 8823
rect 13538 8820 13544 8832
rect 13035 8792 13544 8820
rect 13035 8789 13047 8792
rect 12989 8783 13047 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 16393 8823 16451 8829
rect 16393 8789 16405 8823
rect 16439 8820 16451 8823
rect 16850 8820 16856 8832
rect 16439 8792 16856 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 18233 8823 18291 8829
rect 18233 8789 18245 8823
rect 18279 8820 18291 8823
rect 23566 8820 23572 8832
rect 18279 8792 23572 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 23566 8780 23572 8792
rect 23624 8780 23630 8832
rect 39850 8780 39856 8832
rect 39908 8820 39914 8832
rect 40405 8823 40463 8829
rect 40405 8820 40417 8823
rect 39908 8792 40417 8820
rect 39908 8780 39914 8792
rect 40405 8789 40417 8792
rect 40451 8789 40463 8823
rect 41782 8820 41788 8832
rect 41743 8792 41788 8820
rect 40405 8783 40463 8789
rect 41782 8780 41788 8792
rect 41840 8780 41846 8832
rect 42334 8820 42340 8832
rect 42295 8792 42340 8820
rect 42334 8780 42340 8792
rect 42392 8780 42398 8832
rect 42886 8820 42892 8832
rect 42847 8792 42892 8820
rect 42886 8780 42892 8792
rect 42944 8780 42950 8832
rect 43438 8820 43444 8832
rect 43399 8792 43444 8820
rect 43438 8780 43444 8792
rect 43496 8780 43502 8832
rect 43806 8780 43812 8832
rect 43864 8820 43870 8832
rect 43993 8823 44051 8829
rect 43993 8820 44005 8823
rect 43864 8792 44005 8820
rect 43864 8780 43870 8792
rect 43993 8789 44005 8792
rect 44039 8789 44051 8823
rect 44542 8820 44548 8832
rect 44503 8792 44548 8820
rect 43993 8783 44051 8789
rect 44542 8780 44548 8792
rect 44600 8780 44606 8832
rect 45646 8820 45652 8832
rect 45607 8792 45652 8820
rect 45646 8780 45652 8792
rect 45704 8780 45710 8832
rect 46106 8780 46112 8832
rect 46164 8820 46170 8832
rect 46201 8823 46259 8829
rect 46201 8820 46213 8823
rect 46164 8792 46213 8820
rect 46164 8780 46170 8792
rect 46201 8789 46213 8792
rect 46247 8789 46259 8823
rect 46201 8783 46259 8789
rect 46382 8780 46388 8832
rect 46440 8820 46446 8832
rect 46753 8823 46811 8829
rect 46753 8820 46765 8823
rect 46440 8792 46765 8820
rect 46440 8780 46446 8792
rect 46753 8789 46765 8792
rect 46799 8789 46811 8823
rect 46753 8783 46811 8789
rect 47026 8780 47032 8832
rect 47084 8820 47090 8832
rect 47305 8823 47363 8829
rect 47305 8820 47317 8823
rect 47084 8792 47317 8820
rect 47084 8780 47090 8792
rect 47305 8789 47317 8792
rect 47351 8789 47363 8823
rect 47305 8783 47363 8789
rect 47486 8780 47492 8832
rect 47544 8820 47550 8832
rect 47857 8823 47915 8829
rect 47857 8820 47869 8823
rect 47544 8792 47869 8820
rect 47544 8780 47550 8792
rect 47857 8789 47869 8792
rect 47903 8789 47915 8823
rect 48406 8820 48412 8832
rect 48367 8792 48412 8820
rect 47857 8783 47915 8789
rect 48406 8780 48412 8792
rect 48464 8780 48470 8832
rect 49050 8780 49056 8832
rect 49108 8820 49114 8832
rect 49605 8823 49663 8829
rect 49605 8820 49617 8823
rect 49108 8792 49617 8820
rect 49108 8780 49114 8792
rect 49605 8789 49617 8792
rect 49651 8820 49663 8823
rect 49694 8820 49700 8832
rect 49651 8792 49700 8820
rect 49651 8789 49663 8792
rect 49605 8783 49663 8789
rect 49694 8780 49700 8792
rect 49752 8780 49758 8832
rect 49970 8780 49976 8832
rect 50028 8820 50034 8832
rect 50157 8823 50215 8829
rect 50157 8820 50169 8823
rect 50028 8792 50169 8820
rect 50028 8780 50034 8792
rect 50157 8789 50169 8792
rect 50203 8820 50215 8823
rect 50430 8820 50436 8832
rect 50203 8792 50436 8820
rect 50203 8789 50215 8792
rect 50157 8783 50215 8789
rect 50430 8780 50436 8792
rect 50488 8780 50494 8832
rect 51442 8780 51448 8832
rect 51500 8820 51506 8832
rect 51537 8823 51595 8829
rect 51537 8820 51549 8823
rect 51500 8792 51549 8820
rect 51500 8780 51506 8792
rect 51537 8789 51549 8792
rect 51583 8820 51595 8823
rect 51626 8820 51632 8832
rect 51583 8792 51632 8820
rect 51583 8789 51595 8792
rect 51537 8783 51595 8789
rect 51626 8780 51632 8792
rect 51684 8780 51690 8832
rect 51994 8820 52000 8832
rect 51955 8792 52000 8820
rect 51994 8780 52000 8792
rect 52052 8780 52058 8832
rect 52454 8780 52460 8832
rect 52512 8820 52518 8832
rect 52549 8823 52607 8829
rect 52549 8820 52561 8823
rect 52512 8792 52561 8820
rect 52512 8780 52518 8792
rect 52549 8789 52561 8792
rect 52595 8789 52607 8823
rect 52549 8783 52607 8789
rect 53006 8780 53012 8832
rect 53064 8820 53070 8832
rect 53193 8823 53251 8829
rect 53193 8820 53205 8823
rect 53064 8792 53205 8820
rect 53064 8780 53070 8792
rect 53193 8789 53205 8792
rect 53239 8789 53251 8823
rect 54110 8820 54116 8832
rect 54071 8792 54116 8820
rect 53193 8783 53251 8789
rect 54110 8780 54116 8792
rect 54168 8780 54174 8832
rect 62850 8780 62856 8832
rect 62908 8820 62914 8832
rect 62945 8823 63003 8829
rect 62945 8820 62957 8823
rect 62908 8792 62957 8820
rect 62908 8780 62914 8792
rect 62945 8789 62957 8792
rect 62991 8820 63003 8823
rect 63126 8820 63132 8832
rect 62991 8792 63132 8820
rect 62991 8789 63003 8792
rect 62945 8783 63003 8789
rect 63126 8780 63132 8792
rect 63184 8780 63190 8832
rect 63494 8820 63500 8832
rect 63407 8792 63500 8820
rect 63494 8780 63500 8792
rect 63552 8820 63558 8832
rect 63770 8820 63776 8832
rect 63552 8792 63776 8820
rect 63552 8780 63558 8792
rect 63770 8780 63776 8792
rect 63828 8780 63834 8832
rect 63862 8780 63868 8832
rect 63920 8820 63926 8832
rect 64046 8820 64052 8832
rect 63920 8792 64052 8820
rect 63920 8780 63926 8792
rect 64046 8780 64052 8792
rect 64104 8780 64110 8832
rect 65058 8820 65064 8832
rect 65019 8792 65064 8820
rect 65058 8780 65064 8792
rect 65116 8780 65122 8832
rect 65426 8780 65432 8832
rect 65484 8820 65490 8832
rect 65705 8823 65763 8829
rect 65705 8820 65717 8823
rect 65484 8792 65717 8820
rect 65484 8780 65490 8792
rect 65705 8789 65717 8792
rect 65751 8789 65763 8823
rect 65705 8783 65763 8789
rect 67453 8823 67511 8829
rect 67453 8789 67465 8823
rect 67499 8820 67511 8823
rect 68094 8820 68100 8832
rect 67499 8792 68100 8820
rect 67499 8789 67511 8792
rect 67453 8783 67511 8789
rect 68094 8780 68100 8792
rect 68152 8780 68158 8832
rect 1104 8730 18952 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 14246 8730
rect 14298 8678 14310 8730
rect 14362 8678 14374 8730
rect 14426 8678 14438 8730
rect 14490 8678 18952 8730
rect 1104 8656 18952 8678
rect 37628 8730 68816 8752
rect 37628 8678 44246 8730
rect 44298 8678 44310 8730
rect 44362 8678 44374 8730
rect 44426 8678 44438 8730
rect 44490 8678 54246 8730
rect 54298 8678 54310 8730
rect 54362 8678 54374 8730
rect 54426 8678 54438 8730
rect 54490 8678 64246 8730
rect 64298 8678 64310 8730
rect 64362 8678 64374 8730
rect 64426 8678 64438 8730
rect 64490 8678 68816 8730
rect 37628 8656 68816 8678
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 4614 8616 4620 8628
rect 4479 8588 4620 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 6914 8616 6920 8628
rect 6875 8588 6920 8616
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 10778 8616 10784 8628
rect 9732 8588 10784 8616
rect 9732 8576 9738 8588
rect 10778 8576 10784 8588
rect 10836 8616 10842 8628
rect 15013 8619 15071 8625
rect 15013 8616 15025 8619
rect 10836 8588 15025 8616
rect 10836 8576 10842 8588
rect 15013 8585 15025 8588
rect 15059 8585 15071 8619
rect 15013 8579 15071 8585
rect 15381 8619 15439 8625
rect 15381 8585 15393 8619
rect 15427 8616 15439 8619
rect 17034 8616 17040 8628
rect 15427 8588 17040 8616
rect 15427 8585 15439 8588
rect 15381 8579 15439 8585
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 34425 8619 34483 8625
rect 34425 8585 34437 8619
rect 34471 8616 34483 8619
rect 34471 8588 40264 8616
rect 34471 8585 34483 8588
rect 34425 8579 34483 8585
rect 2682 8508 2688 8560
rect 2740 8548 2746 8560
rect 3145 8551 3203 8557
rect 3145 8548 3157 8551
rect 2740 8520 3157 8548
rect 2740 8508 2746 8520
rect 3145 8517 3157 8520
rect 3191 8517 3203 8551
rect 3145 8511 3203 8517
rect 14902 8551 14960 8557
rect 14902 8517 14914 8551
rect 14948 8548 14960 8551
rect 16298 8548 16304 8560
rect 14948 8520 16304 8548
rect 14948 8517 14960 8520
rect 14902 8511 14960 8517
rect 16298 8508 16304 8520
rect 16356 8508 16362 8560
rect 33597 8551 33655 8557
rect 33597 8517 33609 8551
rect 33643 8548 33655 8551
rect 33643 8520 40172 8548
rect 33643 8517 33655 8520
rect 33597 8511 33655 8517
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 14458 8480 14464 8492
rect 12575 8452 14464 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 15102 8480 15108 8492
rect 15063 8452 15108 8480
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 24486 8480 24492 8492
rect 15344 8452 24492 8480
rect 15344 8440 15350 8452
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 2590 8372 2596 8424
rect 2648 8412 2654 8424
rect 2685 8415 2743 8421
rect 2685 8412 2697 8415
rect 2648 8384 2697 8412
rect 2648 8372 2654 8384
rect 2685 8381 2697 8384
rect 2731 8381 2743 8415
rect 2685 8375 2743 8381
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 13044 8384 13185 8412
rect 13044 8372 13050 8384
rect 13173 8381 13185 8384
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8412 14795 8415
rect 15010 8412 15016 8424
rect 14783 8384 15016 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 1949 8347 2007 8353
rect 1949 8313 1961 8347
rect 1995 8344 2007 8347
rect 3050 8344 3056 8356
rect 1995 8316 3056 8344
rect 1995 8313 2007 8316
rect 1949 8307 2007 8313
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 3326 8304 3332 8356
rect 3384 8344 3390 8356
rect 3697 8347 3755 8353
rect 3697 8344 3709 8347
rect 3384 8316 3709 8344
rect 3384 8304 3390 8316
rect 3697 8313 3709 8316
rect 3743 8313 3755 8347
rect 3697 8307 3755 8313
rect 5537 8347 5595 8353
rect 5537 8313 5549 8347
rect 5583 8344 5595 8347
rect 5718 8344 5724 8356
rect 5583 8316 5724 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 5718 8304 5724 8316
rect 5776 8344 5782 8356
rect 6178 8344 6184 8356
rect 5776 8316 6184 8344
rect 5776 8304 5782 8316
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 7558 8344 7564 8356
rect 7515 8316 7564 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 8110 8344 8116 8356
rect 8071 8316 8116 8344
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 9030 8304 9036 8356
rect 9088 8344 9094 8356
rect 9309 8347 9367 8353
rect 9309 8344 9321 8347
rect 9088 8316 9321 8344
rect 9088 8304 9094 8316
rect 9309 8313 9321 8316
rect 9355 8313 9367 8347
rect 9309 8307 9367 8313
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 9953 8347 10011 8353
rect 9953 8344 9965 8347
rect 9916 8316 9965 8344
rect 9916 8304 9922 8316
rect 9953 8313 9965 8316
rect 9999 8313 10011 8347
rect 10778 8344 10784 8356
rect 10739 8316 10784 8344
rect 9953 8307 10011 8313
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 14292 8344 14320 8375
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 16408 8421 16436 8452
rect 24486 8440 24492 8452
rect 24544 8440 24550 8492
rect 31938 8440 31944 8492
rect 31996 8480 32002 8492
rect 31996 8452 39436 8480
rect 31996 8440 32002 8452
rect 39408 8424 39436 8452
rect 16393 8415 16451 8421
rect 16393 8381 16405 8415
rect 16439 8381 16451 8415
rect 16393 8375 16451 8381
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 14826 8344 14832 8356
rect 14292 8316 14832 8344
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 17512 8344 17540 8375
rect 18046 8372 18052 8424
rect 18104 8412 18110 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 18104 8384 18153 8412
rect 18104 8372 18110 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 37090 8372 37096 8424
rect 37148 8412 37154 8424
rect 38105 8415 38163 8421
rect 38105 8412 38117 8415
rect 37148 8384 38117 8412
rect 37148 8372 37154 8384
rect 38105 8381 38117 8384
rect 38151 8412 38163 8415
rect 38470 8412 38476 8424
rect 38151 8384 38476 8412
rect 38151 8381 38163 8384
rect 38105 8375 38163 8381
rect 38470 8372 38476 8384
rect 38528 8372 38534 8424
rect 38749 8415 38807 8421
rect 38749 8381 38761 8415
rect 38795 8381 38807 8415
rect 39390 8412 39396 8424
rect 39351 8384 39396 8412
rect 38749 8375 38807 8381
rect 17678 8344 17684 8356
rect 17512 8316 17684 8344
rect 17678 8304 17684 8316
rect 17736 8344 17742 8356
rect 21082 8344 21088 8356
rect 17736 8316 21088 8344
rect 17736 8304 17742 8316
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 32950 8304 32956 8356
rect 33008 8344 33014 8356
rect 38654 8344 38660 8356
rect 33008 8316 38660 8344
rect 33008 8304 33014 8316
rect 38654 8304 38660 8316
rect 38712 8344 38718 8356
rect 38764 8344 38792 8375
rect 39390 8372 39396 8384
rect 39448 8372 39454 8424
rect 40034 8412 40040 8424
rect 39995 8384 40040 8412
rect 40034 8372 40040 8384
rect 40092 8372 40098 8424
rect 40144 8412 40172 8520
rect 40236 8480 40264 8588
rect 41046 8576 41052 8628
rect 41104 8616 41110 8628
rect 48406 8616 48412 8628
rect 41104 8588 48412 8616
rect 41104 8576 41110 8588
rect 48406 8576 48412 8588
rect 48464 8576 48470 8628
rect 50341 8619 50399 8625
rect 50341 8585 50353 8619
rect 50387 8616 50399 8619
rect 50614 8616 50620 8628
rect 50387 8588 50620 8616
rect 50387 8585 50399 8588
rect 50341 8579 50399 8585
rect 50614 8576 50620 8588
rect 50672 8576 50678 8628
rect 50706 8576 50712 8628
rect 50764 8616 50770 8628
rect 50801 8619 50859 8625
rect 50801 8616 50813 8619
rect 50764 8588 50813 8616
rect 50764 8576 50770 8588
rect 50801 8585 50813 8588
rect 50847 8616 50859 8619
rect 51442 8616 51448 8628
rect 50847 8588 51448 8616
rect 50847 8585 50859 8588
rect 50801 8579 50859 8585
rect 51442 8576 51448 8588
rect 51500 8576 51506 8628
rect 51537 8619 51595 8625
rect 51537 8585 51549 8619
rect 51583 8616 51595 8619
rect 51810 8616 51816 8628
rect 51583 8588 51816 8616
rect 51583 8585 51595 8588
rect 51537 8579 51595 8585
rect 51810 8576 51816 8588
rect 51868 8576 51874 8628
rect 51902 8576 51908 8628
rect 51960 8616 51966 8628
rect 51997 8619 52055 8625
rect 51997 8616 52009 8619
rect 51960 8588 52009 8616
rect 51960 8576 51966 8588
rect 51997 8585 52009 8588
rect 52043 8585 52055 8619
rect 51997 8579 52055 8585
rect 54018 8576 54024 8628
rect 54076 8616 54082 8628
rect 54113 8619 54171 8625
rect 54113 8616 54125 8619
rect 54076 8588 54125 8616
rect 54076 8576 54082 8588
rect 54113 8585 54125 8588
rect 54159 8616 54171 8619
rect 55030 8616 55036 8628
rect 54159 8588 55036 8616
rect 54159 8585 54171 8588
rect 54113 8579 54171 8585
rect 55030 8576 55036 8588
rect 55088 8576 55094 8628
rect 61378 8616 61384 8628
rect 61339 8588 61384 8616
rect 61378 8576 61384 8588
rect 61436 8576 61442 8628
rect 40494 8508 40500 8560
rect 40552 8548 40558 8560
rect 43530 8548 43536 8560
rect 40552 8520 43536 8548
rect 40552 8508 40558 8520
rect 43530 8508 43536 8520
rect 43588 8508 43594 8560
rect 43714 8508 43720 8560
rect 43772 8548 43778 8560
rect 43990 8548 43996 8560
rect 43772 8520 43996 8548
rect 43772 8508 43778 8520
rect 43990 8508 43996 8520
rect 44048 8508 44054 8560
rect 40236 8452 40632 8480
rect 40310 8412 40316 8424
rect 40144 8384 40316 8412
rect 40310 8372 40316 8384
rect 40368 8412 40374 8424
rect 40497 8415 40555 8421
rect 40497 8412 40509 8415
rect 40368 8384 40509 8412
rect 40368 8372 40374 8384
rect 40497 8381 40509 8384
rect 40543 8381 40555 8415
rect 40604 8412 40632 8452
rect 41414 8412 41420 8424
rect 40604 8384 41420 8412
rect 40497 8375 40555 8381
rect 41414 8372 41420 8384
rect 41472 8412 41478 8424
rect 42245 8415 42303 8421
rect 41472 8384 41517 8412
rect 41472 8372 41478 8384
rect 42245 8381 42257 8415
rect 42291 8412 42303 8415
rect 42610 8412 42616 8424
rect 42291 8384 42616 8412
rect 42291 8381 42303 8384
rect 42245 8375 42303 8381
rect 38712 8316 38792 8344
rect 38712 8304 38718 8316
rect 41322 8304 41328 8356
rect 41380 8344 41386 8356
rect 42260 8344 42288 8375
rect 42610 8372 42616 8384
rect 42668 8372 42674 8424
rect 43530 8412 43536 8424
rect 43491 8384 43536 8412
rect 43530 8372 43536 8384
rect 43588 8372 43594 8424
rect 44637 8415 44695 8421
rect 44637 8381 44649 8415
rect 44683 8412 44695 8415
rect 45094 8412 45100 8424
rect 44683 8384 45100 8412
rect 44683 8381 44695 8384
rect 44637 8375 44695 8381
rect 45094 8372 45100 8384
rect 45152 8372 45158 8424
rect 66257 8415 66315 8421
rect 66257 8381 66269 8415
rect 66303 8412 66315 8415
rect 67082 8412 67088 8424
rect 66303 8384 67088 8412
rect 66303 8381 66315 8384
rect 66257 8375 66315 8381
rect 67082 8372 67088 8384
rect 67140 8372 67146 8424
rect 67450 8412 67456 8424
rect 67363 8384 67456 8412
rect 67450 8372 67456 8384
rect 67508 8372 67514 8424
rect 68094 8412 68100 8424
rect 68055 8384 68100 8412
rect 68094 8372 68100 8384
rect 68152 8372 68158 8424
rect 45738 8344 45744 8356
rect 41380 8316 42288 8344
rect 45699 8316 45744 8344
rect 41380 8304 41386 8316
rect 45738 8304 45744 8316
rect 45796 8304 45802 8356
rect 46658 8304 46664 8356
rect 46716 8344 46722 8356
rect 46753 8347 46811 8353
rect 46753 8344 46765 8347
rect 46716 8316 46765 8344
rect 46716 8304 46722 8316
rect 46753 8313 46765 8316
rect 46799 8313 46811 8347
rect 46753 8307 46811 8313
rect 47118 8304 47124 8356
rect 47176 8344 47182 8356
rect 47305 8347 47363 8353
rect 47305 8344 47317 8347
rect 47176 8316 47317 8344
rect 47176 8304 47182 8316
rect 47305 8313 47317 8316
rect 47351 8313 47363 8347
rect 47305 8307 47363 8313
rect 48130 8304 48136 8356
rect 48188 8344 48194 8356
rect 48317 8347 48375 8353
rect 48317 8344 48329 8347
rect 48188 8316 48329 8344
rect 48188 8304 48194 8316
rect 48317 8313 48329 8316
rect 48363 8313 48375 8347
rect 48317 8307 48375 8313
rect 48498 8304 48504 8356
rect 48556 8344 48562 8356
rect 48777 8347 48835 8353
rect 48777 8344 48789 8347
rect 48556 8316 48789 8344
rect 48556 8304 48562 8316
rect 48777 8313 48789 8316
rect 48823 8313 48835 8347
rect 48777 8307 48835 8313
rect 49050 8304 49056 8356
rect 49108 8344 49114 8356
rect 49329 8347 49387 8353
rect 49329 8344 49341 8347
rect 49108 8316 49341 8344
rect 49108 8304 49114 8316
rect 49329 8313 49341 8316
rect 49375 8313 49387 8347
rect 49329 8307 49387 8313
rect 52270 8304 52276 8356
rect 52328 8344 52334 8356
rect 52549 8347 52607 8353
rect 52549 8344 52561 8347
rect 52328 8316 52561 8344
rect 52328 8304 52334 8316
rect 52549 8313 52561 8316
rect 52595 8313 52607 8347
rect 52549 8307 52607 8313
rect 53374 8304 53380 8356
rect 53432 8344 53438 8356
rect 53469 8347 53527 8353
rect 53469 8344 53481 8347
rect 53432 8316 53481 8344
rect 53432 8304 53438 8316
rect 53469 8313 53481 8316
rect 53515 8313 53527 8347
rect 54662 8344 54668 8356
rect 54623 8316 54668 8344
rect 53469 8307 53527 8313
rect 54662 8304 54668 8316
rect 54720 8304 54726 8356
rect 55214 8344 55220 8356
rect 55175 8316 55220 8344
rect 55214 8304 55220 8316
rect 55272 8304 55278 8356
rect 55674 8344 55680 8356
rect 55635 8316 55680 8344
rect 55674 8304 55680 8316
rect 55732 8304 55738 8356
rect 62206 8344 62212 8356
rect 62167 8316 62212 8344
rect 62206 8304 62212 8316
rect 62264 8304 62270 8356
rect 62574 8304 62580 8356
rect 62632 8344 62638 8356
rect 62945 8347 63003 8353
rect 62945 8344 62957 8347
rect 62632 8316 62957 8344
rect 62632 8304 62638 8316
rect 62945 8313 62957 8316
rect 62991 8313 63003 8347
rect 62945 8307 63003 8313
rect 64509 8347 64567 8353
rect 64509 8313 64521 8347
rect 64555 8344 64567 8347
rect 64598 8344 64604 8356
rect 64555 8316 64604 8344
rect 64555 8313 64567 8316
rect 64509 8307 64567 8313
rect 64598 8304 64604 8316
rect 64656 8304 64662 8356
rect 65610 8344 65616 8356
rect 65571 8316 65616 8344
rect 65610 8304 65616 8316
rect 65668 8304 65674 8356
rect 66438 8304 66444 8356
rect 66496 8344 66502 8356
rect 66717 8347 66775 8353
rect 66717 8344 66729 8347
rect 66496 8316 66729 8344
rect 66496 8304 66502 8316
rect 66717 8313 66729 8316
rect 66763 8313 66775 8347
rect 67468 8344 67496 8372
rect 68186 8344 68192 8356
rect 67468 8316 68192 8344
rect 66717 8307 66775 8313
rect 68186 8304 68192 8316
rect 68244 8304 68250 8356
rect 2866 8236 2872 8288
rect 2924 8276 2930 8288
rect 4890 8276 4896 8288
rect 2924 8248 4896 8276
rect 2924 8236 2930 8248
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 8754 8276 8760 8288
rect 8715 8248 8760 8276
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 11977 8279 12035 8285
rect 11977 8245 11989 8279
rect 12023 8276 12035 8279
rect 12250 8276 12256 8288
rect 12023 8248 12256 8276
rect 12023 8245 12035 8248
rect 11977 8239 12035 8245
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 15378 8276 15384 8288
rect 15252 8248 15384 8276
rect 15252 8236 15258 8248
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 41414 8236 41420 8288
rect 41472 8276 41478 8288
rect 41690 8276 41696 8288
rect 41472 8248 41696 8276
rect 41472 8236 41478 8248
rect 41690 8236 41696 8248
rect 41748 8236 41754 8288
rect 43990 8276 43996 8288
rect 43951 8248 43996 8276
rect 43990 8236 43996 8248
rect 44048 8236 44054 8288
rect 45189 8279 45247 8285
rect 45189 8245 45201 8279
rect 45235 8276 45247 8279
rect 45370 8276 45376 8288
rect 45235 8248 45376 8276
rect 45235 8245 45247 8248
rect 45189 8239 45247 8245
rect 45370 8236 45376 8248
rect 45428 8236 45434 8288
rect 46198 8276 46204 8288
rect 46159 8248 46204 8276
rect 46198 8236 46204 8248
rect 46256 8236 46262 8288
rect 57330 8236 57336 8288
rect 57388 8276 57394 8288
rect 57514 8276 57520 8288
rect 57388 8248 57520 8276
rect 57388 8236 57394 8248
rect 57514 8236 57520 8248
rect 57572 8236 57578 8288
rect 64690 8236 64696 8288
rect 64748 8276 64754 8288
rect 64969 8279 65027 8285
rect 64969 8276 64981 8279
rect 64748 8248 64981 8276
rect 64748 8236 64754 8248
rect 64969 8245 64981 8248
rect 65015 8245 65027 8279
rect 64969 8239 65027 8245
rect 1104 8186 18952 8208
rect 1104 8134 9246 8186
rect 9298 8134 9310 8186
rect 9362 8134 9374 8186
rect 9426 8134 9438 8186
rect 9490 8134 18952 8186
rect 1104 8112 18952 8134
rect 37628 8186 68816 8208
rect 37628 8134 39246 8186
rect 39298 8134 39310 8186
rect 39362 8134 39374 8186
rect 39426 8134 39438 8186
rect 39490 8134 49246 8186
rect 49298 8134 49310 8186
rect 49362 8134 49374 8186
rect 49426 8134 49438 8186
rect 49490 8134 59246 8186
rect 59298 8134 59310 8186
rect 59362 8134 59374 8186
rect 59426 8134 59438 8186
rect 59490 8134 68816 8186
rect 37628 8112 68816 8134
rect 6270 8072 6276 8084
rect 6231 8044 6276 8072
rect 6270 8032 6276 8044
rect 6328 8032 6334 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 15010 8072 15016 8084
rect 14608 8044 15016 8072
rect 14608 8032 14614 8044
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 17034 8072 17040 8084
rect 15396 8044 17040 8072
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7936 11115 7939
rect 11238 7936 11244 7948
rect 11103 7908 11244 7936
rect 11103 7905 11115 7908
rect 11057 7899 11115 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11756 7908 11897 7936
rect 11756 7896 11762 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7905 12587 7939
rect 12529 7899 12587 7905
rect 12544 7868 12572 7899
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12676 7908 13001 7936
rect 12676 7896 12682 7908
rect 12989 7905 13001 7908
rect 13035 7905 13047 7939
rect 12989 7899 13047 7905
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 13906 7936 13912 7948
rect 13863 7908 13912 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 15396 7945 15424 8044
rect 17034 8032 17040 8044
rect 17092 8072 17098 8084
rect 17218 8072 17224 8084
rect 17092 8044 17224 8072
rect 17092 8032 17098 8044
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 36906 8032 36912 8084
rect 36964 8072 36970 8084
rect 36964 8044 40264 8072
rect 36964 8032 36970 8044
rect 16482 8004 16488 8016
rect 16040 7976 16488 8004
rect 16040 7945 16068 7976
rect 16482 7964 16488 7976
rect 16540 8004 16546 8016
rect 23290 8004 23296 8016
rect 16540 7976 23296 8004
rect 16540 7964 16546 7976
rect 23290 7964 23296 7976
rect 23348 7964 23354 8016
rect 34974 7964 34980 8016
rect 35032 8004 35038 8016
rect 38654 8004 38660 8016
rect 35032 7976 38660 8004
rect 35032 7964 35038 7976
rect 38654 7964 38660 7976
rect 38712 8004 38718 8016
rect 38712 7976 38792 8004
rect 38712 7964 38718 7976
rect 15381 7939 15439 7945
rect 15381 7905 15393 7939
rect 15427 7905 15439 7939
rect 15381 7899 15439 7905
rect 16025 7939 16083 7945
rect 16025 7905 16037 7939
rect 16071 7905 16083 7939
rect 16025 7899 16083 7905
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 17126 7936 17132 7948
rect 17087 7908 17132 7936
rect 16669 7899 16727 7905
rect 12710 7868 12716 7880
rect 12544 7840 12716 7868
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 16684 7868 16712 7899
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 18230 7936 18236 7948
rect 18191 7908 18236 7936
rect 18230 7896 18236 7908
rect 18288 7936 18294 7948
rect 23750 7936 23756 7948
rect 18288 7908 23756 7936
rect 18288 7896 18294 7908
rect 23750 7896 23756 7908
rect 23808 7896 23814 7948
rect 32030 7896 32036 7948
rect 32088 7936 32094 7948
rect 37918 7936 37924 7948
rect 32088 7908 37924 7936
rect 32088 7896 32094 7908
rect 37918 7896 37924 7908
rect 37976 7936 37982 7948
rect 38764 7945 38792 7976
rect 39022 7964 39028 8016
rect 39080 8004 39086 8016
rect 40236 8004 40264 8044
rect 40310 8032 40316 8084
rect 40368 8072 40374 8084
rect 42978 8072 42984 8084
rect 40368 8044 42984 8072
rect 40368 8032 40374 8044
rect 42978 8032 42984 8044
rect 43036 8032 43042 8084
rect 55309 8075 55367 8081
rect 55309 8041 55321 8075
rect 55355 8072 55367 8075
rect 55398 8072 55404 8084
rect 55355 8044 55404 8072
rect 55355 8041 55367 8044
rect 55309 8035 55367 8041
rect 55398 8032 55404 8044
rect 55456 8032 55462 8084
rect 56042 8032 56048 8084
rect 56100 8072 56106 8084
rect 56689 8075 56747 8081
rect 56689 8072 56701 8075
rect 56100 8044 56701 8072
rect 56100 8032 56106 8044
rect 56689 8041 56701 8044
rect 56735 8041 56747 8075
rect 56689 8035 56747 8041
rect 57238 8032 57244 8084
rect 57296 8072 57302 8084
rect 57333 8075 57391 8081
rect 57333 8072 57345 8075
rect 57296 8044 57345 8072
rect 57296 8032 57302 8044
rect 57333 8041 57345 8044
rect 57379 8041 57391 8075
rect 57333 8035 57391 8041
rect 57422 8032 57428 8084
rect 57480 8072 57486 8084
rect 57977 8075 58035 8081
rect 57977 8072 57989 8075
rect 57480 8044 57989 8072
rect 57480 8032 57486 8044
rect 57977 8041 57989 8044
rect 58023 8041 58035 8075
rect 57977 8035 58035 8041
rect 46198 8004 46204 8016
rect 39080 7976 39804 8004
rect 40236 7976 46204 8004
rect 39080 7964 39086 7976
rect 38105 7939 38163 7945
rect 38105 7936 38117 7939
rect 37976 7908 38117 7936
rect 37976 7896 37982 7908
rect 38105 7905 38117 7908
rect 38151 7905 38163 7939
rect 38105 7899 38163 7905
rect 38749 7939 38807 7945
rect 38749 7905 38761 7939
rect 38795 7905 38807 7939
rect 38749 7899 38807 7905
rect 39393 7939 39451 7945
rect 39393 7905 39405 7939
rect 39439 7936 39451 7939
rect 39666 7936 39672 7948
rect 39439 7908 39672 7936
rect 39439 7905 39451 7908
rect 39393 7899 39451 7905
rect 16942 7868 16948 7880
rect 16684 7840 16948 7868
rect 16942 7828 16948 7840
rect 17000 7868 17006 7880
rect 20990 7868 20996 7880
rect 17000 7840 20996 7868
rect 17000 7828 17006 7840
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 37461 7871 37519 7877
rect 37461 7837 37473 7871
rect 37507 7868 37519 7871
rect 39408 7868 39436 7899
rect 39666 7896 39672 7908
rect 39724 7896 39730 7948
rect 37507 7840 39436 7868
rect 39776 7868 39804 7976
rect 40957 7939 41015 7945
rect 40957 7905 40969 7939
rect 41003 7936 41015 7939
rect 41414 7936 41420 7948
rect 41003 7908 41420 7936
rect 41003 7905 41015 7908
rect 40957 7899 41015 7905
rect 41414 7896 41420 7908
rect 41472 7896 41478 7948
rect 41601 7939 41659 7945
rect 41601 7905 41613 7939
rect 41647 7936 41659 7939
rect 41874 7936 41880 7948
rect 41647 7908 41880 7936
rect 41647 7905 41659 7908
rect 41601 7899 41659 7905
rect 41874 7896 41880 7908
rect 41932 7896 41938 7948
rect 42245 7939 42303 7945
rect 42245 7905 42257 7939
rect 42291 7936 42303 7939
rect 42794 7936 42800 7948
rect 42291 7908 42800 7936
rect 42291 7905 42303 7908
rect 42245 7899 42303 7905
rect 42260 7868 42288 7899
rect 42794 7896 42800 7908
rect 42852 7896 42858 7948
rect 42889 7939 42947 7945
rect 42889 7905 42901 7939
rect 42935 7936 42947 7939
rect 42978 7936 42984 7948
rect 42935 7908 42984 7936
rect 42935 7905 42947 7908
rect 42889 7899 42947 7905
rect 42978 7896 42984 7908
rect 43036 7896 43042 7948
rect 43548 7945 43576 7976
rect 46198 7964 46204 7976
rect 46256 7964 46262 8016
rect 43533 7939 43591 7945
rect 43533 7905 43545 7939
rect 43579 7905 43591 7939
rect 43533 7899 43591 7905
rect 43898 7896 43904 7948
rect 43956 7936 43962 7948
rect 43993 7939 44051 7945
rect 43993 7936 44005 7939
rect 43956 7908 44005 7936
rect 43956 7896 43962 7908
rect 43993 7905 44005 7908
rect 44039 7936 44051 7939
rect 44082 7936 44088 7948
rect 44039 7908 44088 7936
rect 44039 7905 44051 7908
rect 43993 7899 44051 7905
rect 44082 7896 44088 7908
rect 44140 7896 44146 7948
rect 44637 7939 44695 7945
rect 44637 7905 44649 7939
rect 44683 7936 44695 7939
rect 44910 7936 44916 7948
rect 44683 7908 44916 7936
rect 44683 7905 44695 7908
rect 44637 7899 44695 7905
rect 44910 7896 44916 7908
rect 44968 7896 44974 7948
rect 46934 7896 46940 7948
rect 46992 7936 46998 7948
rect 55950 7936 55956 7948
rect 46992 7908 55956 7936
rect 46992 7896 46998 7908
rect 55950 7896 55956 7908
rect 56008 7896 56014 7948
rect 67174 7896 67180 7948
rect 67232 7936 67238 7948
rect 67361 7939 67419 7945
rect 67361 7936 67373 7939
rect 67232 7908 67373 7936
rect 67232 7896 67238 7908
rect 67361 7905 67373 7908
rect 67407 7905 67419 7939
rect 67361 7899 67419 7905
rect 67634 7896 67640 7948
rect 67692 7936 67698 7948
rect 68002 7936 68008 7948
rect 67692 7908 68008 7936
rect 67692 7896 67698 7908
rect 68002 7896 68008 7908
rect 68060 7896 68066 7948
rect 39776 7840 42288 7868
rect 37507 7837 37519 7840
rect 37461 7831 37519 7837
rect 43622 7828 43628 7880
rect 43680 7868 43686 7880
rect 45554 7868 45560 7880
rect 43680 7840 45560 7868
rect 43680 7828 43686 7840
rect 45554 7828 45560 7840
rect 45612 7828 45618 7880
rect 48406 7828 48412 7880
rect 48464 7868 48470 7880
rect 48961 7871 49019 7877
rect 48961 7868 48973 7871
rect 48464 7840 48973 7868
rect 48464 7828 48470 7840
rect 48961 7837 48973 7840
rect 49007 7837 49019 7871
rect 48961 7831 49019 7837
rect 66622 7828 66628 7880
rect 66680 7868 66686 7880
rect 68278 7868 68284 7880
rect 66680 7840 68284 7868
rect 66680 7828 66686 7840
rect 68278 7828 68284 7840
rect 68336 7828 68342 7880
rect 2777 7803 2835 7809
rect 2777 7769 2789 7803
rect 2823 7800 2835 7803
rect 15194 7800 15200 7812
rect 2823 7772 15200 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 15194 7760 15200 7772
rect 15252 7760 15258 7812
rect 15286 7760 15292 7812
rect 15344 7800 15350 7812
rect 23658 7800 23664 7812
rect 15344 7772 23664 7800
rect 15344 7760 15350 7772
rect 23658 7760 23664 7772
rect 23716 7760 23722 7812
rect 38654 7760 38660 7812
rect 38712 7800 38718 7812
rect 41874 7800 41880 7812
rect 38712 7772 41880 7800
rect 38712 7760 38718 7772
rect 41874 7760 41880 7772
rect 41932 7760 41938 7812
rect 48590 7760 48596 7812
rect 48648 7800 48654 7812
rect 49513 7803 49571 7809
rect 49513 7800 49525 7803
rect 48648 7772 49525 7800
rect 48648 7760 48654 7772
rect 49513 7769 49525 7772
rect 49559 7769 49571 7803
rect 49513 7763 49571 7769
rect 63681 7803 63739 7809
rect 63681 7769 63693 7803
rect 63727 7800 63739 7803
rect 65334 7800 65340 7812
rect 63727 7772 65340 7800
rect 63727 7769 63739 7772
rect 63681 7763 63739 7769
rect 65334 7760 65340 7772
rect 65392 7760 65398 7812
rect 65429 7803 65487 7809
rect 65429 7769 65441 7803
rect 65475 7800 65487 7803
rect 66162 7800 66168 7812
rect 65475 7772 66168 7800
rect 65475 7769 65487 7772
rect 65429 7763 65487 7769
rect 66162 7760 66168 7772
rect 66220 7760 66226 7812
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3878 7732 3884 7744
rect 3839 7704 3884 7732
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4525 7735 4583 7741
rect 4525 7701 4537 7735
rect 4571 7732 4583 7735
rect 4798 7732 4804 7744
rect 4571 7704 4804 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 4948 7704 5181 7732
rect 4948 7692 4954 7704
rect 5169 7701 5181 7704
rect 5215 7701 5227 7735
rect 5169 7695 5227 7701
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5721 7735 5779 7741
rect 5721 7732 5733 7735
rect 5592 7704 5733 7732
rect 5592 7692 5598 7704
rect 5721 7701 5733 7704
rect 5767 7701 5779 7735
rect 5721 7695 5779 7701
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7374 7732 7380 7744
rect 6963 7704 7380 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 7561 7735 7619 7741
rect 7561 7701 7573 7735
rect 7607 7732 7619 7735
rect 7926 7732 7932 7744
rect 7607 7704 7932 7732
rect 7607 7701 7619 7704
rect 7561 7695 7619 7701
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8386 7732 8392 7744
rect 8343 7704 8392 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 8996 7704 9137 7732
rect 8996 7692 9002 7704
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 9674 7732 9680 7744
rect 9635 7704 9680 7732
rect 9125 7695 9183 7701
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10413 7735 10471 7741
rect 10413 7701 10425 7735
rect 10459 7732 10471 7735
rect 11514 7732 11520 7744
rect 10459 7704 11520 7732
rect 10459 7701 10471 7704
rect 10413 7695 10471 7701
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 14737 7735 14795 7741
rect 14737 7701 14749 7735
rect 14783 7732 14795 7735
rect 16482 7732 16488 7744
rect 14783 7704 16488 7732
rect 14783 7701 14795 7704
rect 14737 7695 14795 7701
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 39666 7692 39672 7744
rect 39724 7732 39730 7744
rect 44726 7732 44732 7744
rect 39724 7704 44732 7732
rect 39724 7692 39730 7704
rect 44726 7692 44732 7704
rect 44784 7692 44790 7744
rect 45554 7692 45560 7744
rect 45612 7732 45618 7744
rect 45649 7735 45707 7741
rect 45649 7732 45661 7735
rect 45612 7704 45661 7732
rect 45612 7692 45618 7704
rect 45649 7701 45661 7704
rect 45695 7701 45707 7735
rect 46198 7732 46204 7744
rect 46159 7704 46204 7732
rect 45649 7695 45707 7701
rect 46198 7692 46204 7704
rect 46256 7692 46262 7744
rect 46842 7732 46848 7744
rect 46803 7704 46848 7732
rect 46842 7692 46848 7704
rect 46900 7692 46906 7744
rect 47210 7692 47216 7744
rect 47268 7732 47274 7744
rect 47305 7735 47363 7741
rect 47305 7732 47317 7735
rect 47268 7704 47317 7732
rect 47268 7692 47274 7704
rect 47305 7701 47317 7704
rect 47351 7701 47363 7735
rect 47854 7732 47860 7744
rect 47815 7704 47860 7732
rect 47305 7695 47363 7701
rect 47854 7692 47860 7704
rect 47912 7692 47918 7744
rect 48314 7692 48320 7744
rect 48372 7732 48378 7744
rect 48409 7735 48467 7741
rect 48409 7732 48421 7735
rect 48372 7704 48421 7732
rect 48372 7692 48378 7704
rect 48409 7701 48421 7704
rect 48455 7701 48467 7735
rect 48409 7695 48467 7701
rect 50157 7735 50215 7741
rect 50157 7701 50169 7735
rect 50203 7732 50215 7735
rect 50338 7732 50344 7744
rect 50203 7704 50344 7732
rect 50203 7701 50215 7704
rect 50157 7695 50215 7701
rect 50338 7692 50344 7704
rect 50396 7692 50402 7744
rect 50890 7732 50896 7744
rect 50851 7704 50896 7732
rect 50890 7692 50896 7704
rect 50948 7692 50954 7744
rect 51442 7732 51448 7744
rect 51403 7704 51448 7732
rect 51442 7692 51448 7704
rect 51500 7692 51506 7744
rect 52086 7732 52092 7744
rect 52047 7704 52092 7732
rect 52086 7692 52092 7704
rect 52144 7692 52150 7744
rect 52362 7692 52368 7744
rect 52420 7732 52426 7744
rect 52549 7735 52607 7741
rect 52549 7732 52561 7735
rect 52420 7704 52561 7732
rect 52420 7692 52426 7704
rect 52549 7701 52561 7704
rect 52595 7701 52607 7735
rect 52549 7695 52607 7701
rect 52822 7692 52828 7744
rect 52880 7732 52886 7744
rect 53101 7735 53159 7741
rect 53101 7732 53113 7735
rect 52880 7704 53113 7732
rect 52880 7692 52886 7704
rect 53101 7701 53113 7704
rect 53147 7701 53159 7735
rect 53101 7695 53159 7701
rect 53466 7692 53472 7744
rect 53524 7732 53530 7744
rect 53653 7735 53711 7741
rect 53653 7732 53665 7735
rect 53524 7704 53665 7732
rect 53524 7692 53530 7704
rect 53653 7701 53665 7704
rect 53699 7732 53711 7735
rect 53742 7732 53748 7744
rect 53699 7704 53748 7732
rect 53699 7701 53711 7704
rect 53653 7695 53711 7701
rect 53742 7692 53748 7704
rect 53800 7692 53806 7744
rect 54573 7735 54631 7741
rect 54573 7701 54585 7735
rect 54619 7732 54631 7735
rect 54846 7732 54852 7744
rect 54619 7704 54852 7732
rect 54619 7701 54631 7704
rect 54573 7695 54631 7701
rect 54846 7692 54852 7704
rect 54904 7692 54910 7744
rect 55950 7692 55956 7744
rect 56008 7732 56014 7744
rect 56137 7735 56195 7741
rect 56137 7732 56149 7735
rect 56008 7704 56149 7732
rect 56008 7692 56014 7704
rect 56137 7701 56149 7704
rect 56183 7701 56195 7735
rect 60826 7732 60832 7744
rect 60787 7704 60832 7732
rect 56137 7695 56195 7701
rect 60826 7692 60832 7704
rect 60884 7692 60890 7744
rect 61930 7732 61936 7744
rect 61891 7704 61936 7732
rect 61930 7692 61936 7704
rect 61988 7692 61994 7744
rect 62482 7732 62488 7744
rect 62443 7704 62488 7732
rect 62482 7692 62488 7704
rect 62540 7692 62546 7744
rect 63034 7732 63040 7744
rect 62995 7704 63040 7732
rect 63034 7692 63040 7704
rect 63092 7692 63098 7744
rect 63862 7692 63868 7744
rect 63920 7732 63926 7744
rect 64141 7735 64199 7741
rect 64141 7732 64153 7735
rect 63920 7704 64153 7732
rect 63920 7692 63926 7704
rect 64141 7701 64153 7704
rect 64187 7701 64199 7735
rect 64141 7695 64199 7701
rect 64877 7735 64935 7741
rect 64877 7701 64889 7735
rect 64923 7732 64935 7735
rect 65150 7732 65156 7744
rect 64923 7704 65156 7732
rect 64923 7701 64935 7704
rect 64877 7695 64935 7701
rect 65150 7692 65156 7704
rect 65208 7692 65214 7744
rect 65886 7732 65892 7744
rect 65847 7704 65892 7732
rect 65886 7692 65892 7704
rect 65944 7692 65950 7744
rect 66622 7732 66628 7744
rect 66583 7704 66628 7732
rect 66622 7692 66628 7704
rect 66680 7692 66686 7744
rect 1104 7642 18952 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 14246 7642
rect 14298 7590 14310 7642
rect 14362 7590 14374 7642
rect 14426 7590 14438 7642
rect 14490 7590 18952 7642
rect 1104 7568 18952 7590
rect 37628 7642 68816 7664
rect 37628 7590 44246 7642
rect 44298 7590 44310 7642
rect 44362 7590 44374 7642
rect 44426 7590 44438 7642
rect 44490 7590 54246 7642
rect 54298 7590 54310 7642
rect 54362 7590 54374 7642
rect 54426 7590 54438 7642
rect 54490 7590 64246 7642
rect 64298 7590 64310 7642
rect 64362 7590 64374 7642
rect 64426 7590 64438 7642
rect 64490 7590 68816 7642
rect 37628 7568 68816 7590
rect 4062 7528 4068 7540
rect 2608 7500 4068 7528
rect 2608 7401 2636 7500
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7528 4215 7531
rect 6822 7528 6828 7540
rect 4203 7500 6828 7528
rect 4203 7497 4215 7500
rect 4157 7491 4215 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7006 7528 7012 7540
rect 6963 7500 7012 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 35250 7488 35256 7540
rect 35308 7528 35314 7540
rect 39666 7528 39672 7540
rect 35308 7500 39672 7528
rect 35308 7488 35314 7500
rect 39666 7488 39672 7500
rect 39724 7488 39730 7540
rect 56778 7528 56784 7540
rect 56739 7500 56784 7528
rect 56778 7488 56784 7500
rect 56836 7488 56842 7540
rect 57146 7488 57152 7540
rect 57204 7528 57210 7540
rect 57425 7531 57483 7537
rect 57425 7528 57437 7531
rect 57204 7500 57437 7528
rect 57204 7488 57210 7500
rect 57425 7497 57437 7500
rect 57471 7528 57483 7531
rect 57514 7528 57520 7540
rect 57471 7500 57520 7528
rect 57471 7497 57483 7500
rect 57425 7491 57483 7497
rect 57514 7488 57520 7500
rect 57572 7488 57578 7540
rect 57974 7528 57980 7540
rect 57935 7500 57980 7528
rect 57974 7488 57980 7500
rect 58032 7488 58038 7540
rect 60182 7528 60188 7540
rect 60143 7500 60188 7528
rect 60182 7488 60188 7500
rect 60240 7488 60246 7540
rect 60734 7488 60740 7540
rect 60792 7528 60798 7540
rect 61102 7528 61108 7540
rect 60792 7500 61108 7528
rect 60792 7488 60798 7500
rect 61102 7488 61108 7500
rect 61160 7488 61166 7540
rect 61654 7528 61660 7540
rect 61615 7500 61660 7528
rect 61654 7488 61660 7500
rect 61712 7528 61718 7540
rect 61838 7528 61844 7540
rect 61712 7500 61844 7528
rect 61712 7488 61718 7500
rect 61838 7488 61844 7500
rect 61896 7488 61902 7540
rect 17678 7460 17684 7472
rect 14936 7432 17684 7460
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 4614 7392 4620 7404
rect 2915 7364 4620 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9171 7364 14504 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 1854 7324 1860 7336
rect 1627 7296 1860 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 2498 7324 2504 7336
rect 1912 7296 2504 7324
rect 1912 7284 1918 7296
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 6972 7296 7113 7324
rect 6972 7284 6978 7296
rect 7101 7293 7113 7296
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 7466 7324 7472 7336
rect 7423 7296 7472 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10870 7324 10876 7336
rect 10468 7296 10876 7324
rect 10468 7284 10474 7296
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 12253 7327 12311 7333
rect 12253 7324 12265 7327
rect 11388 7296 12265 7324
rect 11388 7284 11394 7296
rect 12253 7293 12265 7296
rect 12299 7293 12311 7327
rect 12253 7287 12311 7293
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 12952 7296 13093 7324
rect 12952 7284 12958 7296
rect 13081 7293 13093 7296
rect 13127 7293 13139 7327
rect 13081 7287 13139 7293
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 14476 7333 14504 7364
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13320 7296 13553 7324
rect 13320 7284 13326 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 13541 7287 13599 7293
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 14936 7324 14964 7432
rect 17678 7420 17684 7432
rect 17736 7420 17742 7472
rect 35618 7420 35624 7472
rect 35676 7460 35682 7472
rect 40310 7460 40316 7472
rect 35676 7432 40316 7460
rect 35676 7420 35682 7432
rect 40310 7420 40316 7432
rect 40368 7420 40374 7472
rect 60200 7460 60228 7488
rect 61194 7460 61200 7472
rect 60200 7432 61200 7460
rect 61194 7420 61200 7432
rect 61252 7420 61258 7472
rect 16666 7392 16672 7404
rect 16408 7364 16672 7392
rect 14507 7296 14964 7324
rect 15105 7327 15163 7333
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 15286 7324 15292 7336
rect 15151 7296 15292 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15378 7284 15384 7336
rect 15436 7324 15442 7336
rect 16408 7333 16436 7364
rect 16666 7352 16672 7364
rect 16724 7392 16730 7404
rect 19518 7392 19524 7404
rect 16724 7364 19524 7392
rect 16724 7352 16730 7364
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 36262 7352 36268 7404
rect 36320 7392 36326 7404
rect 40126 7392 40132 7404
rect 36320 7364 40132 7392
rect 36320 7352 36326 7364
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 15436 7296 15761 7324
rect 15436 7284 15442 7296
rect 15749 7293 15761 7296
rect 15795 7324 15807 7327
rect 16393 7327 16451 7333
rect 15795 7296 16344 7324
rect 15795 7293 15807 7296
rect 15749 7287 15807 7293
rect 6270 7216 6276 7268
rect 6328 7256 6334 7268
rect 7285 7259 7343 7265
rect 7285 7256 7297 7259
rect 6328 7228 7297 7256
rect 6328 7216 6334 7228
rect 7285 7225 7297 7228
rect 7331 7225 7343 7259
rect 7285 7219 7343 7225
rect 9677 7259 9735 7265
rect 9677 7225 9689 7259
rect 9723 7256 9735 7259
rect 11422 7256 11428 7268
rect 9723 7228 11428 7256
rect 9723 7225 9735 7228
rect 9677 7219 9735 7225
rect 11422 7216 11428 7228
rect 11480 7216 11486 7268
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2222 7188 2228 7200
rect 2179 7160 2228 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4120 7160 4721 7188
rect 4120 7148 4126 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 4709 7151 4767 7157
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5442 7188 5448 7200
rect 5399 7160 5448 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5776 7160 5825 7188
rect 5776 7148 5782 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 8018 7188 8024 7200
rect 7979 7160 8024 7188
rect 5813 7151 5871 7157
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 11882 7188 11888 7200
rect 10275 7160 11888 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 16316 7188 16344 7296
rect 16393 7293 16405 7327
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 17589 7327 17647 7333
rect 17589 7293 17601 7327
rect 17635 7293 17647 7327
rect 18230 7324 18236 7336
rect 18191 7296 18236 7324
rect 17589 7287 17647 7293
rect 17604 7256 17632 7287
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 38102 7324 38108 7336
rect 38063 7296 38108 7324
rect 38102 7284 38108 7296
rect 38160 7284 38166 7336
rect 38746 7324 38752 7336
rect 38212 7296 38654 7324
rect 38707 7296 38752 7324
rect 17770 7256 17776 7268
rect 17604 7228 17776 7256
rect 17770 7216 17776 7228
rect 17828 7256 17834 7268
rect 21726 7256 21732 7268
rect 17828 7228 21732 7256
rect 17828 7216 17834 7228
rect 21726 7216 21732 7228
rect 21784 7216 21790 7268
rect 33042 7216 33048 7268
rect 33100 7256 33106 7268
rect 38212 7256 38240 7296
rect 33100 7228 38240 7256
rect 38626 7256 38654 7296
rect 38746 7284 38752 7296
rect 38804 7284 38810 7336
rect 40052 7333 40080 7364
rect 40126 7352 40132 7364
rect 40184 7352 40190 7404
rect 40328 7364 41460 7392
rect 40328 7336 40356 7364
rect 39393 7327 39451 7333
rect 39393 7293 39405 7327
rect 39439 7293 39451 7327
rect 39393 7287 39451 7293
rect 40037 7327 40095 7333
rect 40037 7293 40049 7327
rect 40083 7293 40095 7327
rect 40037 7287 40095 7293
rect 39114 7256 39120 7268
rect 38626 7228 39120 7256
rect 33100 7216 33106 7228
rect 39114 7216 39120 7228
rect 39172 7256 39178 7268
rect 39408 7256 39436 7287
rect 40310 7284 40316 7336
rect 40368 7284 40374 7336
rect 40770 7324 40776 7336
rect 40683 7296 40776 7324
rect 40770 7284 40776 7296
rect 40828 7284 40834 7336
rect 41432 7333 41460 7364
rect 44082 7352 44088 7404
rect 44140 7392 44146 7404
rect 46382 7392 46388 7404
rect 44140 7364 46388 7392
rect 44140 7352 44146 7364
rect 41417 7327 41475 7333
rect 41417 7293 41429 7327
rect 41463 7324 41475 7327
rect 41506 7324 41512 7336
rect 41463 7296 41512 7324
rect 41463 7293 41475 7296
rect 41417 7287 41475 7293
rect 41506 7284 41512 7296
rect 41564 7284 41570 7336
rect 41690 7284 41696 7336
rect 41748 7324 41754 7336
rect 42245 7327 42303 7333
rect 42245 7324 42257 7327
rect 41748 7296 42257 7324
rect 41748 7284 41754 7296
rect 42245 7293 42257 7296
rect 42291 7324 42303 7327
rect 43070 7324 43076 7336
rect 42291 7296 43076 7324
rect 42291 7293 42303 7296
rect 42245 7287 42303 7293
rect 43070 7284 43076 7296
rect 43128 7284 43134 7336
rect 43346 7324 43352 7336
rect 43307 7296 43352 7324
rect 43346 7284 43352 7296
rect 43404 7284 43410 7336
rect 44177 7327 44235 7333
rect 44177 7293 44189 7327
rect 44223 7324 44235 7327
rect 44726 7324 44732 7336
rect 44223 7296 44732 7324
rect 44223 7293 44235 7296
rect 44177 7287 44235 7293
rect 44726 7284 44732 7296
rect 44784 7284 44790 7336
rect 45480 7333 45508 7364
rect 46382 7352 46388 7364
rect 46440 7352 46446 7404
rect 65242 7352 65248 7404
rect 65300 7392 65306 7404
rect 69290 7392 69296 7404
rect 65300 7364 69296 7392
rect 65300 7352 65306 7364
rect 44821 7327 44879 7333
rect 44821 7293 44833 7327
rect 44867 7293 44879 7327
rect 44821 7287 44879 7293
rect 45465 7327 45523 7333
rect 45465 7293 45477 7327
rect 45511 7293 45523 7327
rect 45465 7287 45523 7293
rect 47121 7327 47179 7333
rect 47121 7293 47133 7327
rect 47167 7324 47179 7327
rect 47578 7324 47584 7336
rect 47167 7296 47584 7324
rect 47167 7293 47179 7296
rect 47121 7287 47179 7293
rect 39172 7228 39436 7256
rect 39172 7216 39178 7228
rect 40126 7216 40132 7268
rect 40184 7256 40190 7268
rect 40788 7256 40816 7284
rect 40184 7228 40816 7256
rect 40184 7216 40190 7228
rect 44358 7216 44364 7268
rect 44416 7256 44422 7268
rect 44836 7256 44864 7287
rect 47578 7284 47584 7296
rect 47636 7284 47642 7336
rect 50154 7284 50160 7336
rect 50212 7324 50218 7336
rect 65444 7333 65472 7364
rect 69290 7352 69296 7364
rect 69348 7352 69354 7404
rect 50985 7327 51043 7333
rect 50985 7324 50997 7327
rect 50212 7296 50997 7324
rect 50212 7284 50218 7296
rect 50985 7293 50997 7296
rect 51031 7293 51043 7327
rect 50985 7287 51043 7293
rect 65429 7327 65487 7333
rect 65429 7293 65441 7327
rect 65475 7293 65487 7327
rect 65429 7287 65487 7293
rect 65978 7284 65984 7336
rect 66036 7324 66042 7336
rect 66073 7327 66131 7333
rect 66073 7324 66085 7327
rect 66036 7296 66085 7324
rect 66036 7284 66042 7296
rect 66073 7293 66085 7296
rect 66119 7293 66131 7327
rect 66073 7287 66131 7293
rect 66254 7284 66260 7336
rect 66312 7324 66318 7336
rect 66714 7324 66720 7336
rect 66312 7296 66720 7324
rect 66312 7284 66318 7296
rect 66714 7284 66720 7296
rect 66772 7284 66778 7336
rect 67177 7327 67235 7333
rect 67177 7293 67189 7327
rect 67223 7293 67235 7327
rect 67177 7287 67235 7293
rect 46106 7256 46112 7268
rect 44416 7228 46112 7256
rect 44416 7216 44422 7228
rect 46106 7216 46112 7228
rect 46164 7216 46170 7268
rect 49970 7216 49976 7268
rect 50028 7256 50034 7268
rect 51537 7259 51595 7265
rect 51537 7256 51549 7259
rect 50028 7228 51549 7256
rect 50028 7216 50034 7228
rect 51537 7225 51549 7228
rect 51583 7225 51595 7259
rect 51537 7219 51595 7225
rect 51718 7216 51724 7268
rect 51776 7256 51782 7268
rect 52641 7259 52699 7265
rect 52641 7256 52653 7259
rect 51776 7228 52653 7256
rect 51776 7216 51782 7228
rect 52641 7225 52653 7228
rect 52687 7225 52699 7259
rect 52641 7219 52699 7225
rect 53834 7216 53840 7268
rect 53892 7256 53898 7268
rect 54573 7259 54631 7265
rect 54573 7256 54585 7259
rect 53892 7228 54585 7256
rect 53892 7216 53898 7228
rect 54573 7225 54585 7228
rect 54619 7225 54631 7259
rect 66990 7256 66996 7268
rect 54573 7219 54631 7225
rect 66732 7228 66996 7256
rect 66732 7200 66760 7228
rect 66990 7216 66996 7228
rect 67048 7256 67054 7268
rect 67192 7256 67220 7287
rect 67818 7284 67824 7336
rect 67876 7324 67882 7336
rect 67913 7327 67971 7333
rect 67913 7324 67925 7327
rect 67876 7296 67925 7324
rect 67876 7284 67882 7296
rect 67913 7293 67925 7296
rect 67959 7293 67971 7327
rect 67913 7287 67971 7293
rect 68094 7256 68100 7268
rect 67048 7228 67220 7256
rect 68055 7228 68100 7256
rect 67048 7216 67054 7228
rect 68094 7216 68100 7228
rect 68152 7216 68158 7268
rect 19426 7188 19432 7200
rect 16316 7160 19432 7188
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 32490 7148 32496 7200
rect 32548 7188 32554 7200
rect 38746 7188 38752 7200
rect 32548 7160 38752 7188
rect 32548 7148 32554 7160
rect 38746 7148 38752 7160
rect 38804 7148 38810 7200
rect 40770 7148 40776 7200
rect 40828 7188 40834 7200
rect 41230 7188 41236 7200
rect 40828 7160 41236 7188
rect 40828 7148 40834 7160
rect 41230 7148 41236 7160
rect 41288 7148 41294 7200
rect 45922 7188 45928 7200
rect 45883 7160 45928 7188
rect 45922 7148 45928 7160
rect 45980 7148 45986 7200
rect 46382 7148 46388 7200
rect 46440 7188 46446 7200
rect 46477 7191 46535 7197
rect 46477 7188 46489 7191
rect 46440 7160 46489 7188
rect 46440 7148 46446 7160
rect 46477 7157 46489 7160
rect 46523 7157 46535 7191
rect 46477 7151 46535 7157
rect 47394 7148 47400 7200
rect 47452 7188 47458 7200
rect 47581 7191 47639 7197
rect 47581 7188 47593 7191
rect 47452 7160 47593 7188
rect 47452 7148 47458 7160
rect 47581 7157 47593 7160
rect 47627 7157 47639 7191
rect 48222 7188 48228 7200
rect 48183 7160 48228 7188
rect 47581 7151 47639 7157
rect 48222 7148 48228 7160
rect 48280 7148 48286 7200
rect 48869 7191 48927 7197
rect 48869 7157 48881 7191
rect 48915 7188 48927 7191
rect 48958 7188 48964 7200
rect 48915 7160 48964 7188
rect 48915 7157 48927 7160
rect 48869 7151 48927 7157
rect 48958 7148 48964 7160
rect 49016 7148 49022 7200
rect 49142 7148 49148 7200
rect 49200 7188 49206 7200
rect 49329 7191 49387 7197
rect 49329 7188 49341 7191
rect 49200 7160 49341 7188
rect 49200 7148 49206 7160
rect 49329 7157 49341 7160
rect 49375 7157 49387 7191
rect 49878 7188 49884 7200
rect 49839 7160 49884 7188
rect 49329 7151 49387 7157
rect 49878 7148 49884 7160
rect 49936 7148 49942 7200
rect 50525 7191 50583 7197
rect 50525 7157 50537 7191
rect 50571 7188 50583 7191
rect 50798 7188 50804 7200
rect 50571 7160 50804 7188
rect 50571 7157 50583 7160
rect 50525 7151 50583 7157
rect 50798 7148 50804 7160
rect 50856 7148 50862 7200
rect 52178 7188 52184 7200
rect 52139 7160 52184 7188
rect 52178 7148 52184 7160
rect 52236 7148 52242 7200
rect 52914 7148 52920 7200
rect 52972 7188 52978 7200
rect 53469 7191 53527 7197
rect 53469 7188 53481 7191
rect 52972 7160 53481 7188
rect 52972 7148 52978 7160
rect 53469 7157 53481 7160
rect 53515 7157 53527 7191
rect 53469 7151 53527 7157
rect 53742 7148 53748 7200
rect 53800 7188 53806 7200
rect 54021 7191 54079 7197
rect 54021 7188 54033 7191
rect 53800 7160 54033 7188
rect 53800 7148 53806 7160
rect 54021 7157 54033 7160
rect 54067 7157 54079 7191
rect 54021 7151 54079 7157
rect 55030 7148 55036 7200
rect 55088 7188 55094 7200
rect 55217 7191 55275 7197
rect 55217 7188 55229 7191
rect 55088 7160 55229 7188
rect 55088 7148 55094 7160
rect 55217 7157 55229 7160
rect 55263 7157 55275 7191
rect 55217 7151 55275 7157
rect 55490 7148 55496 7200
rect 55548 7188 55554 7200
rect 55677 7191 55735 7197
rect 55677 7188 55689 7191
rect 55548 7160 55689 7188
rect 55548 7148 55554 7160
rect 55677 7157 55689 7160
rect 55723 7157 55735 7191
rect 56226 7188 56232 7200
rect 56187 7160 56232 7188
rect 55677 7151 55735 7157
rect 56226 7148 56232 7160
rect 56284 7148 56290 7200
rect 59538 7148 59544 7200
rect 59596 7188 59602 7200
rect 59633 7191 59691 7197
rect 59633 7188 59645 7191
rect 59596 7160 59645 7188
rect 59596 7148 59602 7160
rect 59633 7157 59645 7160
rect 59679 7157 59691 7191
rect 59633 7151 59691 7157
rect 62301 7191 62359 7197
rect 62301 7157 62313 7191
rect 62347 7188 62359 7191
rect 62390 7188 62396 7200
rect 62347 7160 62396 7188
rect 62347 7157 62359 7160
rect 62301 7151 62359 7157
rect 62390 7148 62396 7160
rect 62448 7148 62454 7200
rect 62758 7188 62764 7200
rect 62719 7160 62764 7188
rect 62758 7148 62764 7160
rect 62816 7148 62822 7200
rect 63310 7188 63316 7200
rect 63271 7160 63316 7188
rect 63310 7148 63316 7160
rect 63368 7148 63374 7200
rect 63494 7148 63500 7200
rect 63552 7188 63558 7200
rect 63957 7191 64015 7197
rect 63957 7188 63969 7191
rect 63552 7160 63969 7188
rect 63552 7148 63558 7160
rect 63957 7157 63969 7160
rect 64003 7157 64015 7191
rect 64782 7188 64788 7200
rect 64743 7160 64788 7188
rect 63957 7151 64015 7157
rect 64782 7148 64788 7160
rect 64840 7148 64846 7200
rect 66714 7148 66720 7200
rect 66772 7148 66778 7200
rect 1104 7098 18952 7120
rect 1104 7046 9246 7098
rect 9298 7046 9310 7098
rect 9362 7046 9374 7098
rect 9426 7046 9438 7098
rect 9490 7046 18952 7098
rect 1104 7024 18952 7046
rect 37628 7098 68816 7120
rect 37628 7046 39246 7098
rect 39298 7046 39310 7098
rect 39362 7046 39374 7098
rect 39426 7046 39438 7098
rect 39490 7046 49246 7098
rect 49298 7046 49310 7098
rect 49362 7046 49374 7098
rect 49426 7046 49438 7098
rect 49490 7046 59246 7098
rect 59298 7046 59310 7098
rect 59362 7046 59374 7098
rect 59426 7046 59438 7098
rect 59490 7046 68816 7098
rect 37628 7024 68816 7046
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 13078 6984 13084 6996
rect 12216 6956 13084 6984
rect 12216 6944 12222 6956
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 31754 6944 31760 6996
rect 31812 6984 31818 6996
rect 40310 6984 40316 6996
rect 31812 6956 40316 6984
rect 31812 6944 31818 6956
rect 40310 6944 40316 6956
rect 40368 6944 40374 6996
rect 41414 6944 41420 6996
rect 41472 6984 41478 6996
rect 44358 6984 44364 6996
rect 41472 6956 44364 6984
rect 41472 6944 41478 6956
rect 44358 6944 44364 6956
rect 44416 6944 44422 6996
rect 62482 6944 62488 6996
rect 62540 6984 62546 6996
rect 67818 6984 67824 6996
rect 62540 6956 67824 6984
rect 62540 6944 62546 6956
rect 67818 6944 67824 6956
rect 67876 6944 67882 6996
rect 38470 6876 38476 6928
rect 38528 6916 38534 6928
rect 40126 6916 40132 6928
rect 38528 6888 40132 6916
rect 38528 6876 38534 6888
rect 40126 6876 40132 6888
rect 40184 6876 40190 6928
rect 43162 6916 43168 6928
rect 42812 6888 43168 6916
rect 1578 6848 1584 6860
rect 1491 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6848 1642 6860
rect 2041 6851 2099 6857
rect 2041 6848 2053 6851
rect 1636 6820 2053 6848
rect 1636 6808 1642 6820
rect 2041 6817 2053 6820
rect 2087 6817 2099 6851
rect 10226 6848 10232 6860
rect 10187 6820 10232 6848
rect 2041 6811 2099 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 11149 6851 11207 6857
rect 11149 6817 11161 6851
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11164 6780 11192 6811
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11664 6820 11805 6848
rect 11664 6808 11670 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12897 6851 12955 6857
rect 12492 6820 12537 6848
rect 12492 6808 12498 6820
rect 12897 6817 12909 6851
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 11974 6780 11980 6792
rect 11164 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 12912 6780 12940 6811
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13780 6820 13829 6848
rect 13780 6808 13786 6820
rect 13817 6817 13829 6820
rect 13863 6817 13875 6851
rect 15378 6848 15384 6860
rect 15339 6820 15384 6848
rect 13817 6811 13875 6817
rect 12584 6752 12940 6780
rect 12584 6740 12590 6752
rect 2498 6672 2504 6724
rect 2556 6712 2562 6724
rect 4433 6715 4491 6721
rect 4433 6712 4445 6715
rect 2556 6684 4445 6712
rect 2556 6672 2562 6684
rect 4433 6681 4445 6684
rect 4479 6681 4491 6715
rect 4433 6675 4491 6681
rect 5994 6672 6000 6724
rect 6052 6712 6058 6724
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 6052 6684 6193 6712
rect 6052 6672 6058 6684
rect 6181 6681 6193 6684
rect 6227 6681 6239 6715
rect 13832 6712 13860 6811
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15896 6820 16037 6848
rect 15896 6808 15902 6820
rect 16025 6817 16037 6820
rect 16071 6848 16083 6851
rect 16114 6848 16120 6860
rect 16071 6820 16120 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 16632 6820 16957 6848
rect 16632 6808 16638 6820
rect 16945 6817 16957 6820
rect 16991 6817 17003 6851
rect 17586 6848 17592 6860
rect 17547 6820 17592 6848
rect 16945 6811 17003 6817
rect 16960 6780 16988 6811
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 18233 6851 18291 6857
rect 18233 6848 18245 6851
rect 18196 6820 18245 6848
rect 18196 6808 18202 6820
rect 18233 6817 18245 6820
rect 18279 6848 18291 6851
rect 19058 6848 19064 6860
rect 18279 6820 19064 6848
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 37369 6851 37427 6857
rect 37369 6817 37381 6851
rect 37415 6848 37427 6851
rect 38105 6851 38163 6857
rect 38105 6848 38117 6851
rect 37415 6820 38117 6848
rect 37415 6817 37427 6820
rect 37369 6811 37427 6817
rect 38105 6817 38117 6820
rect 38151 6817 38163 6851
rect 38562 6848 38568 6860
rect 38523 6820 38568 6848
rect 38105 6811 38163 6817
rect 22646 6780 22652 6792
rect 16960 6752 22652 6780
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 38120 6780 38148 6811
rect 38562 6808 38568 6820
rect 38620 6808 38626 6860
rect 38746 6808 38752 6860
rect 38804 6848 38810 6860
rect 39393 6851 39451 6857
rect 39393 6848 39405 6851
rect 38804 6820 39405 6848
rect 38804 6808 38810 6820
rect 39393 6817 39405 6820
rect 39439 6817 39451 6851
rect 41138 6848 41144 6860
rect 39393 6811 39451 6817
rect 39960 6820 41144 6848
rect 39850 6780 39856 6792
rect 38120 6752 39856 6780
rect 39850 6740 39856 6752
rect 39908 6740 39914 6792
rect 13832 6684 17172 6712
rect 6181 6675 6239 6681
rect 2590 6644 2596 6656
rect 2551 6616 2596 6644
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 3142 6644 3148 6656
rect 3103 6616 3148 6644
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3844 6616 3893 6644
rect 3844 6604 3850 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 5074 6644 5080 6656
rect 5035 6616 5080 6644
rect 3881 6607 3939 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5721 6647 5779 6653
rect 5721 6613 5733 6647
rect 5767 6644 5779 6647
rect 6086 6644 6092 6656
rect 5767 6616 6092 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 7650 6644 7656 6656
rect 7515 6616 7656 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 8202 6644 8208 6656
rect 8163 6616 8208 6644
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6644 9643 6647
rect 13722 6644 13728 6656
rect 9631 6616 13728 6644
rect 9631 6613 9643 6616
rect 9585 6607 9643 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 17034 6644 17040 6656
rect 14783 6616 17040 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 17144 6644 17172 6684
rect 17586 6672 17592 6724
rect 17644 6712 17650 6724
rect 20898 6712 20904 6724
rect 17644 6684 20904 6712
rect 17644 6672 17650 6684
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 36998 6672 37004 6724
rect 37056 6712 37062 6724
rect 39960 6712 39988 6820
rect 41138 6808 41144 6820
rect 41196 6848 41202 6860
rect 41325 6851 41383 6857
rect 41325 6848 41337 6851
rect 41196 6820 41337 6848
rect 41196 6808 41202 6820
rect 41325 6817 41337 6820
rect 41371 6817 41383 6851
rect 41325 6811 41383 6817
rect 41414 6808 41420 6860
rect 41472 6848 41478 6860
rect 42150 6848 42156 6860
rect 41472 6820 42156 6848
rect 41472 6808 41478 6820
rect 42150 6808 42156 6820
rect 42208 6808 42214 6860
rect 42812 6857 42840 6888
rect 43162 6876 43168 6888
rect 43220 6876 43226 6928
rect 45554 6916 45560 6928
rect 43456 6888 43668 6916
rect 42797 6851 42855 6857
rect 42797 6817 42809 6851
rect 42843 6817 42855 6851
rect 42797 6811 42855 6817
rect 42886 6808 42892 6860
rect 42944 6848 42950 6860
rect 43456 6848 43484 6888
rect 42944 6820 43484 6848
rect 43533 6851 43591 6857
rect 42944 6808 42950 6820
rect 43533 6817 43545 6851
rect 43579 6817 43591 6851
rect 43640 6848 43668 6888
rect 45296 6888 45560 6916
rect 43993 6851 44051 6857
rect 43993 6848 44005 6851
rect 43640 6820 44005 6848
rect 43533 6811 43591 6817
rect 43993 6817 44005 6820
rect 44039 6848 44051 6851
rect 44726 6848 44732 6860
rect 44039 6820 44732 6848
rect 44039 6817 44051 6820
rect 43993 6811 44051 6817
rect 40126 6740 40132 6792
rect 40184 6780 40190 6792
rect 43548 6780 43576 6811
rect 44726 6808 44732 6820
rect 44784 6808 44790 6860
rect 44821 6851 44879 6857
rect 44821 6817 44833 6851
rect 44867 6848 44879 6851
rect 45186 6848 45192 6860
rect 44867 6820 45192 6848
rect 44867 6817 44879 6820
rect 44821 6811 44879 6817
rect 44542 6780 44548 6792
rect 40184 6752 44548 6780
rect 40184 6740 40190 6752
rect 44542 6740 44548 6752
rect 44600 6740 44606 6792
rect 44836 6712 44864 6811
rect 45186 6808 45192 6820
rect 45244 6808 45250 6860
rect 37056 6684 39988 6712
rect 40052 6684 44864 6712
rect 37056 6672 37062 6684
rect 18966 6644 18972 6656
rect 17144 6616 18972 6644
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 37826 6604 37832 6656
rect 37884 6644 37890 6656
rect 40052 6644 40080 6684
rect 45186 6672 45192 6724
rect 45244 6712 45250 6724
rect 45296 6712 45324 6888
rect 45554 6876 45560 6888
rect 45612 6876 45618 6928
rect 65334 6916 65340 6928
rect 64984 6888 65340 6916
rect 45830 6808 45836 6860
rect 45888 6848 45894 6860
rect 46017 6851 46075 6857
rect 46017 6848 46029 6851
rect 45888 6820 46029 6848
rect 45888 6808 45894 6820
rect 46017 6817 46029 6820
rect 46063 6817 46075 6851
rect 46017 6811 46075 6817
rect 46661 6851 46719 6857
rect 46661 6817 46673 6851
rect 46707 6817 46719 6851
rect 47486 6848 47492 6860
rect 47447 6820 47492 6848
rect 46661 6811 46719 6817
rect 45554 6740 45560 6792
rect 45612 6780 45618 6792
rect 46566 6780 46572 6792
rect 45612 6752 46572 6780
rect 45612 6740 45618 6752
rect 46566 6740 46572 6752
rect 46624 6780 46630 6792
rect 46676 6780 46704 6811
rect 47486 6808 47492 6820
rect 47544 6808 47550 6860
rect 59357 6851 59415 6857
rect 59357 6817 59369 6851
rect 59403 6848 59415 6851
rect 59630 6848 59636 6860
rect 59403 6820 59636 6848
rect 59403 6817 59415 6820
rect 59357 6811 59415 6817
rect 59630 6808 59636 6820
rect 59688 6808 59694 6860
rect 64984 6857 65012 6888
rect 65334 6876 65340 6888
rect 65392 6916 65398 6928
rect 65392 6888 65748 6916
rect 65392 6876 65398 6888
rect 64969 6851 65027 6857
rect 64969 6817 64981 6851
rect 65015 6817 65027 6851
rect 64969 6811 65027 6817
rect 65426 6808 65432 6860
rect 65484 6848 65490 6860
rect 65613 6851 65671 6857
rect 65613 6848 65625 6851
rect 65484 6820 65625 6848
rect 65484 6808 65490 6820
rect 65613 6817 65625 6820
rect 65659 6817 65671 6851
rect 65613 6811 65671 6817
rect 46624 6752 46704 6780
rect 46624 6740 46630 6752
rect 47118 6740 47124 6792
rect 47176 6740 47182 6792
rect 47302 6740 47308 6792
rect 47360 6780 47366 6792
rect 48501 6783 48559 6789
rect 48501 6780 48513 6783
rect 47360 6752 48513 6780
rect 47360 6740 47366 6752
rect 48501 6749 48513 6752
rect 48547 6749 48559 6783
rect 48501 6743 48559 6749
rect 64138 6740 64144 6792
rect 64196 6780 64202 6792
rect 65334 6780 65340 6792
rect 64196 6752 65340 6780
rect 64196 6740 64202 6752
rect 65334 6740 65340 6752
rect 65392 6740 65398 6792
rect 65720 6780 65748 6888
rect 67266 6808 67272 6860
rect 67324 6848 67330 6860
rect 67453 6851 67511 6857
rect 67453 6848 67465 6851
rect 67324 6820 67465 6848
rect 67324 6808 67330 6820
rect 67453 6817 67465 6820
rect 67499 6817 67511 6851
rect 67453 6811 67511 6817
rect 67726 6808 67732 6860
rect 67784 6848 67790 6860
rect 67913 6851 67971 6857
rect 67913 6848 67925 6851
rect 67784 6820 67925 6848
rect 67784 6808 67790 6820
rect 67913 6817 67925 6820
rect 67959 6817 67971 6851
rect 67913 6811 67971 6817
rect 68462 6780 68468 6792
rect 65720 6752 68468 6780
rect 68462 6740 68468 6752
rect 68520 6740 68526 6792
rect 45244 6684 45324 6712
rect 45244 6672 45250 6684
rect 46106 6672 46112 6724
rect 46164 6712 46170 6724
rect 47136 6712 47164 6740
rect 46164 6684 47164 6712
rect 46164 6672 46170 6684
rect 48038 6672 48044 6724
rect 48096 6712 48102 6724
rect 49053 6715 49111 6721
rect 49053 6712 49065 6715
rect 48096 6684 49065 6712
rect 48096 6672 48102 6684
rect 49053 6681 49065 6684
rect 49099 6681 49111 6715
rect 49053 6675 49111 6681
rect 57606 6672 57612 6724
rect 57664 6712 57670 6724
rect 58345 6715 58403 6721
rect 58345 6712 58357 6715
rect 57664 6684 58357 6712
rect 57664 6672 57670 6684
rect 58345 6681 58357 6684
rect 58391 6681 58403 6715
rect 58345 6675 58403 6681
rect 64046 6672 64052 6724
rect 64104 6712 64110 6724
rect 65794 6712 65800 6724
rect 64104 6684 65800 6712
rect 64104 6672 64110 6684
rect 65794 6672 65800 6684
rect 65852 6672 65858 6724
rect 37884 6616 40080 6644
rect 37884 6604 37890 6616
rect 40310 6604 40316 6656
rect 40368 6644 40374 6656
rect 40405 6647 40463 6653
rect 40405 6644 40417 6647
rect 40368 6616 40417 6644
rect 40368 6604 40374 6616
rect 40405 6613 40417 6616
rect 40451 6613 40463 6647
rect 40405 6607 40463 6613
rect 46382 6604 46388 6656
rect 46440 6644 46446 6656
rect 46566 6644 46572 6656
rect 46440 6616 46572 6644
rect 46440 6604 46446 6616
rect 46566 6604 46572 6616
rect 46624 6604 46630 6656
rect 47118 6604 47124 6656
rect 47176 6644 47182 6656
rect 47949 6647 48007 6653
rect 47949 6644 47961 6647
rect 47176 6616 47961 6644
rect 47176 6604 47182 6616
rect 47949 6613 47961 6616
rect 47995 6613 48007 6647
rect 47949 6607 48007 6613
rect 49697 6647 49755 6653
rect 49697 6613 49709 6647
rect 49743 6644 49755 6647
rect 49786 6644 49792 6656
rect 49743 6616 49792 6644
rect 49743 6613 49755 6616
rect 49697 6607 49755 6613
rect 49786 6604 49792 6616
rect 49844 6604 49850 6656
rect 50062 6604 50068 6656
rect 50120 6644 50126 6656
rect 50157 6647 50215 6653
rect 50157 6644 50169 6647
rect 50120 6616 50169 6644
rect 50120 6604 50126 6616
rect 50157 6613 50169 6616
rect 50203 6613 50215 6647
rect 50157 6607 50215 6613
rect 50706 6604 50712 6656
rect 50764 6644 50770 6656
rect 50893 6647 50951 6653
rect 50893 6644 50905 6647
rect 50764 6616 50905 6644
rect 50764 6604 50770 6616
rect 50893 6613 50905 6616
rect 50939 6613 50951 6647
rect 50893 6607 50951 6613
rect 51258 6604 51264 6656
rect 51316 6644 51322 6656
rect 51445 6647 51503 6653
rect 51445 6644 51457 6647
rect 51316 6616 51457 6644
rect 51316 6604 51322 6616
rect 51445 6613 51457 6616
rect 51491 6613 51503 6647
rect 51445 6607 51503 6613
rect 51810 6604 51816 6656
rect 51868 6644 51874 6656
rect 51997 6647 52055 6653
rect 51997 6644 52009 6647
rect 51868 6616 52009 6644
rect 51868 6604 51874 6616
rect 51997 6613 52009 6616
rect 52043 6613 52055 6647
rect 52546 6644 52552 6656
rect 52507 6616 52552 6644
rect 51997 6607 52055 6613
rect 52546 6604 52552 6616
rect 52604 6604 52610 6656
rect 53190 6644 53196 6656
rect 53151 6616 53196 6644
rect 53190 6604 53196 6616
rect 53248 6604 53254 6656
rect 53926 6644 53932 6656
rect 53887 6616 53932 6644
rect 53926 6604 53932 6616
rect 53984 6604 53990 6656
rect 54570 6644 54576 6656
rect 54531 6616 54576 6644
rect 54570 6604 54576 6616
rect 54628 6604 54634 6656
rect 54938 6604 54944 6656
rect 54996 6644 55002 6656
rect 55033 6647 55091 6653
rect 55033 6644 55045 6647
rect 54996 6616 55045 6644
rect 54996 6604 55002 6616
rect 55033 6613 55045 6616
rect 55079 6613 55091 6647
rect 55033 6607 55091 6613
rect 55398 6604 55404 6656
rect 55456 6644 55462 6656
rect 56137 6647 56195 6653
rect 56137 6644 56149 6647
rect 55456 6616 56149 6644
rect 55456 6604 55462 6616
rect 56137 6613 56149 6616
rect 56183 6613 56195 6647
rect 56137 6607 56195 6613
rect 56318 6604 56324 6656
rect 56376 6644 56382 6656
rect 56689 6647 56747 6653
rect 56689 6644 56701 6647
rect 56376 6616 56701 6644
rect 56376 6604 56382 6616
rect 56689 6613 56701 6616
rect 56735 6613 56747 6647
rect 57238 6644 57244 6656
rect 57199 6616 57244 6644
rect 56689 6607 56747 6613
rect 57238 6604 57244 6616
rect 57296 6604 57302 6656
rect 57882 6644 57888 6656
rect 57843 6616 57888 6644
rect 57882 6604 57888 6616
rect 57940 6604 57946 6656
rect 59909 6647 59967 6653
rect 59909 6613 59921 6647
rect 59955 6644 59967 6647
rect 60182 6644 60188 6656
rect 59955 6616 60188 6644
rect 59955 6613 59967 6616
rect 59909 6607 59967 6613
rect 60182 6604 60188 6616
rect 60240 6604 60246 6656
rect 60366 6644 60372 6656
rect 60327 6616 60372 6644
rect 60366 6604 60372 6616
rect 60424 6604 60430 6656
rect 61378 6644 61384 6656
rect 61339 6616 61384 6644
rect 61378 6604 61384 6616
rect 61436 6604 61442 6656
rect 62022 6644 62028 6656
rect 61983 6616 62028 6644
rect 62022 6604 62028 6616
rect 62080 6604 62086 6656
rect 62850 6644 62856 6656
rect 62811 6616 62856 6644
rect 62850 6604 62856 6616
rect 62908 6604 62914 6656
rect 63402 6644 63408 6656
rect 63363 6616 63408 6644
rect 63402 6604 63408 6616
rect 63460 6604 63466 6656
rect 64138 6644 64144 6656
rect 64099 6616 64144 6644
rect 64138 6604 64144 6616
rect 64196 6604 64202 6656
rect 66809 6647 66867 6653
rect 66809 6613 66821 6647
rect 66855 6644 66867 6647
rect 67542 6644 67548 6656
rect 66855 6616 67548 6644
rect 66855 6613 66867 6616
rect 66809 6607 66867 6613
rect 67542 6604 67548 6616
rect 67600 6604 67606 6656
rect 1104 6554 18952 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 14246 6554
rect 14298 6502 14310 6554
rect 14362 6502 14374 6554
rect 14426 6502 14438 6554
rect 14490 6502 18952 6554
rect 1104 6480 18952 6502
rect 37628 6554 68816 6576
rect 37628 6502 44246 6554
rect 44298 6502 44310 6554
rect 44362 6502 44374 6554
rect 44426 6502 44438 6554
rect 44490 6502 54246 6554
rect 54298 6502 54310 6554
rect 54362 6502 54374 6554
rect 54426 6502 54438 6554
rect 54490 6502 64246 6554
rect 64298 6502 64310 6554
rect 64362 6502 64374 6554
rect 64426 6502 64438 6554
rect 64490 6502 68816 6554
rect 37628 6480 68816 6502
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 16298 6440 16304 6452
rect 15436 6412 16304 6440
rect 15436 6400 15442 6412
rect 16298 6400 16304 6412
rect 16356 6440 16362 6452
rect 20438 6440 20444 6452
rect 16356 6412 20444 6440
rect 16356 6400 16362 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 39577 6443 39635 6449
rect 39577 6409 39589 6443
rect 39623 6440 39635 6443
rect 39758 6440 39764 6452
rect 39623 6412 39764 6440
rect 39623 6409 39635 6412
rect 39577 6403 39635 6409
rect 39758 6400 39764 6412
rect 39816 6400 39822 6452
rect 39850 6400 39856 6452
rect 39908 6440 39914 6452
rect 40037 6443 40095 6449
rect 40037 6440 40049 6443
rect 39908 6412 40049 6440
rect 39908 6400 39914 6412
rect 40037 6409 40049 6412
rect 40083 6409 40095 6443
rect 45646 6440 45652 6452
rect 40037 6403 40095 6409
rect 40236 6412 45652 6440
rect 22554 6372 22560 6384
rect 16408 6344 22560 6372
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 7006 6304 7012 6316
rect 5132 6276 7012 6304
rect 5132 6264 5138 6276
rect 7006 6264 7012 6276
rect 7064 6304 7070 6316
rect 16114 6304 16120 6316
rect 7064 6276 8616 6304
rect 7064 6264 7070 6276
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 1728 6208 2053 6236
rect 1728 6196 1734 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 8588 6245 8616 6276
rect 15120 6276 16120 6304
rect 3145 6239 3203 6245
rect 3145 6236 3157 6239
rect 3016 6208 3157 6236
rect 3016 6196 3022 6208
rect 3145 6205 3157 6208
rect 3191 6205 3203 6239
rect 3145 6199 3203 6205
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 9180 6208 9413 6236
rect 9180 6196 9186 6208
rect 9401 6205 9413 6208
rect 9447 6236 9459 6239
rect 9582 6236 9588 6248
rect 9447 6208 9588 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9824 6208 9873 6236
rect 9824 6196 9830 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 11112 6208 11161 6236
rect 11112 6196 11118 6208
rect 11149 6205 11161 6208
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 13170 6236 13176 6248
rect 13131 6208 13176 6236
rect 12529 6199 12587 6205
rect 4249 6171 4307 6177
rect 4249 6137 4261 6171
rect 4295 6168 4307 6171
rect 5074 6168 5080 6180
rect 4295 6140 5080 6168
rect 4295 6137 4307 6140
rect 4249 6131 4307 6137
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 7377 6171 7435 6177
rect 7377 6137 7389 6171
rect 7423 6168 7435 6171
rect 12544 6168 12572 6199
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6205 13875 6239
rect 14458 6236 14464 6248
rect 14419 6208 14464 6236
rect 13817 6199 13875 6205
rect 13630 6168 13636 6180
rect 7423 6140 13636 6168
rect 7423 6137 7435 6140
rect 7377 6131 7435 6137
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 13832 6168 13860 6199
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 15120 6245 15148 6276
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6205 15163 6239
rect 15105 6199 15163 6205
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 15749 6239 15807 6245
rect 15749 6236 15761 6239
rect 15620 6208 15761 6236
rect 15620 6196 15626 6208
rect 15749 6205 15761 6208
rect 15795 6236 15807 6239
rect 16206 6236 16212 6248
rect 15795 6208 16212 6236
rect 15795 6205 15807 6208
rect 15749 6199 15807 6205
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 16298 6196 16304 6248
rect 16356 6236 16362 6248
rect 16408 6245 16436 6344
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 36538 6332 36544 6384
rect 36596 6372 36602 6384
rect 40236 6372 40264 6412
rect 45646 6400 45652 6412
rect 45704 6400 45710 6452
rect 42794 6372 42800 6384
rect 36596 6344 40264 6372
rect 40328 6344 42800 6372
rect 36596 6332 36602 6344
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 19150 6304 19156 6316
rect 16908 6276 19156 6304
rect 16908 6264 16914 6276
rect 17604 6245 17632 6276
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 35526 6264 35532 6316
rect 35584 6304 35590 6316
rect 37918 6304 37924 6316
rect 35584 6276 37504 6304
rect 37879 6276 37924 6304
rect 35584 6264 35590 6276
rect 16393 6239 16451 6245
rect 16393 6236 16405 6239
rect 16356 6208 16405 6236
rect 16356 6196 16362 6208
rect 16393 6205 16405 6208
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 19334 6236 19340 6248
rect 18279 6208 19340 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 19334 6196 19340 6208
rect 19392 6236 19398 6248
rect 19886 6236 19892 6248
rect 19392 6208 19892 6236
rect 19392 6196 19398 6208
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 31573 6239 31631 6245
rect 31573 6205 31585 6239
rect 31619 6236 31631 6239
rect 37369 6239 37427 6245
rect 37369 6236 37381 6239
rect 31619 6208 37381 6236
rect 31619 6205 31631 6208
rect 31573 6199 31631 6205
rect 37369 6205 37381 6208
rect 37415 6205 37427 6239
rect 37476 6236 37504 6276
rect 37918 6264 37924 6276
rect 37976 6264 37982 6316
rect 38749 6307 38807 6313
rect 38749 6273 38761 6307
rect 38795 6304 38807 6307
rect 39850 6304 39856 6316
rect 38795 6276 39856 6304
rect 38795 6273 38807 6276
rect 38749 6267 38807 6273
rect 39850 6264 39856 6276
rect 39908 6264 39914 6316
rect 40328 6236 40356 6344
rect 42794 6332 42800 6344
rect 42852 6332 42858 6384
rect 47210 6372 47216 6384
rect 46124 6344 47216 6372
rect 44174 6264 44180 6316
rect 44232 6304 44238 6316
rect 46124 6304 46152 6344
rect 47210 6332 47216 6344
rect 47268 6332 47274 6384
rect 48777 6307 48835 6313
rect 48777 6304 48789 6307
rect 44232 6276 46152 6304
rect 44232 6264 44238 6276
rect 40681 6239 40739 6245
rect 40681 6236 40693 6239
rect 37476 6208 40356 6236
rect 40420 6208 40693 6236
rect 37369 6199 37427 6205
rect 14090 6168 14096 6180
rect 13832 6140 14096 6168
rect 14090 6128 14096 6140
rect 14148 6168 14154 6180
rect 23382 6168 23388 6180
rect 14148 6140 23388 6168
rect 14148 6128 14154 6140
rect 23382 6128 23388 6140
rect 23440 6128 23446 6180
rect 35342 6128 35348 6180
rect 35400 6168 35406 6180
rect 40420 6168 40448 6208
rect 40681 6205 40693 6208
rect 40727 6236 40739 6239
rect 40862 6236 40868 6248
rect 40727 6208 40868 6236
rect 40727 6205 40739 6208
rect 40681 6199 40739 6205
rect 40862 6196 40868 6208
rect 40920 6196 40926 6248
rect 41417 6239 41475 6245
rect 41417 6205 41429 6239
rect 41463 6236 41475 6239
rect 41598 6236 41604 6248
rect 41463 6208 41604 6236
rect 41463 6205 41475 6208
rect 41417 6199 41475 6205
rect 41432 6168 41460 6199
rect 41598 6196 41604 6208
rect 41656 6196 41662 6248
rect 42058 6236 42064 6248
rect 42019 6208 42064 6236
rect 42058 6196 42064 6208
rect 42116 6196 42122 6248
rect 43070 6196 43076 6248
rect 43128 6236 43134 6248
rect 43349 6239 43407 6245
rect 43349 6236 43361 6239
rect 43128 6208 43361 6236
rect 43128 6196 43134 6208
rect 43349 6205 43361 6208
rect 43395 6236 43407 6239
rect 43438 6236 43444 6248
rect 43395 6208 43444 6236
rect 43395 6205 43407 6208
rect 43349 6199 43407 6205
rect 43438 6196 43444 6208
rect 43496 6196 43502 6248
rect 43993 6239 44051 6245
rect 43993 6205 44005 6239
rect 44039 6205 44051 6239
rect 43993 6199 44051 6205
rect 35400 6140 40448 6168
rect 40604 6140 41460 6168
rect 35400 6128 35406 6140
rect 3602 6100 3608 6112
rect 3563 6072 3608 6100
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4672 6072 4721 6100
rect 4672 6060 4678 6072
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 4709 6063 4767 6069
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 5261 6103 5319 6109
rect 5261 6100 5273 6103
rect 5040 6072 5273 6100
rect 5040 6060 5046 6072
rect 5261 6069 5273 6072
rect 5307 6069 5319 6103
rect 5261 6063 5319 6069
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 5813 6103 5871 6109
rect 5813 6100 5825 6103
rect 5776 6072 5825 6100
rect 5776 6060 5782 6072
rect 5813 6069 5825 6072
rect 5859 6069 5871 6103
rect 6730 6100 6736 6112
rect 6691 6072 6736 6100
rect 5813 6063 5871 6069
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 10870 6100 10876 6112
rect 7975 6072 10876 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11885 6103 11943 6109
rect 11885 6069 11897 6103
rect 11931 6100 11943 6103
rect 16574 6100 16580 6112
rect 11931 6072 16580 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 35434 6060 35440 6112
rect 35492 6100 35498 6112
rect 40604 6100 40632 6140
rect 42978 6128 42984 6180
rect 43036 6168 43042 6180
rect 43806 6168 43812 6180
rect 43036 6140 43812 6168
rect 43036 6128 43042 6140
rect 43806 6128 43812 6140
rect 43864 6168 43870 6180
rect 44008 6168 44036 6199
rect 44726 6196 44732 6248
rect 44784 6236 44790 6248
rect 44821 6239 44879 6245
rect 44821 6236 44833 6239
rect 44784 6208 44833 6236
rect 44784 6196 44790 6208
rect 44821 6205 44833 6208
rect 44867 6205 44879 6239
rect 44821 6199 44879 6205
rect 45465 6239 45523 6245
rect 45465 6205 45477 6239
rect 45511 6236 45523 6239
rect 45646 6236 45652 6248
rect 45511 6208 45652 6236
rect 45511 6205 45523 6208
rect 45465 6199 45523 6205
rect 43864 6140 44036 6168
rect 44836 6168 44864 6199
rect 45646 6196 45652 6208
rect 45704 6196 45710 6248
rect 46124 6245 46152 6276
rect 46216 6276 48789 6304
rect 46109 6239 46167 6245
rect 46109 6205 46121 6239
rect 46155 6205 46167 6239
rect 46109 6199 46167 6205
rect 46216 6168 46244 6276
rect 48777 6273 48789 6276
rect 48823 6273 48835 6307
rect 48777 6267 48835 6273
rect 46753 6239 46811 6245
rect 46753 6205 46765 6239
rect 46799 6205 46811 6239
rect 46753 6199 46811 6205
rect 44836 6140 46244 6168
rect 46768 6168 46796 6199
rect 47026 6196 47032 6248
rect 47084 6236 47090 6248
rect 47213 6239 47271 6245
rect 47213 6236 47225 6239
rect 47084 6208 47225 6236
rect 47084 6196 47090 6208
rect 47213 6205 47225 6208
rect 47259 6205 47271 6239
rect 47213 6199 47271 6205
rect 49970 6196 49976 6248
rect 50028 6236 50034 6248
rect 50249 6239 50307 6245
rect 50249 6236 50261 6239
rect 50028 6208 50261 6236
rect 50028 6196 50034 6208
rect 50249 6205 50261 6208
rect 50295 6205 50307 6239
rect 50890 6236 50896 6248
rect 50851 6208 50896 6236
rect 50249 6199 50307 6205
rect 50890 6196 50896 6208
rect 50948 6196 50954 6248
rect 51997 6239 52055 6245
rect 51997 6205 52009 6239
rect 52043 6236 52055 6239
rect 55858 6236 55864 6248
rect 52043 6208 55864 6236
rect 52043 6205 52055 6208
rect 51997 6199 52055 6205
rect 55858 6196 55864 6208
rect 55916 6196 55922 6248
rect 64690 6196 64696 6248
rect 64748 6236 64754 6248
rect 64785 6239 64843 6245
rect 64785 6236 64797 6239
rect 64748 6208 64797 6236
rect 64748 6196 64754 6208
rect 64785 6205 64797 6208
rect 64831 6205 64843 6239
rect 64785 6199 64843 6205
rect 65058 6196 65064 6248
rect 65116 6236 65122 6248
rect 65245 6239 65303 6245
rect 65245 6236 65257 6239
rect 65116 6208 65257 6236
rect 65116 6196 65122 6208
rect 65245 6205 65257 6208
rect 65291 6205 65303 6239
rect 65245 6199 65303 6205
rect 66438 6196 66444 6248
rect 66496 6236 66502 6248
rect 66625 6239 66683 6245
rect 66625 6236 66637 6239
rect 66496 6208 66637 6236
rect 66496 6196 66502 6208
rect 66625 6205 66637 6208
rect 66671 6205 66683 6239
rect 66625 6199 66683 6205
rect 66898 6196 66904 6248
rect 66956 6236 66962 6248
rect 67082 6236 67088 6248
rect 66956 6208 67088 6236
rect 66956 6196 66962 6208
rect 67082 6196 67088 6208
rect 67140 6196 67146 6248
rect 67542 6196 67548 6248
rect 67600 6236 67606 6248
rect 68097 6239 68155 6245
rect 68097 6236 68109 6239
rect 67600 6208 68109 6236
rect 67600 6196 67606 6208
rect 68097 6205 68109 6208
rect 68143 6205 68155 6239
rect 68097 6199 68155 6205
rect 47854 6168 47860 6180
rect 46768 6140 47860 6168
rect 43864 6128 43870 6140
rect 35492 6072 40632 6100
rect 35492 6060 35498 6072
rect 41138 6060 41144 6112
rect 41196 6100 41202 6112
rect 46768 6100 46796 6140
rect 47854 6128 47860 6140
rect 47912 6128 47918 6180
rect 47946 6128 47952 6180
rect 48004 6168 48010 6180
rect 49329 6171 49387 6177
rect 49329 6168 49341 6171
rect 48004 6140 49341 6168
rect 48004 6128 48010 6140
rect 49329 6137 49341 6140
rect 49375 6137 49387 6171
rect 49329 6131 49387 6137
rect 56410 6128 56416 6180
rect 56468 6168 56474 6180
rect 58069 6171 58127 6177
rect 58069 6168 58081 6171
rect 56468 6140 58081 6168
rect 56468 6128 56474 6140
rect 58069 6137 58081 6140
rect 58115 6137 58127 6171
rect 58069 6131 58127 6137
rect 59906 6128 59912 6180
rect 59964 6168 59970 6180
rect 60737 6171 60795 6177
rect 60737 6168 60749 6171
rect 59964 6140 60749 6168
rect 59964 6128 59970 6140
rect 60737 6137 60749 6140
rect 60783 6137 60795 6171
rect 60737 6131 60795 6137
rect 41196 6072 46796 6100
rect 41196 6060 41202 6072
rect 46934 6060 46940 6112
rect 46992 6100 46998 6112
rect 48225 6103 48283 6109
rect 48225 6100 48237 6103
rect 46992 6072 48237 6100
rect 46992 6060 46998 6072
rect 48225 6069 48237 6072
rect 48271 6069 48283 6103
rect 48225 6063 48283 6069
rect 52549 6103 52607 6109
rect 52549 6069 52561 6103
rect 52595 6100 52607 6103
rect 52638 6100 52644 6112
rect 52595 6072 52644 6100
rect 52595 6069 52607 6072
rect 52549 6063 52607 6069
rect 52638 6060 52644 6072
rect 52696 6060 52702 6112
rect 53282 6060 53288 6112
rect 53340 6100 53346 6112
rect 53653 6103 53711 6109
rect 53653 6100 53665 6103
rect 53340 6072 53665 6100
rect 53340 6060 53346 6072
rect 53653 6069 53665 6072
rect 53699 6069 53711 6103
rect 53653 6063 53711 6069
rect 54389 6103 54447 6109
rect 54389 6069 54401 6103
rect 54435 6100 54447 6103
rect 54754 6100 54760 6112
rect 54435 6072 54760 6100
rect 54435 6069 54447 6072
rect 54389 6063 54447 6069
rect 54754 6060 54760 6072
rect 54812 6060 54818 6112
rect 55033 6103 55091 6109
rect 55033 6069 55045 6103
rect 55079 6100 55091 6103
rect 55122 6100 55128 6112
rect 55079 6072 55128 6100
rect 55079 6069 55091 6072
rect 55033 6063 55091 6069
rect 55122 6060 55128 6072
rect 55180 6060 55186 6112
rect 55582 6100 55588 6112
rect 55543 6072 55588 6100
rect 55582 6060 55588 6072
rect 55640 6060 55646 6112
rect 56134 6100 56140 6112
rect 56095 6072 56140 6100
rect 56134 6060 56140 6072
rect 56192 6060 56198 6112
rect 56870 6060 56876 6112
rect 56928 6100 56934 6112
rect 56965 6103 57023 6109
rect 56965 6100 56977 6103
rect 56928 6072 56977 6100
rect 56928 6060 56934 6072
rect 56965 6069 56977 6072
rect 57011 6069 57023 6103
rect 57514 6100 57520 6112
rect 57475 6072 57520 6100
rect 56965 6063 57023 6069
rect 57514 6060 57520 6072
rect 57572 6060 57578 6112
rect 58894 6100 58900 6112
rect 58855 6072 58900 6100
rect 58894 6060 58900 6072
rect 58952 6060 58958 6112
rect 59633 6103 59691 6109
rect 59633 6069 59645 6103
rect 59679 6100 59691 6103
rect 59814 6100 59820 6112
rect 59679 6072 59820 6100
rect 59679 6069 59691 6072
rect 59633 6063 59691 6069
rect 59814 6060 59820 6072
rect 59872 6060 59878 6112
rect 60090 6100 60096 6112
rect 60051 6072 60096 6100
rect 60090 6060 60096 6072
rect 60148 6060 60154 6112
rect 61654 6100 61660 6112
rect 61615 6072 61660 6100
rect 61654 6060 61660 6072
rect 61712 6060 61718 6112
rect 62298 6100 62304 6112
rect 62259 6072 62304 6100
rect 62298 6060 62304 6072
rect 62356 6060 62362 6112
rect 62945 6103 63003 6109
rect 62945 6069 62957 6103
rect 62991 6100 63003 6103
rect 63218 6100 63224 6112
rect 62991 6072 63224 6100
rect 62991 6069 63003 6072
rect 62945 6063 63003 6069
rect 63218 6060 63224 6072
rect 63276 6060 63282 6112
rect 63678 6060 63684 6112
rect 63736 6100 63742 6112
rect 64049 6103 64107 6109
rect 64049 6100 64061 6103
rect 63736 6072 64061 6100
rect 63736 6060 63742 6072
rect 64049 6069 64061 6072
rect 64095 6069 64107 6103
rect 64049 6063 64107 6069
rect 64506 6060 64512 6112
rect 64564 6100 64570 6112
rect 65889 6103 65947 6109
rect 65889 6100 65901 6103
rect 64564 6072 65901 6100
rect 64564 6060 64570 6072
rect 65889 6069 65901 6072
rect 65935 6069 65947 6103
rect 65889 6063 65947 6069
rect 1104 6010 18952 6032
rect 1104 5958 9246 6010
rect 9298 5958 9310 6010
rect 9362 5958 9374 6010
rect 9426 5958 9438 6010
rect 9490 5958 18952 6010
rect 1104 5936 18952 5958
rect 37628 6010 68816 6032
rect 37628 5958 39246 6010
rect 39298 5958 39310 6010
rect 39362 5958 39374 6010
rect 39426 5958 39438 6010
rect 39490 5958 49246 6010
rect 49298 5958 49310 6010
rect 49362 5958 49374 6010
rect 49426 5958 49438 6010
rect 49490 5958 59246 6010
rect 59298 5958 59310 6010
rect 59362 5958 59374 6010
rect 59426 5958 59438 6010
rect 59490 5958 68816 6010
rect 37628 5936 68816 5958
rect 10042 5856 10048 5908
rect 10100 5856 10106 5908
rect 13354 5896 13360 5908
rect 13188 5868 13360 5896
rect 1762 5828 1768 5840
rect 1723 5800 1768 5828
rect 1762 5788 1768 5800
rect 1820 5788 1826 5840
rect 1949 5831 2007 5837
rect 1949 5797 1961 5831
rect 1995 5828 2007 5831
rect 2774 5828 2780 5840
rect 1995 5800 2780 5828
rect 1995 5797 2007 5800
rect 1949 5791 2007 5797
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 2038 5720 2044 5772
rect 2096 5760 2102 5772
rect 2682 5760 2688 5772
rect 2096 5732 2688 5760
rect 2096 5720 2102 5732
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 3326 5760 3332 5772
rect 3287 5732 3332 5760
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 4948 5732 5089 5760
rect 4948 5720 4954 5732
rect 5077 5729 5089 5732
rect 5123 5729 5135 5763
rect 5077 5723 5135 5729
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 5721 5763 5779 5769
rect 5721 5760 5733 5763
rect 5592 5732 5733 5760
rect 5592 5720 5598 5732
rect 5721 5729 5733 5732
rect 5767 5729 5779 5763
rect 5721 5723 5779 5729
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8352 5732 8401 5760
rect 8352 5720 8358 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 10060 5760 10088 5856
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 8389 5723 8447 5729
rect 9968 5732 10149 5760
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 9493 5695 9551 5701
rect 9493 5692 9505 5695
rect 3108 5664 9505 5692
rect 3108 5652 3114 5664
rect 9493 5661 9505 5664
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 9968 5636 9996 5732
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10318 5720 10324 5772
rect 10376 5760 10382 5772
rect 10686 5760 10692 5772
rect 10376 5732 10692 5760
rect 10376 5720 10382 5732
rect 10686 5720 10692 5732
rect 10744 5760 10750 5772
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10744 5732 10793 5760
rect 10744 5720 10750 5732
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 12066 5760 12072 5772
rect 11931 5732 12072 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 13188 5769 13216 5868
rect 13354 5856 13360 5868
rect 13412 5896 13418 5908
rect 20346 5896 20352 5908
rect 13412 5868 20352 5896
rect 13412 5856 13418 5868
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 35986 5856 35992 5908
rect 36044 5896 36050 5908
rect 42058 5896 42064 5908
rect 36044 5868 42064 5896
rect 36044 5856 36050 5868
rect 42058 5856 42064 5868
rect 42116 5856 42122 5908
rect 42702 5856 42708 5908
rect 42760 5896 42766 5908
rect 42760 5868 44312 5896
rect 42760 5856 42766 5868
rect 15286 5828 15292 5840
rect 14936 5800 15292 5828
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 13173 5763 13231 5769
rect 12575 5732 12609 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 13173 5729 13185 5763
rect 13219 5729 13231 5763
rect 13173 5723 13231 5729
rect 12544 5692 12572 5723
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 14936 5769 14964 5800
rect 15286 5788 15292 5800
rect 15344 5788 15350 5840
rect 38378 5788 38384 5840
rect 38436 5828 38442 5840
rect 38473 5831 38531 5837
rect 38473 5828 38485 5831
rect 38436 5800 38485 5828
rect 38436 5788 38442 5800
rect 38473 5797 38485 5800
rect 38519 5797 38531 5831
rect 38473 5791 38531 5797
rect 43806 5788 43812 5840
rect 43864 5828 43870 5840
rect 44082 5828 44088 5840
rect 43864 5800 44088 5828
rect 43864 5788 43870 5800
rect 44082 5788 44088 5800
rect 44140 5788 44146 5840
rect 44284 5828 44312 5868
rect 44450 5856 44456 5908
rect 44508 5896 44514 5908
rect 46106 5896 46112 5908
rect 44508 5868 46112 5896
rect 44508 5856 44514 5868
rect 46106 5856 46112 5868
rect 46164 5896 46170 5908
rect 46164 5868 47256 5896
rect 46164 5856 46170 5868
rect 46934 5828 46940 5840
rect 44284 5800 46940 5828
rect 13817 5763 13875 5769
rect 13817 5760 13829 5763
rect 13780 5732 13829 5760
rect 13780 5720 13786 5732
rect 13817 5729 13829 5732
rect 13863 5729 13875 5763
rect 13817 5723 13875 5729
rect 14921 5763 14979 5769
rect 14921 5729 14933 5763
rect 14967 5729 14979 5763
rect 15378 5760 15384 5772
rect 15339 5732 15384 5760
rect 14921 5723 14979 5729
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 15470 5692 15476 5704
rect 12406 5664 15476 5692
rect 7377 5627 7435 5633
rect 7377 5593 7389 5627
rect 7423 5624 7435 5627
rect 7423 5596 9904 5624
rect 7423 5593 7435 5596
rect 7377 5587 7435 5593
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 2372 5528 3893 5556
rect 2372 5516 2378 5528
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 6270 5556 6276 5568
rect 6231 5528 6276 5556
rect 3881 5519 3939 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 7742 5556 7748 5568
rect 6871 5528 7748 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 7929 5559 7987 5565
rect 7929 5525 7941 5559
rect 7975 5556 7987 5559
rect 9398 5556 9404 5568
rect 7975 5528 9404 5556
rect 7975 5525 7987 5528
rect 7929 5519 7987 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 9876 5556 9904 5596
rect 9950 5584 9956 5636
rect 10008 5584 10014 5636
rect 12406 5556 12434 5664
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 16316 5692 16344 5723
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16540 5732 16957 5760
rect 16540 5720 16546 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 16574 5692 16580 5704
rect 16316 5664 16580 5692
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16960 5692 16988 5723
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 17092 5732 17601 5760
rect 17092 5720 17098 5732
rect 17589 5729 17601 5732
rect 17635 5760 17647 5763
rect 20070 5760 20076 5772
rect 17635 5732 20076 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 33962 5720 33968 5772
rect 34020 5760 34026 5772
rect 39853 5763 39911 5769
rect 39853 5760 39865 5763
rect 34020 5732 39865 5760
rect 34020 5720 34026 5732
rect 39853 5729 39865 5732
rect 39899 5760 39911 5763
rect 40310 5760 40316 5772
rect 39899 5732 40316 5760
rect 39899 5729 39911 5732
rect 39853 5723 39911 5729
rect 40310 5720 40316 5732
rect 40368 5720 40374 5772
rect 41049 5763 41107 5769
rect 41049 5729 41061 5763
rect 41095 5760 41107 5763
rect 41322 5760 41328 5772
rect 41095 5732 41328 5760
rect 41095 5729 41107 5732
rect 41049 5723 41107 5729
rect 41322 5720 41328 5732
rect 41380 5720 41386 5772
rect 41693 5763 41751 5769
rect 41693 5729 41705 5763
rect 41739 5760 41751 5763
rect 41782 5760 41788 5772
rect 41739 5732 41788 5760
rect 41739 5729 41751 5732
rect 41693 5723 41751 5729
rect 41782 5720 41788 5732
rect 41840 5720 41846 5772
rect 42334 5760 42340 5772
rect 42295 5732 42340 5760
rect 42334 5720 42340 5732
rect 42392 5720 42398 5772
rect 42794 5760 42800 5772
rect 42755 5732 42800 5760
rect 42794 5720 42800 5732
rect 42852 5720 42858 5772
rect 43625 5763 43683 5769
rect 43625 5729 43637 5763
rect 43671 5760 43683 5763
rect 43990 5760 43996 5772
rect 43671 5732 43996 5760
rect 43671 5729 43683 5732
rect 43625 5723 43683 5729
rect 19334 5692 19340 5704
rect 16960 5664 19340 5692
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 37918 5652 37924 5704
rect 37976 5692 37982 5704
rect 43640 5692 43668 5723
rect 43990 5720 43996 5732
rect 44048 5720 44054 5772
rect 44284 5769 44312 5800
rect 46934 5788 46940 5800
rect 46992 5788 46998 5840
rect 44269 5763 44327 5769
rect 44269 5729 44281 5763
rect 44315 5729 44327 5763
rect 44913 5763 44971 5769
rect 44913 5760 44925 5763
rect 44269 5723 44327 5729
rect 44376 5732 44925 5760
rect 37976 5664 43668 5692
rect 37976 5652 37982 5664
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 19610 5624 19616 5636
rect 14516 5596 19616 5624
rect 14516 5584 14522 5596
rect 19610 5584 19616 5596
rect 19668 5584 19674 5636
rect 31938 5624 31944 5636
rect 31899 5596 31944 5624
rect 31938 5584 31944 5596
rect 31996 5584 32002 5636
rect 36814 5584 36820 5636
rect 36872 5624 36878 5636
rect 38289 5627 38347 5633
rect 38289 5624 38301 5627
rect 36872 5596 38301 5624
rect 36872 5584 36878 5596
rect 38289 5593 38301 5596
rect 38335 5593 38347 5627
rect 39206 5624 39212 5636
rect 39167 5596 39212 5624
rect 38289 5587 38347 5593
rect 39206 5584 39212 5596
rect 39264 5584 39270 5636
rect 40310 5584 40316 5636
rect 40368 5624 40374 5636
rect 40770 5624 40776 5636
rect 40368 5596 40776 5624
rect 40368 5584 40374 5596
rect 40770 5584 40776 5596
rect 40828 5584 40834 5636
rect 42150 5624 42156 5636
rect 41616 5596 42156 5624
rect 9876 5528 12434 5556
rect 18049 5559 18107 5565
rect 18049 5525 18061 5559
rect 18095 5556 18107 5559
rect 18138 5556 18144 5568
rect 18095 5528 18144 5556
rect 18095 5525 18107 5528
rect 18049 5519 18107 5525
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 24486 5556 24492 5568
rect 24447 5528 24492 5556
rect 24486 5516 24492 5528
rect 24544 5516 24550 5568
rect 24946 5516 24952 5568
rect 25004 5556 25010 5568
rect 25225 5559 25283 5565
rect 25225 5556 25237 5559
rect 25004 5528 25237 5556
rect 25004 5516 25010 5528
rect 25225 5525 25237 5528
rect 25271 5525 25283 5559
rect 25225 5519 25283 5525
rect 31754 5516 31760 5568
rect 31812 5556 31818 5568
rect 32030 5556 32036 5568
rect 31812 5528 31857 5556
rect 31991 5528 32036 5556
rect 31812 5516 31818 5528
rect 32030 5516 32036 5528
rect 32088 5516 32094 5568
rect 32306 5556 32312 5568
rect 32267 5528 32312 5556
rect 32306 5516 32312 5528
rect 32364 5516 32370 5568
rect 32490 5556 32496 5568
rect 32451 5528 32496 5556
rect 32490 5516 32496 5528
rect 32548 5516 32554 5568
rect 37734 5516 37740 5568
rect 37792 5556 37798 5568
rect 38562 5556 38568 5568
rect 37792 5528 38568 5556
rect 37792 5516 37798 5528
rect 38562 5516 38568 5528
rect 38620 5516 38626 5568
rect 39850 5516 39856 5568
rect 39908 5556 39914 5568
rect 41616 5556 41644 5596
rect 42150 5584 42156 5596
rect 42208 5584 42214 5636
rect 42794 5584 42800 5636
rect 42852 5624 42858 5636
rect 44376 5624 44404 5732
rect 44913 5729 44925 5732
rect 44959 5760 44971 5763
rect 45370 5760 45376 5772
rect 44959 5732 45376 5760
rect 44959 5729 44971 5732
rect 44913 5723 44971 5729
rect 45370 5720 45376 5732
rect 45428 5720 45434 5772
rect 46658 5720 46664 5772
rect 46716 5760 46722 5772
rect 47228 5769 47256 5868
rect 47670 5856 47676 5908
rect 47728 5896 47734 5908
rect 47854 5896 47860 5908
rect 47728 5868 47860 5896
rect 47728 5856 47734 5868
rect 47854 5856 47860 5868
rect 47912 5856 47918 5908
rect 66530 5788 66536 5840
rect 66588 5828 66594 5840
rect 67177 5831 67235 5837
rect 67177 5828 67189 5831
rect 66588 5800 67189 5828
rect 66588 5788 66594 5800
rect 67177 5797 67189 5800
rect 67223 5797 67235 5831
rect 67177 5791 67235 5797
rect 67818 5788 67824 5840
rect 67876 5828 67882 5840
rect 67913 5831 67971 5837
rect 67913 5828 67925 5831
rect 67876 5800 67925 5828
rect 67876 5788 67882 5800
rect 67913 5797 67925 5800
rect 67959 5797 67971 5831
rect 67913 5791 67971 5797
rect 46753 5763 46811 5769
rect 46753 5760 46765 5763
rect 46716 5732 46765 5760
rect 46716 5720 46722 5732
rect 46753 5729 46765 5732
rect 46799 5729 46811 5763
rect 46753 5723 46811 5729
rect 47213 5763 47271 5769
rect 47213 5729 47225 5763
rect 47259 5729 47271 5763
rect 47213 5723 47271 5729
rect 48041 5763 48099 5769
rect 48041 5729 48053 5763
rect 48087 5760 48099 5763
rect 48130 5760 48136 5772
rect 48087 5732 48136 5760
rect 48087 5729 48099 5732
rect 48041 5723 48099 5729
rect 48056 5692 48084 5723
rect 48130 5720 48136 5732
rect 48188 5720 48194 5772
rect 48498 5720 48504 5772
rect 48556 5760 48562 5772
rect 48685 5763 48743 5769
rect 48685 5760 48697 5763
rect 48556 5732 48697 5760
rect 48556 5720 48562 5732
rect 48685 5729 48697 5732
rect 48731 5729 48743 5763
rect 48685 5723 48743 5729
rect 49050 5720 49056 5772
rect 49108 5760 49114 5772
rect 49329 5763 49387 5769
rect 49329 5760 49341 5763
rect 49108 5732 49341 5760
rect 49108 5720 49114 5732
rect 49329 5729 49341 5732
rect 49375 5729 49387 5763
rect 49329 5723 49387 5729
rect 49973 5763 50031 5769
rect 49973 5729 49985 5763
rect 50019 5760 50031 5763
rect 50154 5760 50160 5772
rect 50019 5732 50160 5760
rect 50019 5729 50031 5732
rect 49973 5723 50031 5729
rect 50154 5720 50160 5732
rect 50212 5720 50218 5772
rect 51166 5720 51172 5772
rect 51224 5760 51230 5772
rect 51445 5763 51503 5769
rect 51445 5760 51457 5763
rect 51224 5732 51457 5760
rect 51224 5720 51230 5732
rect 51445 5729 51457 5732
rect 51491 5760 51503 5763
rect 51718 5760 51724 5772
rect 51491 5732 51724 5760
rect 51491 5729 51503 5732
rect 51445 5723 51503 5729
rect 51718 5720 51724 5732
rect 51776 5720 51782 5772
rect 52089 5763 52147 5769
rect 52089 5729 52101 5763
rect 52135 5760 52147 5763
rect 52362 5760 52368 5772
rect 52135 5732 52368 5760
rect 52135 5729 52147 5732
rect 52089 5723 52147 5729
rect 52104 5692 52132 5723
rect 52362 5720 52368 5732
rect 52420 5720 52426 5772
rect 52733 5763 52791 5769
rect 52733 5729 52745 5763
rect 52779 5729 52791 5763
rect 52733 5723 52791 5729
rect 45388 5664 48084 5692
rect 51736 5664 52132 5692
rect 52748 5692 52776 5723
rect 52822 5720 52828 5772
rect 52880 5760 52886 5772
rect 53193 5763 53251 5769
rect 53193 5760 53205 5763
rect 52880 5732 53205 5760
rect 52880 5720 52886 5732
rect 53193 5729 53205 5732
rect 53239 5729 53251 5763
rect 53193 5723 53251 5729
rect 54021 5763 54079 5769
rect 54021 5729 54033 5763
rect 54067 5729 54079 5763
rect 54021 5723 54079 5729
rect 54665 5763 54723 5769
rect 54665 5729 54677 5763
rect 54711 5760 54723 5763
rect 55030 5760 55036 5772
rect 54711 5732 55036 5760
rect 54711 5729 54723 5732
rect 54665 5723 54723 5729
rect 52914 5692 52920 5704
rect 52748 5664 52920 5692
rect 45388 5636 45416 5664
rect 51736 5636 51764 5664
rect 52914 5652 52920 5664
rect 52972 5652 52978 5704
rect 53098 5652 53104 5704
rect 53156 5692 53162 5704
rect 54036 5692 54064 5723
rect 55030 5720 55036 5732
rect 55088 5720 55094 5772
rect 55309 5763 55367 5769
rect 55309 5729 55321 5763
rect 55355 5760 55367 5763
rect 55490 5760 55496 5772
rect 55355 5732 55496 5760
rect 55355 5729 55367 5732
rect 55309 5723 55367 5729
rect 55490 5720 55496 5732
rect 55548 5720 55554 5772
rect 56410 5720 56416 5772
rect 56468 5760 56474 5772
rect 56689 5763 56747 5769
rect 56689 5760 56701 5763
rect 56468 5732 56701 5760
rect 56468 5720 56474 5732
rect 56689 5729 56701 5732
rect 56735 5729 56747 5763
rect 56689 5723 56747 5729
rect 62574 5720 62580 5772
rect 62632 5760 62638 5772
rect 62853 5763 62911 5769
rect 62853 5760 62865 5763
rect 62632 5732 62865 5760
rect 62632 5720 62638 5732
rect 62853 5729 62865 5732
rect 62899 5729 62911 5763
rect 63494 5760 63500 5772
rect 63455 5732 63500 5760
rect 62853 5723 62911 5729
rect 63494 5720 63500 5732
rect 63552 5720 63558 5772
rect 64046 5720 64052 5772
rect 64104 5760 64110 5772
rect 64325 5763 64383 5769
rect 64325 5760 64337 5763
rect 64104 5732 64337 5760
rect 64104 5720 64110 5732
rect 64325 5729 64337 5732
rect 64371 5760 64383 5763
rect 64598 5760 64604 5772
rect 64371 5732 64604 5760
rect 64371 5729 64383 5732
rect 64325 5723 64383 5729
rect 64598 5720 64604 5732
rect 64656 5720 64662 5772
rect 65429 5763 65487 5769
rect 65429 5729 65441 5763
rect 65475 5729 65487 5763
rect 65429 5723 65487 5729
rect 66073 5763 66131 5769
rect 66073 5729 66085 5763
rect 66119 5760 66131 5763
rect 66162 5760 66168 5772
rect 66119 5732 66168 5760
rect 66119 5729 66131 5732
rect 66073 5723 66131 5729
rect 54938 5692 54944 5704
rect 53156 5664 54944 5692
rect 53156 5652 53162 5664
rect 54938 5652 54944 5664
rect 54996 5652 55002 5704
rect 65444 5692 65472 5723
rect 66162 5720 66168 5732
rect 66220 5720 66226 5772
rect 68094 5760 68100 5772
rect 68055 5732 68100 5760
rect 68094 5720 68100 5732
rect 68152 5720 68158 5772
rect 65610 5692 65616 5704
rect 65444 5664 65616 5692
rect 65610 5652 65616 5664
rect 65668 5692 65674 5704
rect 69014 5692 69020 5704
rect 65668 5664 69020 5692
rect 65668 5652 65674 5664
rect 69014 5652 69020 5664
rect 69072 5652 69078 5704
rect 42852 5596 44404 5624
rect 42852 5584 42858 5596
rect 44450 5584 44456 5636
rect 44508 5584 44514 5636
rect 45370 5584 45376 5636
rect 45428 5584 45434 5636
rect 51718 5584 51724 5636
rect 51776 5584 51782 5636
rect 51994 5584 52000 5636
rect 52052 5624 52058 5636
rect 52362 5624 52368 5636
rect 52052 5596 52368 5624
rect 52052 5584 52058 5596
rect 52362 5584 52368 5596
rect 52420 5584 52426 5636
rect 60550 5584 60556 5636
rect 60608 5624 60614 5636
rect 60737 5627 60795 5633
rect 60737 5624 60749 5627
rect 60608 5596 60749 5624
rect 60608 5584 60614 5596
rect 60737 5593 60749 5596
rect 60783 5593 60795 5627
rect 60737 5587 60795 5593
rect 64506 5584 64512 5636
rect 64564 5584 64570 5636
rect 67361 5627 67419 5633
rect 67361 5593 67373 5627
rect 67407 5624 67419 5627
rect 69842 5624 69848 5636
rect 67407 5596 69848 5624
rect 67407 5593 67419 5596
rect 67361 5587 67419 5593
rect 69842 5584 69848 5596
rect 69900 5584 69906 5636
rect 39908 5528 41644 5556
rect 39908 5516 39914 5528
rect 41690 5516 41696 5568
rect 41748 5556 41754 5568
rect 44468 5556 44496 5584
rect 41748 5528 44496 5556
rect 41748 5516 41754 5528
rect 44542 5516 44548 5568
rect 44600 5556 44606 5568
rect 45649 5559 45707 5565
rect 45649 5556 45661 5559
rect 44600 5528 45661 5556
rect 44600 5516 44606 5528
rect 45649 5525 45661 5528
rect 45695 5525 45707 5559
rect 45649 5519 45707 5525
rect 56778 5516 56784 5568
rect 56836 5556 56842 5568
rect 57149 5559 57207 5565
rect 57149 5556 57161 5559
rect 56836 5528 57161 5556
rect 56836 5516 56842 5528
rect 57149 5525 57161 5528
rect 57195 5525 57207 5559
rect 57698 5556 57704 5568
rect 57659 5528 57704 5556
rect 57149 5519 57207 5525
rect 57698 5516 57704 5528
rect 57756 5516 57762 5568
rect 58802 5556 58808 5568
rect 58763 5528 58808 5556
rect 58802 5516 58808 5528
rect 58860 5516 58866 5568
rect 59357 5559 59415 5565
rect 59357 5525 59369 5559
rect 59403 5556 59415 5559
rect 59998 5556 60004 5568
rect 59403 5528 60004 5556
rect 59403 5525 59415 5528
rect 59357 5519 59415 5525
rect 59998 5516 60004 5528
rect 60056 5516 60062 5568
rect 60274 5556 60280 5568
rect 60235 5528 60280 5556
rect 60274 5516 60280 5528
rect 60332 5516 60338 5568
rect 60458 5516 60464 5568
rect 60516 5556 60522 5568
rect 61381 5559 61439 5565
rect 61381 5556 61393 5559
rect 60516 5528 61393 5556
rect 60516 5516 60522 5528
rect 61381 5525 61393 5528
rect 61427 5525 61439 5559
rect 61381 5519 61439 5525
rect 61746 5516 61752 5568
rect 61804 5556 61810 5568
rect 61933 5559 61991 5565
rect 61933 5556 61945 5559
rect 61804 5528 61945 5556
rect 61804 5516 61810 5528
rect 61933 5525 61945 5528
rect 61979 5525 61991 5559
rect 64524 5556 64552 5584
rect 64690 5556 64696 5568
rect 64524 5528 64696 5556
rect 61933 5519 61991 5525
rect 64690 5516 64696 5528
rect 64748 5516 64754 5568
rect 37274 5488 37280 5500
rect 1104 5466 18952 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 14246 5466
rect 14298 5414 14310 5466
rect 14362 5414 14374 5466
rect 14426 5414 14438 5466
rect 14490 5414 18952 5466
rect 1104 5392 18952 5414
rect 31726 5460 37280 5488
rect 12158 5312 12164 5364
rect 12216 5352 12222 5364
rect 31726 5352 31754 5460
rect 37274 5448 37280 5460
rect 37332 5448 37338 5500
rect 37628 5466 68816 5488
rect 37628 5414 44246 5466
rect 44298 5414 44310 5466
rect 44362 5414 44374 5466
rect 44426 5414 44438 5466
rect 44490 5414 54246 5466
rect 54298 5414 54310 5466
rect 54362 5414 54374 5466
rect 54426 5414 54438 5466
rect 54490 5414 64246 5466
rect 64298 5414 64310 5466
rect 64362 5414 64374 5466
rect 64426 5414 64438 5466
rect 64490 5414 68816 5466
rect 37628 5392 68816 5414
rect 12216 5324 31754 5352
rect 12216 5312 12222 5324
rect 36170 5312 36176 5364
rect 36228 5352 36234 5364
rect 39853 5355 39911 5361
rect 39853 5352 39865 5355
rect 36228 5324 39865 5352
rect 36228 5312 36234 5324
rect 39853 5321 39865 5324
rect 39899 5321 39911 5355
rect 39853 5315 39911 5321
rect 40218 5312 40224 5364
rect 40276 5352 40282 5364
rect 46198 5352 46204 5364
rect 40276 5324 46204 5352
rect 40276 5312 40282 5324
rect 46198 5312 46204 5324
rect 46256 5312 46262 5364
rect 48314 5352 48320 5364
rect 48148 5324 48320 5352
rect 4798 5244 4804 5296
rect 4856 5244 4862 5296
rect 5442 5284 5448 5296
rect 4908 5256 5448 5284
rect 4062 5216 4068 5228
rect 2884 5188 4068 5216
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1486 5148 1492 5160
rect 1443 5120 1492 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1486 5108 1492 5120
rect 1544 5108 1550 5160
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 1946 5148 1952 5160
rect 1636 5120 1952 5148
rect 1636 5108 1642 5120
rect 1946 5108 1952 5120
rect 2004 5148 2010 5160
rect 2041 5151 2099 5157
rect 2041 5148 2053 5151
rect 2004 5120 2053 5148
rect 2004 5108 2010 5120
rect 2041 5117 2053 5120
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 2884 5157 2912 5188
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4816 5216 4844 5244
rect 4172 5188 4844 5216
rect 4172 5160 4200 5188
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 2832 5120 2881 5148
rect 2832 5108 2838 5120
rect 2869 5117 2881 5120
rect 2915 5117 2927 5151
rect 2869 5111 2927 5117
rect 3326 5108 3332 5160
rect 3384 5148 3390 5160
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 3384 5120 3525 5148
rect 3384 5108 3390 5120
rect 3513 5117 3525 5120
rect 3559 5148 3571 5151
rect 3878 5148 3884 5160
rect 3559 5120 3884 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 4154 5148 4160 5160
rect 4067 5120 4160 5148
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4798 5148 4804 5160
rect 4711 5120 4804 5148
rect 4798 5108 4804 5120
rect 4856 5148 4862 5160
rect 4908 5148 4936 5256
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 9030 5244 9036 5296
rect 9088 5244 9094 5296
rect 9398 5244 9404 5296
rect 9456 5284 9462 5296
rect 20714 5284 20720 5296
rect 9456 5256 20720 5284
rect 9456 5244 9462 5256
rect 9048 5216 9076 5244
rect 9048 5188 9536 5216
rect 5442 5148 5448 5160
rect 4856 5120 4936 5148
rect 5403 5120 5448 5148
rect 4856 5108 4862 5120
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 6638 5148 6644 5160
rect 6144 5120 6644 5148
rect 6144 5108 6150 5120
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6696 5120 6837 5148
rect 6696 5108 6702 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 7558 5148 7564 5160
rect 7340 5120 7564 5148
rect 7340 5108 7346 5120
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 8110 5148 8116 5160
rect 7668 5120 8116 5148
rect 7466 5040 7472 5092
rect 7524 5080 7530 5092
rect 7668 5080 7696 5120
rect 8110 5108 8116 5120
rect 8168 5148 8174 5160
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 8168 5120 8217 5148
rect 8168 5108 8174 5120
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 8846 5108 8852 5160
rect 8904 5148 8910 5160
rect 9508 5157 9536 5188
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8904 5120 9045 5148
rect 8904 5108 8910 5120
rect 9033 5117 9045 5120
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5117 9551 5151
rect 9493 5111 9551 5117
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 9858 5148 9864 5160
rect 9732 5120 9864 5148
rect 9732 5108 9738 5120
rect 9858 5108 9864 5120
rect 9916 5148 9922 5160
rect 12728 5157 12756 5256
rect 20714 5244 20720 5256
rect 20772 5244 20778 5296
rect 23566 5244 23572 5296
rect 23624 5284 23630 5296
rect 42334 5284 42340 5296
rect 23624 5256 42340 5284
rect 23624 5244 23630 5256
rect 42334 5244 42340 5256
rect 42392 5284 42398 5296
rect 42610 5284 42616 5296
rect 42392 5256 42616 5284
rect 42392 5244 42398 5256
rect 42610 5244 42616 5256
rect 42668 5244 42674 5296
rect 44174 5244 44180 5296
rect 44232 5284 44238 5296
rect 45094 5284 45100 5296
rect 44232 5256 45100 5284
rect 44232 5244 44238 5256
rect 14550 5216 14556 5228
rect 14016 5188 14556 5216
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 9916 5120 10149 5148
rect 9916 5108 9922 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5117 12771 5151
rect 13354 5148 13360 5160
rect 13315 5120 13360 5148
rect 12713 5111 12771 5117
rect 7524 5052 7696 5080
rect 7524 5040 7530 5052
rect 7742 5040 7748 5092
rect 7800 5080 7806 5092
rect 11164 5080 11192 5111
rect 13354 5108 13360 5120
rect 13412 5148 13418 5160
rect 13538 5148 13544 5160
rect 13412 5120 13544 5148
rect 13412 5108 13418 5120
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 14016 5157 14044 5188
rect 14550 5176 14556 5188
rect 14608 5216 14614 5228
rect 14918 5216 14924 5228
rect 14608 5188 14924 5216
rect 14608 5176 14614 5188
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 21818 5216 21824 5228
rect 15028 5188 21824 5216
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5117 14059 5151
rect 15028 5148 15056 5188
rect 14001 5111 14059 5117
rect 14292 5120 15056 5148
rect 15381 5151 15439 5157
rect 7800 5052 11192 5080
rect 7800 5040 7806 5052
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10962 5012 10968 5024
rect 9916 4984 10968 5012
rect 9916 4972 9922 4984
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11164 5012 11192 5052
rect 12069 5083 12127 5089
rect 12069 5049 12081 5083
rect 12115 5080 12127 5083
rect 14292 5080 14320 5120
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 15562 5148 15568 5160
rect 15427 5120 15568 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 16408 5157 16436 5188
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 32953 5219 33011 5225
rect 32953 5185 32965 5219
rect 32999 5216 33011 5219
rect 33042 5216 33048 5228
rect 32999 5188 33048 5216
rect 32999 5185 33011 5188
rect 32953 5179 33011 5185
rect 33042 5176 33048 5188
rect 33100 5176 33106 5228
rect 34977 5219 35035 5225
rect 34977 5185 34989 5219
rect 35023 5216 35035 5219
rect 44542 5216 44548 5228
rect 35023 5188 44548 5216
rect 35023 5185 35035 5188
rect 34977 5179 35035 5185
rect 16393 5151 16451 5157
rect 16393 5117 16405 5151
rect 16439 5117 16451 5151
rect 17862 5148 17868 5160
rect 17823 5120 17868 5148
rect 16393 5111 16451 5117
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 37734 5108 37740 5160
rect 37792 5148 37798 5160
rect 37792 5120 38608 5148
rect 37792 5108 37798 5120
rect 12115 5052 14320 5080
rect 12115 5049 12127 5052
rect 12069 5043 12127 5049
rect 14458 5040 14464 5092
rect 14516 5080 14522 5092
rect 14516 5052 14561 5080
rect 14516 5040 14522 5052
rect 14642 5040 14648 5092
rect 14700 5080 14706 5092
rect 15580 5080 15608 5108
rect 16945 5083 17003 5089
rect 16945 5080 16957 5083
rect 14700 5052 14745 5080
rect 15580 5052 16957 5080
rect 14700 5040 14706 5052
rect 16945 5049 16957 5052
rect 16991 5049 17003 5083
rect 17678 5080 17684 5092
rect 17639 5052 17684 5080
rect 16945 5043 17003 5049
rect 17678 5040 17684 5052
rect 17736 5040 17742 5092
rect 33413 5083 33471 5089
rect 33413 5049 33425 5083
rect 33459 5080 33471 5083
rect 38289 5083 38347 5089
rect 38289 5080 38301 5083
rect 33459 5052 38301 5080
rect 33459 5049 33471 5052
rect 33413 5043 33471 5049
rect 38289 5049 38301 5052
rect 38335 5049 38347 5083
rect 38289 5043 38347 5049
rect 38378 5040 38384 5092
rect 38436 5080 38442 5092
rect 38473 5083 38531 5089
rect 38473 5080 38485 5083
rect 38436 5052 38485 5080
rect 38436 5040 38442 5052
rect 38473 5049 38485 5052
rect 38519 5049 38531 5083
rect 38580 5080 38608 5120
rect 38838 5108 38844 5160
rect 38896 5148 38902 5160
rect 39209 5151 39267 5157
rect 39209 5148 39221 5151
rect 38896 5120 39221 5148
rect 38896 5108 38902 5120
rect 39209 5117 39221 5120
rect 39255 5117 39267 5151
rect 39209 5111 39267 5117
rect 39758 5108 39764 5160
rect 39816 5148 39822 5160
rect 41233 5151 41291 5157
rect 41233 5148 41245 5151
rect 39816 5120 41245 5148
rect 39816 5108 39822 5120
rect 41233 5117 41245 5120
rect 41279 5117 41291 5151
rect 41233 5111 41291 5117
rect 41417 5151 41475 5157
rect 41417 5117 41429 5151
rect 41463 5148 41475 5151
rect 41966 5148 41972 5160
rect 41463 5120 41972 5148
rect 41463 5117 41475 5120
rect 41417 5111 41475 5117
rect 41966 5108 41972 5120
rect 42024 5108 42030 5160
rect 42168 5157 42196 5188
rect 44542 5176 44548 5188
rect 44600 5176 44606 5228
rect 42153 5151 42211 5157
rect 42153 5117 42165 5151
rect 42199 5117 42211 5151
rect 42153 5111 42211 5117
rect 43346 5108 43352 5160
rect 43404 5148 43410 5160
rect 43533 5151 43591 5157
rect 43533 5148 43545 5151
rect 43404 5120 43545 5148
rect 43404 5108 43410 5120
rect 43533 5117 43545 5120
rect 43579 5148 43591 5151
rect 44177 5151 44235 5157
rect 43579 5120 44128 5148
rect 43579 5117 43591 5120
rect 43533 5111 43591 5117
rect 39945 5083 40003 5089
rect 38580 5052 39252 5080
rect 38473 5043 38531 5049
rect 17494 5012 17500 5024
rect 11164 4984 17500 5012
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 37182 4972 37188 5024
rect 37240 5012 37246 5024
rect 39117 5015 39175 5021
rect 39117 5012 39129 5015
rect 37240 4984 39129 5012
rect 37240 4972 37246 4984
rect 39117 4981 39129 4984
rect 39163 4981 39175 5015
rect 39224 5012 39252 5052
rect 39945 5049 39957 5083
rect 39991 5080 40003 5083
rect 40218 5080 40224 5092
rect 39991 5052 40224 5080
rect 39991 5049 40003 5052
rect 39945 5043 40003 5049
rect 40218 5040 40224 5052
rect 40276 5040 40282 5092
rect 40681 5083 40739 5089
rect 40681 5049 40693 5083
rect 40727 5080 40739 5083
rect 42518 5080 42524 5092
rect 40727 5052 42524 5080
rect 40727 5049 40739 5052
rect 40681 5043 40739 5049
rect 42518 5040 42524 5052
rect 42576 5040 42582 5092
rect 42610 5040 42616 5092
rect 42668 5080 42674 5092
rect 44100 5080 44128 5120
rect 44177 5117 44189 5151
rect 44223 5148 44235 5151
rect 44450 5148 44456 5160
rect 44223 5120 44456 5148
rect 44223 5117 44235 5120
rect 44177 5111 44235 5117
rect 44450 5108 44456 5120
rect 44508 5108 44514 5160
rect 44652 5157 44680 5256
rect 45094 5244 45100 5256
rect 45152 5244 45158 5296
rect 47946 5216 47952 5228
rect 46124 5188 47952 5216
rect 44637 5151 44695 5157
rect 44637 5117 44649 5151
rect 44683 5117 44695 5151
rect 44637 5111 44695 5117
rect 45465 5151 45523 5157
rect 45465 5117 45477 5151
rect 45511 5148 45523 5151
rect 45646 5148 45652 5160
rect 45511 5120 45652 5148
rect 45511 5117 45523 5120
rect 45465 5111 45523 5117
rect 45646 5108 45652 5120
rect 45704 5108 45710 5160
rect 45830 5108 45836 5160
rect 45888 5148 45894 5160
rect 46124 5157 46152 5188
rect 47946 5176 47952 5188
rect 48004 5176 48010 5228
rect 46109 5151 46167 5157
rect 46109 5148 46121 5151
rect 45888 5120 46121 5148
rect 45888 5108 45894 5120
rect 46109 5117 46121 5120
rect 46155 5117 46167 5151
rect 46750 5148 46756 5160
rect 46711 5120 46756 5148
rect 46109 5111 46167 5117
rect 46750 5108 46756 5120
rect 46808 5108 46814 5160
rect 47302 5108 47308 5160
rect 47360 5148 47366 5160
rect 47397 5151 47455 5157
rect 47397 5148 47409 5151
rect 47360 5120 47409 5148
rect 47360 5108 47366 5120
rect 47397 5117 47409 5120
rect 47443 5117 47455 5151
rect 47397 5111 47455 5117
rect 46382 5080 46388 5092
rect 42668 5052 43760 5080
rect 44100 5052 46388 5080
rect 42668 5040 42674 5052
rect 40589 5015 40647 5021
rect 40589 5012 40601 5015
rect 39224 4984 40601 5012
rect 39117 4975 39175 4981
rect 40589 4981 40601 4984
rect 40635 4981 40647 5015
rect 43732 5012 43760 5052
rect 46382 5040 46388 5052
rect 46440 5040 46446 5092
rect 48148 5024 48176 5324
rect 48314 5312 48320 5324
rect 48372 5312 48378 5364
rect 50522 5244 50528 5296
rect 50580 5284 50586 5296
rect 51169 5287 51227 5293
rect 51169 5284 51181 5287
rect 50580 5256 51181 5284
rect 50580 5244 50586 5256
rect 51169 5253 51181 5256
rect 51215 5253 51227 5287
rect 51169 5247 51227 5253
rect 63586 5244 63592 5296
rect 63644 5284 63650 5296
rect 64230 5284 64236 5296
rect 63644 5256 64236 5284
rect 63644 5244 63650 5256
rect 64230 5244 64236 5256
rect 64288 5244 64294 5296
rect 48314 5176 48320 5228
rect 48372 5216 48378 5228
rect 49421 5219 49479 5225
rect 49421 5216 49433 5219
rect 48372 5188 49433 5216
rect 48372 5176 48378 5188
rect 49421 5185 49433 5188
rect 49467 5185 49479 5219
rect 49421 5179 49479 5185
rect 51074 5176 51080 5228
rect 51132 5216 51138 5228
rect 51132 5188 52132 5216
rect 51132 5176 51138 5188
rect 52104 5160 52132 5188
rect 60826 5176 60832 5228
rect 60884 5216 60890 5228
rect 60884 5188 67956 5216
rect 60884 5176 60890 5188
rect 48590 5108 48596 5160
rect 48648 5148 48654 5160
rect 48777 5151 48835 5157
rect 48777 5148 48789 5151
rect 48648 5120 48789 5148
rect 48648 5108 48654 5120
rect 48777 5117 48789 5120
rect 48823 5117 48835 5151
rect 48777 5111 48835 5117
rect 50065 5151 50123 5157
rect 50065 5117 50077 5151
rect 50111 5148 50123 5151
rect 50338 5148 50344 5160
rect 50111 5120 50344 5148
rect 50111 5117 50123 5120
rect 50065 5111 50123 5117
rect 50338 5108 50344 5120
rect 50396 5148 50402 5160
rect 50522 5148 50528 5160
rect 50396 5120 50528 5148
rect 50396 5108 50402 5120
rect 50522 5108 50528 5120
rect 50580 5108 50586 5160
rect 50614 5108 50620 5160
rect 50672 5148 50678 5160
rect 51721 5151 51779 5157
rect 50672 5120 51488 5148
rect 50672 5108 50678 5120
rect 51350 5080 51356 5092
rect 51311 5052 51356 5080
rect 51350 5040 51356 5052
rect 51408 5040 51414 5092
rect 48130 5012 48136 5024
rect 43732 4984 48136 5012
rect 40589 4975 40647 4981
rect 48130 4972 48136 4984
rect 48188 4972 48194 5024
rect 51460 5021 51488 5120
rect 51721 5117 51733 5151
rect 51767 5148 51779 5151
rect 51902 5148 51908 5160
rect 51767 5120 51908 5148
rect 51767 5117 51779 5120
rect 51721 5111 51779 5117
rect 51902 5108 51908 5120
rect 51960 5108 51966 5160
rect 52086 5108 52092 5160
rect 52144 5148 52150 5160
rect 52181 5151 52239 5157
rect 52181 5148 52193 5151
rect 52144 5120 52193 5148
rect 52144 5108 52150 5120
rect 52181 5117 52193 5120
rect 52227 5117 52239 5151
rect 52181 5111 52239 5117
rect 53742 5108 53748 5160
rect 53800 5148 53806 5160
rect 54021 5151 54079 5157
rect 54021 5148 54033 5151
rect 53800 5120 54033 5148
rect 53800 5108 53806 5120
rect 54021 5117 54033 5120
rect 54067 5117 54079 5151
rect 54021 5111 54079 5117
rect 54481 5151 54539 5157
rect 54481 5117 54493 5151
rect 54527 5117 54539 5151
rect 54481 5111 54539 5117
rect 53834 5040 53840 5092
rect 53892 5080 53898 5092
rect 54496 5080 54524 5111
rect 54938 5108 54944 5160
rect 54996 5148 55002 5160
rect 55309 5151 55367 5157
rect 55309 5148 55321 5151
rect 54996 5120 55321 5148
rect 54996 5108 55002 5120
rect 55309 5117 55321 5120
rect 55355 5148 55367 5151
rect 55398 5148 55404 5160
rect 55355 5120 55404 5148
rect 55355 5117 55367 5120
rect 55309 5111 55367 5117
rect 55398 5108 55404 5120
rect 55456 5108 55462 5160
rect 55950 5148 55956 5160
rect 55863 5120 55956 5148
rect 55950 5108 55956 5120
rect 56008 5148 56014 5160
rect 56318 5148 56324 5160
rect 56008 5120 56324 5148
rect 56008 5108 56014 5120
rect 56318 5108 56324 5120
rect 56376 5108 56382 5160
rect 56413 5151 56471 5157
rect 56413 5117 56425 5151
rect 56459 5117 56471 5151
rect 56413 5111 56471 5117
rect 53892 5052 54524 5080
rect 53892 5040 53898 5052
rect 55766 5040 55772 5092
rect 55824 5080 55830 5092
rect 56226 5080 56232 5092
rect 55824 5052 56232 5080
rect 55824 5040 55830 5052
rect 56226 5040 56232 5052
rect 56284 5080 56290 5092
rect 56428 5080 56456 5111
rect 56594 5108 56600 5160
rect 56652 5148 56658 5160
rect 57238 5148 57244 5160
rect 56652 5120 57244 5148
rect 56652 5108 56658 5120
rect 57238 5108 57244 5120
rect 57296 5108 57302 5160
rect 57606 5108 57612 5160
rect 57664 5148 57670 5160
rect 57885 5151 57943 5157
rect 57885 5148 57897 5151
rect 57664 5120 57897 5148
rect 57664 5108 57670 5120
rect 57885 5117 57897 5120
rect 57931 5117 57943 5151
rect 57885 5111 57943 5117
rect 59906 5108 59912 5160
rect 59964 5148 59970 5160
rect 60093 5151 60151 5157
rect 60093 5148 60105 5151
rect 59964 5120 60105 5148
rect 59964 5108 59970 5120
rect 60093 5117 60105 5120
rect 60139 5117 60151 5151
rect 60093 5111 60151 5117
rect 60366 5108 60372 5160
rect 60424 5148 60430 5160
rect 60553 5151 60611 5157
rect 60553 5148 60565 5151
rect 60424 5120 60565 5148
rect 60424 5108 60430 5120
rect 60553 5117 60565 5120
rect 60599 5117 60611 5151
rect 60553 5111 60611 5117
rect 60734 5108 60740 5160
rect 60792 5148 60798 5160
rect 61378 5148 61384 5160
rect 60792 5120 61384 5148
rect 60792 5108 60798 5120
rect 61378 5108 61384 5120
rect 61436 5108 61442 5160
rect 61841 5151 61899 5157
rect 61841 5117 61853 5151
rect 61887 5148 61899 5151
rect 62022 5148 62028 5160
rect 61887 5120 62028 5148
rect 61887 5117 61899 5120
rect 61841 5111 61899 5117
rect 56284 5052 56456 5080
rect 56284 5040 56290 5052
rect 61286 5040 61292 5092
rect 61344 5080 61350 5092
rect 61856 5080 61884 5111
rect 62022 5108 62028 5120
rect 62080 5108 62086 5160
rect 62114 5108 62120 5160
rect 62172 5148 62178 5160
rect 62669 5151 62727 5157
rect 62669 5148 62681 5151
rect 62172 5120 62681 5148
rect 62172 5108 62178 5120
rect 62669 5117 62681 5120
rect 62715 5148 62727 5151
rect 62758 5148 62764 5160
rect 62715 5120 62764 5148
rect 62715 5117 62727 5120
rect 62669 5111 62727 5117
rect 62758 5108 62764 5120
rect 62816 5108 62822 5160
rect 63034 5108 63040 5160
rect 63092 5148 63098 5160
rect 63129 5151 63187 5157
rect 63129 5148 63141 5151
rect 63092 5120 63141 5148
rect 63092 5108 63098 5120
rect 63129 5117 63141 5120
rect 63175 5117 63187 5151
rect 63129 5111 63187 5117
rect 63586 5108 63592 5160
rect 63644 5148 63650 5160
rect 63862 5148 63868 5160
rect 63644 5120 63868 5148
rect 63644 5108 63650 5120
rect 63862 5108 63868 5120
rect 63920 5148 63926 5160
rect 64325 5151 64383 5157
rect 64325 5148 64337 5151
rect 63920 5120 64337 5148
rect 63920 5108 63926 5120
rect 64325 5117 64337 5120
rect 64371 5117 64383 5151
rect 65150 5148 65156 5160
rect 65063 5120 65156 5148
rect 64325 5111 64383 5117
rect 65150 5108 65156 5120
rect 65208 5108 65214 5160
rect 65610 5108 65616 5160
rect 65668 5148 65674 5160
rect 65797 5151 65855 5157
rect 65797 5148 65809 5151
rect 65668 5120 65809 5148
rect 65668 5108 65674 5120
rect 65797 5117 65809 5120
rect 65843 5148 65855 5151
rect 65886 5148 65892 5160
rect 65843 5120 65892 5148
rect 65843 5117 65855 5120
rect 65797 5111 65855 5117
rect 65886 5108 65892 5120
rect 65944 5108 65950 5160
rect 66441 5151 66499 5157
rect 66441 5117 66453 5151
rect 66487 5148 66499 5151
rect 66622 5148 66628 5160
rect 66487 5120 66628 5148
rect 66487 5117 66499 5120
rect 66441 5111 66499 5117
rect 66622 5108 66628 5120
rect 66680 5108 66686 5160
rect 67928 5157 67956 5188
rect 67913 5151 67971 5157
rect 67913 5117 67925 5151
rect 67959 5117 67971 5151
rect 67913 5111 67971 5117
rect 61344 5052 61884 5080
rect 61344 5040 61350 5052
rect 51445 5015 51503 5021
rect 51445 4981 51457 5015
rect 51491 4981 51503 5015
rect 51445 4975 51503 4981
rect 51534 4972 51540 5024
rect 51592 5012 51598 5024
rect 51592 4984 51637 5012
rect 51592 4972 51598 4984
rect 51994 4972 52000 5024
rect 52052 5012 52058 5024
rect 52825 5015 52883 5021
rect 52825 5012 52837 5015
rect 52052 4984 52837 5012
rect 52052 4972 52058 4984
rect 52825 4981 52837 4984
rect 52871 4981 52883 5015
rect 58710 5012 58716 5024
rect 58671 4984 58716 5012
rect 52825 4975 52883 4981
rect 58710 4972 58716 4984
rect 58768 4972 58774 5024
rect 59357 5015 59415 5021
rect 59357 4981 59369 5015
rect 59403 5012 59415 5015
rect 59538 5012 59544 5024
rect 59403 4984 59544 5012
rect 59403 4981 59415 4984
rect 59357 4975 59415 4981
rect 59538 4972 59544 4984
rect 59596 4972 59602 5024
rect 65168 5012 65196 5108
rect 66346 5040 66352 5092
rect 66404 5080 66410 5092
rect 67177 5083 67235 5089
rect 67177 5080 67189 5083
rect 66404 5052 67189 5080
rect 66404 5040 66410 5052
rect 67177 5049 67189 5052
rect 67223 5049 67235 5083
rect 67177 5043 67235 5049
rect 68097 5083 68155 5089
rect 68097 5049 68109 5083
rect 68143 5080 68155 5083
rect 68738 5080 68744 5092
rect 68143 5052 68744 5080
rect 68143 5049 68155 5052
rect 68097 5043 68155 5049
rect 68738 5040 68744 5052
rect 68796 5040 68802 5092
rect 66990 5012 66996 5024
rect 65168 4984 66996 5012
rect 66990 4972 66996 4984
rect 67048 4972 67054 5024
rect 67269 5015 67327 5021
rect 67269 4981 67281 5015
rect 67315 5012 67327 5015
rect 69658 5012 69664 5024
rect 67315 4984 69664 5012
rect 67315 4981 67327 4984
rect 67269 4975 67327 4981
rect 69658 4972 69664 4984
rect 69716 4972 69722 5024
rect 1104 4922 18952 4944
rect 1104 4870 9246 4922
rect 9298 4870 9310 4922
rect 9362 4870 9374 4922
rect 9426 4870 9438 4922
rect 9490 4870 18952 4922
rect 23842 4904 23848 4956
rect 23900 4944 23906 4956
rect 33042 4944 33048 4956
rect 23900 4916 33048 4944
rect 23900 4904 23906 4916
rect 33042 4904 33048 4916
rect 33100 4904 33106 4956
rect 37628 4922 68816 4944
rect 24486 4876 24492 4888
rect 1104 4848 18952 4870
rect 24447 4848 24492 4876
rect 24486 4836 24492 4848
rect 24544 4836 24550 4888
rect 31754 4836 31760 4888
rect 31812 4876 31818 4888
rect 32030 4876 32036 4888
rect 31812 4848 31857 4876
rect 31991 4848 32036 4876
rect 31812 4836 31818 4848
rect 32030 4836 32036 4848
rect 32088 4836 32094 4888
rect 32306 4876 32312 4888
rect 32267 4848 32312 4876
rect 32306 4836 32312 4848
rect 32364 4836 32370 4888
rect 32490 4876 32496 4888
rect 32451 4848 32496 4876
rect 32490 4836 32496 4848
rect 32548 4836 32554 4888
rect 37628 4870 39246 4922
rect 39298 4870 39310 4922
rect 39362 4870 39374 4922
rect 39426 4870 39438 4922
rect 39490 4870 49246 4922
rect 49298 4870 49310 4922
rect 49362 4870 49374 4922
rect 49426 4870 49438 4922
rect 49490 4870 59246 4922
rect 59298 4870 59310 4922
rect 59362 4870 59374 4922
rect 59426 4870 59438 4922
rect 59490 4870 68816 4922
rect 37628 4848 68816 4870
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7742 4808 7748 4820
rect 7064 4780 7748 4808
rect 7064 4768 7070 4780
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 10836 4780 14412 4808
rect 10836 4768 10842 4780
rect 1949 4743 2007 4749
rect 1949 4709 1961 4743
rect 1995 4740 2007 4743
rect 3970 4740 3976 4752
rect 1995 4712 3976 4740
rect 1995 4709 2007 4712
rect 1949 4703 2007 4709
rect 3970 4700 3976 4712
rect 4028 4700 4034 4752
rect 13630 4740 13636 4752
rect 11900 4712 13636 4740
rect 11900 4684 11928 4712
rect 13630 4700 13636 4712
rect 13688 4700 13694 4752
rect 2498 4672 2504 4684
rect 1964 4644 2504 4672
rect 1964 4616 1992 4644
rect 2498 4632 2504 4644
rect 2556 4672 2562 4684
rect 2685 4675 2743 4681
rect 2685 4672 2697 4675
rect 2556 4644 2697 4672
rect 2556 4632 2562 4644
rect 2685 4641 2697 4644
rect 2731 4641 2743 4675
rect 2685 4635 2743 4641
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 3234 4672 3240 4684
rect 3191 4644 3240 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 4614 4672 4620 4684
rect 4575 4644 4620 4672
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 5040 4644 5273 4672
rect 5040 4632 5046 4644
rect 5261 4641 5273 4644
rect 5307 4641 5319 4675
rect 5718 4672 5724 4684
rect 5679 4644 5724 4672
rect 5261 4635 5319 4641
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 6052 4644 6377 4672
rect 6052 4632 6058 4644
rect 6365 4641 6377 4644
rect 6411 4641 6423 4675
rect 7006 4672 7012 4684
rect 6919 4644 7012 4672
rect 6365 4635 6423 4641
rect 7006 4632 7012 4644
rect 7064 4672 7070 4684
rect 7374 4672 7380 4684
rect 7064 4644 7380 4672
rect 7064 4632 7070 4644
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 7616 4644 7665 4672
rect 7616 4632 7622 4644
rect 7653 4641 7665 4644
rect 7699 4672 7711 4675
rect 7926 4672 7932 4684
rect 7699 4644 7932 4672
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 8754 4672 8760 4684
rect 8619 4644 8760 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 8754 4632 8760 4644
rect 8812 4672 8818 4684
rect 9214 4672 9220 4684
rect 8812 4644 9220 4672
rect 8812 4632 8818 4644
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9582 4632 9588 4684
rect 9640 4672 9646 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9640 4644 9689 4672
rect 9640 4632 9646 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 10778 4672 10784 4684
rect 10643 4644 10784 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 11241 4675 11299 4681
rect 11241 4641 11253 4675
rect 11287 4672 11299 4675
rect 11422 4672 11428 4684
rect 11287 4644 11428 4672
rect 11287 4641 11299 4644
rect 11241 4635 11299 4641
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 11882 4672 11888 4684
rect 11843 4644 11888 4672
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12308 4644 12541 4672
rect 12308 4632 12314 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13538 4672 13544 4684
rect 13219 4644 13544 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 1946 4564 1952 4616
rect 2004 4564 2010 4616
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 3878 4468 3884 4480
rect 3839 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 12544 4468 12572 4635
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 13817 4675 13875 4681
rect 13817 4641 13829 4675
rect 13863 4672 13875 4675
rect 14090 4672 14096 4684
rect 13863 4644 14096 4672
rect 13863 4641 13875 4644
rect 13817 4635 13875 4641
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 14384 4672 14412 4780
rect 14660 4780 16160 4808
rect 14660 4672 14688 4780
rect 14921 4743 14979 4749
rect 14921 4709 14933 4743
rect 14967 4740 14979 4743
rect 16022 4740 16028 4752
rect 14967 4712 16028 4740
rect 14967 4709 14979 4712
rect 14921 4703 14979 4709
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 16132 4740 16160 4780
rect 16482 4768 16488 4820
rect 16540 4808 16546 4820
rect 51902 4808 51908 4820
rect 16540 4780 51908 4808
rect 16540 4768 16546 4780
rect 51902 4768 51908 4780
rect 51960 4808 51966 4820
rect 52270 4808 52276 4820
rect 51960 4780 52276 4808
rect 51960 4768 51966 4780
rect 52270 4768 52276 4780
rect 52328 4768 52334 4820
rect 62666 4768 62672 4820
rect 62724 4808 62730 4820
rect 62724 4780 68048 4808
rect 62724 4768 62730 4780
rect 16132 4712 16988 4740
rect 14384 4644 14688 4672
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15252 4644 15669 4672
rect 15252 4632 15258 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 16356 4644 16405 4672
rect 16356 4632 16362 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 16666 4604 16672 4616
rect 13412 4576 16672 4604
rect 13412 4564 13418 4576
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 14642 4496 14648 4548
rect 14700 4536 14706 4548
rect 14737 4539 14795 4545
rect 14737 4536 14749 4539
rect 14700 4508 14749 4536
rect 14700 4496 14706 4508
rect 14737 4505 14749 4508
rect 14783 4505 14795 4539
rect 14737 4499 14795 4505
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 15473 4539 15531 4545
rect 15473 4536 15485 4539
rect 15252 4508 15485 4536
rect 15252 4496 15258 4508
rect 15473 4505 15485 4508
rect 15519 4505 15531 4539
rect 16850 4536 16856 4548
rect 16811 4508 16856 4536
rect 15473 4499 15531 4505
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 16960 4536 16988 4712
rect 17218 4700 17224 4752
rect 17276 4740 17282 4752
rect 59354 4740 59360 4752
rect 17276 4712 59360 4740
rect 17276 4700 17282 4712
rect 59354 4700 59360 4712
rect 59412 4700 59418 4752
rect 60642 4700 60648 4752
rect 60700 4740 60706 4752
rect 68020 4749 68048 4780
rect 67177 4743 67235 4749
rect 67177 4740 67189 4743
rect 60700 4712 67189 4740
rect 60700 4700 60706 4712
rect 67177 4709 67189 4712
rect 67223 4709 67235 4743
rect 67177 4703 67235 4709
rect 68005 4743 68063 4749
rect 68005 4709 68017 4743
rect 68051 4709 68063 4743
rect 68005 4703 68063 4709
rect 17037 4675 17095 4681
rect 17037 4641 17049 4675
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 18782 4672 18788 4684
rect 18095 4644 18788 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 17052 4604 17080 4635
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 23750 4632 23756 4684
rect 23808 4672 23814 4684
rect 24394 4672 24400 4684
rect 23808 4644 24400 4672
rect 23808 4632 23814 4644
rect 24394 4632 24400 4644
rect 24452 4632 24458 4684
rect 31938 4672 31944 4684
rect 31899 4644 31944 4672
rect 31938 4632 31944 4644
rect 31996 4632 32002 4684
rect 37550 4632 37556 4684
rect 37608 4672 37614 4684
rect 38473 4675 38531 4681
rect 38473 4672 38485 4675
rect 37608 4644 38485 4672
rect 37608 4632 37614 4644
rect 38473 4641 38485 4644
rect 38519 4641 38531 4675
rect 38473 4635 38531 4641
rect 39209 4675 39267 4681
rect 39209 4641 39221 4675
rect 39255 4672 39267 4675
rect 39666 4672 39672 4684
rect 39255 4644 39672 4672
rect 39255 4641 39267 4644
rect 39209 4635 39267 4641
rect 39666 4632 39672 4644
rect 39724 4632 39730 4684
rect 39850 4672 39856 4684
rect 39811 4644 39856 4672
rect 39850 4632 39856 4644
rect 39908 4632 39914 4684
rect 40957 4675 41015 4681
rect 40957 4641 40969 4675
rect 41003 4672 41015 4675
rect 41046 4672 41052 4684
rect 41003 4644 41052 4672
rect 41003 4641 41015 4644
rect 40957 4635 41015 4641
rect 41046 4632 41052 4644
rect 41104 4632 41110 4684
rect 42153 4675 42211 4681
rect 42153 4641 42165 4675
rect 42199 4672 42211 4675
rect 42610 4672 42616 4684
rect 42199 4644 42616 4672
rect 42199 4641 42211 4644
rect 42153 4635 42211 4641
rect 42610 4632 42616 4644
rect 42668 4632 42674 4684
rect 42886 4672 42892 4684
rect 42847 4644 42892 4672
rect 42886 4632 42892 4644
rect 42944 4632 42950 4684
rect 44729 4675 44787 4681
rect 44729 4672 44741 4675
rect 44008 4644 44741 4672
rect 18506 4604 18512 4616
rect 17052 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 34606 4564 34612 4616
rect 34664 4604 34670 4616
rect 44008 4604 44036 4644
rect 44729 4641 44741 4644
rect 44775 4672 44787 4675
rect 45922 4672 45928 4684
rect 44775 4644 45928 4672
rect 44775 4641 44787 4644
rect 44729 4635 44787 4641
rect 45922 4632 45928 4644
rect 45980 4632 45986 4684
rect 46106 4632 46112 4684
rect 46164 4672 46170 4684
rect 46201 4675 46259 4681
rect 46201 4672 46213 4675
rect 46164 4644 46213 4672
rect 46164 4632 46170 4644
rect 46201 4641 46213 4644
rect 46247 4641 46259 4675
rect 46201 4635 46259 4641
rect 46382 4632 46388 4684
rect 46440 4672 46446 4684
rect 46661 4675 46719 4681
rect 46661 4672 46673 4675
rect 46440 4644 46673 4672
rect 46440 4632 46446 4644
rect 46661 4641 46673 4644
rect 46707 4641 46719 4675
rect 47394 4672 47400 4684
rect 47355 4644 47400 4672
rect 46661 4635 46719 4641
rect 47394 4632 47400 4644
rect 47452 4632 47458 4684
rect 48038 4672 48044 4684
rect 47999 4644 48044 4672
rect 48038 4632 48044 4644
rect 48096 4632 48102 4684
rect 48130 4632 48136 4684
rect 48188 4672 48194 4684
rect 48501 4675 48559 4681
rect 48501 4672 48513 4675
rect 48188 4644 48513 4672
rect 48188 4632 48194 4644
rect 48501 4641 48513 4644
rect 48547 4641 48559 4675
rect 48501 4635 48559 4641
rect 49145 4675 49203 4681
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49234 4672 49240 4684
rect 49191 4644 49240 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49234 4632 49240 4644
rect 49292 4632 49298 4684
rect 49973 4675 50031 4681
rect 49973 4641 49985 4675
rect 50019 4672 50031 4675
rect 50338 4672 50344 4684
rect 50019 4644 50344 4672
rect 50019 4641 50031 4644
rect 49973 4635 50031 4641
rect 50338 4632 50344 4644
rect 50396 4672 50402 4684
rect 50798 4672 50804 4684
rect 50396 4644 50804 4672
rect 50396 4632 50402 4644
rect 50798 4632 50804 4644
rect 50856 4632 50862 4684
rect 51442 4672 51448 4684
rect 51403 4644 51448 4672
rect 51442 4632 51448 4644
rect 51500 4632 51506 4684
rect 52089 4675 52147 4681
rect 52089 4641 52101 4675
rect 52135 4672 52147 4675
rect 52178 4672 52184 4684
rect 52135 4644 52184 4672
rect 52135 4641 52147 4644
rect 52089 4635 52147 4641
rect 52178 4632 52184 4644
rect 52236 4632 52242 4684
rect 52822 4632 52828 4684
rect 52880 4672 52886 4684
rect 53190 4672 53196 4684
rect 52880 4644 53196 4672
rect 52880 4632 52886 4644
rect 53190 4632 53196 4644
rect 53248 4672 53254 4684
rect 53377 4675 53435 4681
rect 53377 4672 53389 4675
rect 53248 4644 53389 4672
rect 53248 4632 53254 4644
rect 53377 4641 53389 4644
rect 53423 4641 53435 4675
rect 53377 4635 53435 4641
rect 53926 4632 53932 4684
rect 53984 4672 53990 4684
rect 54021 4675 54079 4681
rect 54021 4672 54033 4675
rect 53984 4644 54033 4672
rect 53984 4632 53990 4644
rect 54021 4641 54033 4644
rect 54067 4641 54079 4675
rect 54021 4635 54079 4641
rect 54570 4632 54576 4684
rect 54628 4672 54634 4684
rect 54665 4675 54723 4681
rect 54665 4672 54677 4675
rect 54628 4644 54677 4672
rect 54628 4632 54634 4644
rect 54665 4641 54677 4644
rect 54711 4641 54723 4675
rect 54665 4635 54723 4641
rect 55398 4632 55404 4684
rect 55456 4672 55462 4684
rect 55585 4675 55643 4681
rect 55585 4672 55597 4675
rect 55456 4644 55597 4672
rect 55456 4632 55462 4644
rect 55585 4641 55597 4644
rect 55631 4672 55643 4675
rect 56134 4672 56140 4684
rect 55631 4644 56140 4672
rect 55631 4641 55643 4644
rect 55585 4635 55643 4641
rect 56134 4632 56140 4644
rect 56192 4632 56198 4684
rect 56686 4632 56692 4684
rect 56744 4672 56750 4684
rect 56870 4672 56876 4684
rect 56744 4644 56876 4672
rect 56744 4632 56750 4644
rect 56870 4632 56876 4644
rect 56928 4632 56934 4684
rect 57054 4632 57060 4684
rect 57112 4672 57118 4684
rect 57514 4672 57520 4684
rect 57112 4644 57520 4672
rect 57112 4632 57118 4644
rect 57514 4632 57520 4644
rect 57572 4632 57578 4684
rect 57882 4632 57888 4684
rect 57940 4672 57946 4684
rect 57977 4675 58035 4681
rect 57977 4672 57989 4675
rect 57940 4644 57989 4672
rect 57940 4632 57946 4644
rect 57977 4641 57989 4644
rect 58023 4641 58035 4675
rect 57977 4635 58035 4641
rect 58618 4632 58624 4684
rect 58676 4672 58682 4684
rect 58805 4675 58863 4681
rect 58805 4672 58817 4675
rect 58676 4644 58817 4672
rect 58676 4632 58682 4644
rect 58805 4641 58817 4644
rect 58851 4672 58863 4675
rect 58894 4672 58900 4684
rect 58851 4644 58900 4672
rect 58851 4641 58863 4644
rect 58805 4635 58863 4641
rect 58894 4632 58900 4644
rect 58952 4632 58958 4684
rect 59722 4672 59728 4684
rect 59635 4644 59728 4672
rect 59722 4632 59728 4644
rect 59780 4672 59786 4684
rect 60090 4672 60096 4684
rect 59780 4644 60096 4672
rect 59780 4632 59786 4644
rect 60090 4632 60096 4644
rect 60148 4632 60154 4684
rect 62390 4672 62396 4684
rect 62351 4644 62396 4672
rect 62390 4632 62396 4644
rect 62448 4632 62454 4684
rect 62482 4632 62488 4684
rect 62540 4672 62546 4684
rect 63221 4675 63279 4681
rect 63221 4672 63233 4675
rect 62540 4644 63233 4672
rect 62540 4632 62546 4644
rect 63221 4641 63233 4644
rect 63267 4672 63279 4675
rect 63310 4672 63316 4684
rect 63267 4644 63316 4672
rect 63267 4641 63279 4644
rect 63221 4635 63279 4641
rect 63310 4632 63316 4644
rect 63368 4632 63374 4684
rect 63862 4632 63868 4684
rect 63920 4672 63926 4684
rect 64049 4675 64107 4681
rect 64049 4672 64061 4675
rect 63920 4644 64061 4672
rect 63920 4632 63926 4644
rect 64049 4641 64061 4644
rect 64095 4672 64107 4675
rect 64138 4672 64144 4684
rect 64095 4644 64144 4672
rect 64095 4641 64107 4644
rect 64049 4635 64107 4641
rect 64138 4632 64144 4644
rect 64196 4632 64202 4684
rect 64690 4672 64696 4684
rect 64651 4644 64696 4672
rect 64690 4632 64696 4644
rect 64748 4632 64754 4684
rect 64782 4632 64788 4684
rect 64840 4672 64846 4684
rect 65153 4675 65211 4681
rect 65153 4672 65165 4675
rect 64840 4644 65165 4672
rect 64840 4632 64846 4644
rect 65153 4641 65165 4644
rect 65199 4641 65211 4675
rect 65153 4635 65211 4641
rect 65242 4632 65248 4684
rect 65300 4672 65306 4684
rect 65981 4675 66039 4681
rect 65981 4672 65993 4675
rect 65300 4644 65993 4672
rect 65300 4632 65306 4644
rect 65981 4641 65993 4644
rect 66027 4641 66039 4675
rect 65981 4635 66039 4641
rect 34664 4576 44036 4604
rect 44085 4607 44143 4613
rect 34664 4564 34670 4576
rect 44085 4573 44097 4607
rect 44131 4604 44143 4607
rect 60182 4604 60188 4616
rect 44131 4576 60188 4604
rect 44131 4573 44143 4576
rect 44085 4567 44143 4573
rect 60182 4564 60188 4576
rect 60240 4604 60246 4616
rect 60642 4604 60648 4616
rect 60240 4576 60648 4604
rect 60240 4564 60246 4576
rect 60642 4564 60648 4576
rect 60700 4564 60706 4616
rect 17034 4536 17040 4548
rect 16960 4508 17040 4536
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 17218 4496 17224 4548
rect 17276 4536 17282 4548
rect 17586 4536 17592 4548
rect 17276 4508 17592 4536
rect 17276 4496 17282 4508
rect 17586 4496 17592 4508
rect 17644 4496 17650 4548
rect 18233 4539 18291 4545
rect 18233 4505 18245 4539
rect 18279 4536 18291 4539
rect 21450 4536 21456 4548
rect 18279 4508 21456 4536
rect 18279 4505 18291 4508
rect 18233 4499 18291 4505
rect 21450 4496 21456 4508
rect 21508 4496 21514 4548
rect 28629 4539 28687 4545
rect 28629 4505 28641 4539
rect 28675 4536 28687 4539
rect 34977 4539 35035 4545
rect 34977 4536 34989 4539
rect 28675 4508 34989 4536
rect 28675 4505 28687 4508
rect 28629 4499 28687 4505
rect 34977 4505 34989 4508
rect 35023 4505 35035 4539
rect 34977 4499 35035 4505
rect 35066 4496 35072 4548
rect 35124 4536 35130 4548
rect 38289 4539 38347 4545
rect 38289 4536 38301 4539
rect 35124 4508 38301 4536
rect 35124 4496 35130 4508
rect 38289 4505 38301 4508
rect 38335 4505 38347 4539
rect 38289 4499 38347 4505
rect 38838 4496 38844 4548
rect 38896 4536 38902 4548
rect 38896 4508 39896 4536
rect 38896 4496 38902 4508
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 12544 4440 19257 4468
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 34333 4471 34391 4477
rect 34333 4437 34345 4471
rect 34379 4468 34391 4471
rect 39117 4471 39175 4477
rect 39117 4468 39129 4471
rect 34379 4440 39129 4468
rect 34379 4437 34391 4440
rect 34333 4431 34391 4437
rect 39117 4437 39129 4440
rect 39163 4437 39175 4471
rect 39868 4468 39896 4508
rect 40218 4496 40224 4548
rect 40276 4536 40282 4548
rect 40773 4539 40831 4545
rect 40773 4536 40785 4539
rect 40276 4508 40785 4536
rect 40276 4496 40282 4508
rect 40773 4505 40785 4508
rect 40819 4505 40831 4539
rect 40773 4499 40831 4505
rect 41046 4496 41052 4548
rect 41104 4536 41110 4548
rect 41322 4536 41328 4548
rect 41104 4508 41328 4536
rect 41104 4496 41110 4508
rect 41322 4496 41328 4508
rect 41380 4536 41386 4548
rect 43349 4539 43407 4545
rect 43349 4536 43361 4539
rect 41380 4508 43361 4536
rect 41380 4496 41386 4508
rect 43349 4505 43361 4508
rect 43395 4505 43407 4539
rect 43349 4499 43407 4505
rect 43438 4496 43444 4548
rect 43496 4536 43502 4548
rect 46106 4536 46112 4548
rect 43496 4508 46112 4536
rect 43496 4496 43502 4508
rect 46106 4496 46112 4508
rect 46164 4496 46170 4548
rect 46198 4496 46204 4548
rect 46256 4536 46262 4548
rect 61749 4539 61807 4545
rect 61749 4536 61761 4539
rect 46256 4508 61761 4536
rect 46256 4496 46262 4508
rect 61749 4505 61761 4508
rect 61795 4505 61807 4539
rect 61749 4499 61807 4505
rect 64230 4496 64236 4548
rect 64288 4496 64294 4548
rect 67818 4536 67824 4548
rect 67779 4508 67824 4536
rect 67818 4496 67824 4508
rect 67876 4496 67882 4548
rect 42061 4471 42119 4477
rect 42061 4468 42073 4471
rect 39868 4440 42073 4468
rect 39117 4431 39175 4437
rect 42061 4437 42073 4440
rect 42107 4437 42119 4471
rect 42061 4431 42119 4437
rect 43070 4428 43076 4480
rect 43128 4468 43134 4480
rect 45646 4468 45652 4480
rect 43128 4440 45652 4468
rect 43128 4428 43134 4440
rect 45646 4428 45652 4440
rect 45704 4428 45710 4480
rect 46382 4428 46388 4480
rect 46440 4468 46446 4480
rect 46750 4468 46756 4480
rect 46440 4440 46756 4468
rect 46440 4428 46446 4440
rect 46750 4428 46756 4440
rect 46808 4428 46814 4480
rect 47670 4428 47676 4480
rect 47728 4468 47734 4480
rect 52733 4471 52791 4477
rect 52733 4468 52745 4471
rect 47728 4440 52745 4468
rect 47728 4428 47734 4440
rect 52733 4437 52745 4440
rect 52779 4437 52791 4471
rect 52733 4431 52791 4437
rect 53926 4428 53932 4480
rect 53984 4468 53990 4480
rect 54846 4468 54852 4480
rect 53984 4440 54852 4468
rect 53984 4428 53990 4440
rect 54846 4428 54852 4440
rect 54904 4428 54910 4480
rect 56226 4468 56232 4480
rect 56187 4440 56232 4468
rect 56226 4428 56232 4440
rect 56284 4428 56290 4480
rect 56870 4428 56876 4480
rect 56928 4468 56934 4480
rect 57882 4468 57888 4480
rect 56928 4440 57888 4468
rect 56928 4428 56934 4440
rect 57882 4428 57888 4440
rect 57940 4428 57946 4480
rect 59354 4428 59360 4480
rect 59412 4468 59418 4480
rect 60185 4471 60243 4477
rect 60185 4468 60197 4471
rect 59412 4440 60197 4468
rect 59412 4428 59418 4440
rect 60185 4437 60197 4440
rect 60231 4437 60243 4471
rect 60185 4431 60243 4437
rect 64046 4428 64052 4480
rect 64104 4468 64110 4480
rect 64248 4468 64276 4496
rect 64104 4440 64276 4468
rect 67269 4471 67327 4477
rect 64104 4428 64110 4440
rect 67269 4437 67281 4471
rect 67315 4468 67327 4471
rect 69106 4468 69112 4480
rect 67315 4440 69112 4468
rect 67315 4437 67327 4440
rect 67269 4431 67327 4437
rect 69106 4428 69112 4440
rect 69164 4428 69170 4480
rect 1104 4378 18952 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 14246 4378
rect 14298 4326 14310 4378
rect 14362 4326 14374 4378
rect 14426 4326 14438 4378
rect 14490 4326 18952 4378
rect 33042 4360 33048 4412
rect 33100 4400 33106 4412
rect 35158 4400 35164 4412
rect 33100 4372 35164 4400
rect 33100 4360 33106 4372
rect 35158 4360 35164 4372
rect 35216 4360 35222 4412
rect 37628 4378 68816 4400
rect 1104 4304 18952 4326
rect 37628 4326 44246 4378
rect 44298 4326 44310 4378
rect 44362 4326 44374 4378
rect 44426 4326 44438 4378
rect 44490 4326 54246 4378
rect 54298 4326 54310 4378
rect 54362 4326 54374 4378
rect 54426 4326 54438 4378
rect 54490 4326 64246 4378
rect 64298 4326 64310 4378
rect 64362 4326 64374 4378
rect 64426 4326 64438 4378
rect 64490 4326 68816 4378
rect 37628 4304 68816 4326
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 16574 4264 16580 4276
rect 11480 4236 16580 4264
rect 11480 4224 11486 4236
rect 16574 4224 16580 4236
rect 16632 4224 16638 4276
rect 16666 4224 16672 4276
rect 16724 4264 16730 4276
rect 18322 4264 18328 4276
rect 16724 4236 18328 4264
rect 16724 4224 16730 4236
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 23290 4224 23296 4276
rect 23348 4264 23354 4276
rect 40126 4264 40132 4276
rect 23348 4236 23428 4264
rect 23348 4224 23354 4236
rect 5905 4199 5963 4205
rect 5905 4165 5917 4199
rect 5951 4196 5963 4199
rect 6822 4196 6828 4208
rect 5951 4168 6828 4196
rect 5951 4165 5963 4168
rect 5905 4159 5963 4165
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 10962 4156 10968 4208
rect 11020 4196 11026 4208
rect 12158 4196 12164 4208
rect 11020 4168 12164 4196
rect 11020 4156 11026 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 13630 4156 13636 4208
rect 13688 4196 13694 4208
rect 19978 4196 19984 4208
rect 13688 4168 19984 4196
rect 13688 4156 13694 4168
rect 19978 4156 19984 4168
rect 20036 4156 20042 4208
rect 382 4088 388 4140
rect 440 4128 446 4140
rect 1486 4128 1492 4140
rect 440 4100 1492 4128
rect 440 4088 446 4100
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 3234 4128 3240 4140
rect 2188 4100 3240 4128
rect 2188 4088 2194 4100
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4614 4128 4620 4140
rect 4028 4100 4620 4128
rect 4028 4088 4034 4100
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5074 4128 5080 4140
rect 4724 4100 5080 4128
rect 842 4020 848 4072
rect 900 4060 906 4072
rect 1581 4063 1639 4069
rect 1581 4060 1593 4063
rect 900 4032 1593 4060
rect 900 4020 906 4032
rect 1581 4029 1593 4032
rect 1627 4060 1639 4063
rect 2222 4060 2228 4072
rect 1627 4032 2228 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 2222 4020 2228 4032
rect 2280 4020 2286 4072
rect 2406 4020 2412 4072
rect 2464 4020 2470 4072
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 2556 4032 2697 4060
rect 2556 4020 2562 4032
rect 2685 4029 2697 4032
rect 2731 4060 2743 4063
rect 3142 4060 3148 4072
rect 2731 4032 3148 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 566 3952 572 4004
rect 624 3992 630 4004
rect 1670 3992 1676 4004
rect 624 3964 1676 3992
rect 624 3952 630 3964
rect 1670 3952 1676 3964
rect 1728 3952 1734 4004
rect 2424 3992 2452 4020
rect 2240 3964 2452 3992
rect 2240 3936 2268 3964
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 3344 3992 3372 4023
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3786 4060 3792 4072
rect 3568 4032 3792 4060
rect 3568 4020 3574 4032
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 4724 4060 4752 4100
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 9490 4128 9496 4140
rect 8812 4100 9496 4128
rect 8812 4088 8818 4100
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 11422 4088 11428 4140
rect 11480 4128 11486 4140
rect 11882 4128 11888 4140
rect 11480 4100 11888 4128
rect 11480 4088 11486 4100
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12434 4128 12440 4140
rect 12032 4100 12440 4128
rect 12032 4088 12038 4100
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 12710 4088 12716 4140
rect 12768 4088 12774 4140
rect 18138 4128 18144 4140
rect 13004 4100 18144 4128
rect 5166 4060 5172 4072
rect 3896 4032 4752 4060
rect 5127 4032 5172 4060
rect 3896 3992 3924 4032
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6454 4060 6460 4072
rect 6328 4032 6460 4060
rect 6328 4020 6334 4032
rect 6454 4020 6460 4032
rect 6512 4060 6518 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6512 4032 6837 4060
rect 6512 4020 6518 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 7374 4060 7380 4072
rect 6972 4032 7380 4060
rect 6972 4020 6978 4032
rect 7374 4020 7380 4032
rect 7432 4060 7438 4072
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 7432 4032 7481 4060
rect 7432 4020 7438 4032
rect 7469 4029 7481 4032
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8386 4060 8392 4072
rect 7984 4032 8392 4060
rect 7984 4020 7990 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 9033 4063 9091 4069
rect 9033 4060 9045 4063
rect 8996 4032 9045 4060
rect 8996 4020 9002 4032
rect 9033 4029 9045 4032
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 10686 4060 10692 4072
rect 10551 4032 10692 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 3108 3964 3924 3992
rect 3108 3952 3114 3964
rect 4614 3952 4620 4004
rect 4672 3992 4678 4004
rect 4985 3995 5043 4001
rect 4985 3992 4997 3995
rect 4672 3964 4997 3992
rect 4672 3952 4678 3964
rect 4985 3961 4997 3964
rect 5031 3961 5043 3995
rect 4985 3955 5043 3961
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 8956 3992 8984 4020
rect 8260 3964 8984 3992
rect 8260 3952 8266 3964
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1946 3924 1952 3936
rect 992 3896 1952 3924
rect 992 3884 998 3896
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2222 3884 2228 3936
rect 2280 3884 2286 3936
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 3418 3924 3424 3936
rect 2464 3896 3424 3924
rect 2464 3884 2470 3896
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 9876 3924 9904 4023
rect 10686 4020 10692 4032
rect 10744 4060 10750 4072
rect 10870 4060 10876 4072
rect 10744 4032 10876 4060
rect 10744 4020 10750 4032
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4060 11207 4063
rect 11514 4060 11520 4072
rect 11195 4032 11520 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 12158 4020 12164 4072
rect 12216 4060 12222 4072
rect 12728 4060 12756 4088
rect 13004 4069 13032 4100
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 23290 4128 23296 4140
rect 19107 4100 23296 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 23290 4088 23296 4100
rect 23348 4088 23354 4140
rect 23400 4128 23428 4236
rect 31726 4236 40132 4264
rect 24946 4128 24952 4140
rect 23400 4100 24952 4128
rect 24946 4088 24952 4100
rect 25004 4088 25010 4140
rect 30561 4131 30619 4137
rect 30561 4097 30573 4131
rect 30607 4128 30619 4131
rect 31726 4128 31754 4236
rect 40126 4224 40132 4236
rect 40184 4224 40190 4276
rect 41782 4224 41788 4276
rect 41840 4264 41846 4276
rect 42518 4264 42524 4276
rect 41840 4236 42524 4264
rect 41840 4224 41846 4236
rect 42518 4224 42524 4236
rect 42576 4224 42582 4276
rect 42610 4224 42616 4276
rect 42668 4264 42674 4276
rect 42668 4236 45600 4264
rect 42668 4224 42674 4236
rect 32677 4199 32735 4205
rect 32677 4165 32689 4199
rect 32723 4196 32735 4199
rect 33134 4196 33140 4208
rect 32723 4168 33140 4196
rect 32723 4165 32735 4168
rect 32677 4159 32735 4165
rect 33134 4156 33140 4168
rect 33192 4156 33198 4208
rect 38562 4196 38568 4208
rect 35636 4168 38568 4196
rect 30607 4100 31754 4128
rect 30607 4097 30619 4100
rect 30561 4091 30619 4097
rect 32582 4088 32588 4140
rect 32640 4128 32646 4140
rect 35636 4128 35664 4168
rect 38562 4156 38568 4168
rect 38620 4156 38626 4208
rect 39025 4199 39083 4205
rect 39025 4165 39037 4199
rect 39071 4196 39083 4199
rect 39114 4196 39120 4208
rect 39071 4168 39120 4196
rect 39071 4165 39083 4168
rect 39025 4159 39083 4165
rect 39114 4156 39120 4168
rect 39172 4156 39178 4208
rect 42444 4168 44036 4196
rect 38102 4128 38108 4140
rect 32640 4100 35664 4128
rect 35728 4100 38108 4128
rect 32640 4088 32646 4100
rect 12216 4032 12756 4060
rect 12989 4063 13047 4069
rect 12216 4020 12222 4032
rect 12989 4029 13001 4063
rect 13035 4029 13047 4063
rect 14366 4060 14372 4072
rect 12989 4023 13047 4029
rect 13096 4032 14372 4060
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 11054 3992 11060 4004
rect 10836 3964 11060 3992
rect 10836 3952 10842 3964
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 11882 3952 11888 4004
rect 11940 3992 11946 4004
rect 12069 3995 12127 4001
rect 12069 3992 12081 3995
rect 11940 3964 12081 3992
rect 11940 3952 11946 3964
rect 12069 3961 12081 3964
rect 12115 3961 12127 3995
rect 12250 3992 12256 4004
rect 12211 3964 12256 3992
rect 12069 3955 12127 3961
rect 12250 3952 12256 3964
rect 12308 3952 12314 4004
rect 12710 3952 12716 4004
rect 12768 3992 12774 4004
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 12768 3964 12817 3992
rect 12768 3952 12774 3964
rect 12805 3961 12817 3964
rect 12851 3961 12863 3995
rect 12805 3955 12863 3961
rect 13096 3924 13124 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 15746 4060 15752 4072
rect 15427 4032 15752 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 17402 4060 17408 4072
rect 16255 4032 17408 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4060 17555 4063
rect 17586 4060 17592 4072
rect 17543 4032 17592 4060
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18690 4060 18696 4072
rect 18095 4032 18696 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19153 4063 19211 4069
rect 19153 4029 19165 4063
rect 19199 4060 19211 4063
rect 24670 4060 24676 4072
rect 19199 4032 24676 4060
rect 19199 4029 19211 4032
rect 19153 4023 19211 4029
rect 24670 4020 24676 4032
rect 24728 4020 24734 4072
rect 26881 4063 26939 4069
rect 26881 4029 26893 4063
rect 26927 4060 26939 4063
rect 33962 4060 33968 4072
rect 26927 4032 33968 4060
rect 26927 4029 26939 4032
rect 26881 4023 26939 4029
rect 33962 4020 33968 4032
rect 34020 4020 34026 4072
rect 13170 3952 13176 4004
rect 13228 3992 13234 4004
rect 13541 3995 13599 4001
rect 13541 3992 13553 3995
rect 13228 3964 13553 3992
rect 13228 3952 13234 3964
rect 13541 3961 13553 3964
rect 13587 3961 13599 3995
rect 13541 3955 13599 3961
rect 13725 3995 13783 4001
rect 13725 3961 13737 3995
rect 13771 3992 13783 3995
rect 13998 3992 14004 4004
rect 13771 3964 14004 3992
rect 13771 3961 13783 3964
rect 13725 3955 13783 3961
rect 13998 3952 14004 3964
rect 14056 3952 14062 4004
rect 14458 3992 14464 4004
rect 14419 3964 14464 3992
rect 14458 3952 14464 3964
rect 14516 3952 14522 4004
rect 16022 3992 16028 4004
rect 15983 3964 16028 3992
rect 16022 3952 16028 3964
rect 16080 3952 16086 4004
rect 18233 3995 18291 4001
rect 18233 3961 18245 3995
rect 18279 3992 18291 3995
rect 21542 3992 21548 4004
rect 18279 3964 21548 3992
rect 18279 3961 18291 3964
rect 18233 3955 18291 3961
rect 21542 3952 21548 3964
rect 21600 3952 21606 4004
rect 22646 3952 22652 4004
rect 22704 3992 22710 4004
rect 23842 3992 23848 4004
rect 22704 3964 23848 3992
rect 22704 3952 22710 3964
rect 23842 3952 23848 3964
rect 23900 3952 23906 4004
rect 28997 3995 29055 4001
rect 28997 3961 29009 3995
rect 29043 3992 29055 3995
rect 35728 3992 35756 4100
rect 38102 4088 38108 4100
rect 38160 4088 38166 4140
rect 38286 4088 38292 4140
rect 38344 4128 38350 4140
rect 41969 4131 42027 4137
rect 41969 4128 41981 4131
rect 38344 4100 41981 4128
rect 38344 4088 38350 4100
rect 41969 4097 41981 4100
rect 42015 4097 42027 4131
rect 41969 4091 42027 4097
rect 42058 4088 42064 4140
rect 42116 4128 42122 4140
rect 42444 4128 42472 4168
rect 42116 4100 42472 4128
rect 42116 4088 42122 4100
rect 42518 4088 42524 4140
rect 42576 4128 42582 4140
rect 43898 4128 43904 4140
rect 42576 4100 43904 4128
rect 42576 4088 42582 4100
rect 43898 4088 43904 4100
rect 43956 4088 43962 4140
rect 44008 4128 44036 4168
rect 45112 4168 45508 4196
rect 45112 4128 45140 4168
rect 44008 4100 45140 4128
rect 45186 4088 45192 4140
rect 45244 4128 45250 4140
rect 45244 4100 45416 4128
rect 45244 4088 45250 4100
rect 35805 4063 35863 4069
rect 35805 4029 35817 4063
rect 35851 4060 35863 4063
rect 38654 4060 38660 4072
rect 35851 4032 38660 4060
rect 35851 4029 35863 4032
rect 35805 4023 35863 4029
rect 38654 4020 38660 4032
rect 38712 4020 38718 4072
rect 39206 4060 39212 4072
rect 39167 4032 39212 4060
rect 39206 4020 39212 4032
rect 39264 4020 39270 4072
rect 39390 4020 39396 4072
rect 39448 4060 39454 4072
rect 39761 4063 39819 4069
rect 39761 4060 39773 4063
rect 39448 4032 39773 4060
rect 39448 4020 39454 4032
rect 39761 4029 39773 4032
rect 39807 4029 39819 4063
rect 39761 4023 39819 4029
rect 40126 4020 40132 4072
rect 40184 4060 40190 4072
rect 40310 4060 40316 4072
rect 40184 4032 40316 4060
rect 40184 4020 40190 4032
rect 40310 4020 40316 4032
rect 40368 4020 40374 4072
rect 40586 4020 40592 4072
rect 40644 4060 40650 4072
rect 40681 4063 40739 4069
rect 40681 4060 40693 4063
rect 40644 4032 40693 4060
rect 40644 4020 40650 4032
rect 40681 4029 40693 4032
rect 40727 4029 40739 4063
rect 40681 4023 40739 4029
rect 42153 4063 42211 4069
rect 42153 4029 42165 4063
rect 42199 4060 42211 4063
rect 42426 4060 42432 4072
rect 42199 4032 42432 4060
rect 42199 4029 42211 4032
rect 42153 4023 42211 4029
rect 42426 4020 42432 4032
rect 42484 4020 42490 4072
rect 43346 4020 43352 4072
rect 43404 4060 43410 4072
rect 44637 4063 44695 4069
rect 43404 4032 44588 4060
rect 43404 4020 43410 4032
rect 29043 3964 35756 3992
rect 37277 3995 37335 4001
rect 29043 3961 29055 3964
rect 28997 3955 29055 3961
rect 37277 3961 37289 3995
rect 37323 3992 37335 3995
rect 38289 3995 38347 4001
rect 38289 3992 38301 3995
rect 37323 3964 38301 3992
rect 37323 3961 37335 3964
rect 37277 3955 37335 3961
rect 38289 3961 38301 3964
rect 38335 3961 38347 3995
rect 38470 3992 38476 4004
rect 38431 3964 38476 3992
rect 38289 3955 38347 3961
rect 38470 3952 38476 3964
rect 38528 3952 38534 4004
rect 38562 3952 38568 4004
rect 38620 3992 38626 4004
rect 38620 3964 38884 3992
rect 38620 3952 38626 3964
rect 4571 3896 13124 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 14369 3927 14427 3933
rect 14369 3924 14381 3927
rect 13688 3896 14381 3924
rect 13688 3884 13694 3896
rect 14369 3893 14381 3896
rect 14415 3893 14427 3927
rect 14369 3887 14427 3893
rect 15473 3927 15531 3933
rect 15473 3893 15485 3927
rect 15519 3924 15531 3927
rect 18966 3924 18972 3936
rect 15519 3896 18972 3924
rect 15519 3893 15531 3896
rect 15473 3887 15531 3893
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19610 3884 19616 3936
rect 19668 3924 19674 3936
rect 21266 3924 21272 3936
rect 19668 3896 21272 3924
rect 19668 3884 19674 3896
rect 21266 3884 21272 3896
rect 21324 3884 21330 3936
rect 21726 3884 21732 3936
rect 21784 3924 21790 3936
rect 24762 3924 24768 3936
rect 21784 3896 24768 3924
rect 21784 3884 21790 3896
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 27893 3927 27951 3933
rect 27893 3893 27905 3927
rect 27939 3924 27951 3927
rect 35713 3927 35771 3933
rect 35713 3924 35725 3927
rect 27939 3896 35725 3924
rect 27939 3893 27951 3896
rect 27893 3887 27951 3893
rect 35713 3893 35725 3896
rect 35759 3893 35771 3927
rect 38746 3924 38752 3936
rect 35713 3887 35771 3893
rect 37016 3896 38752 3924
rect 1104 3834 18952 3856
rect 1104 3782 9246 3834
rect 9298 3782 9310 3834
rect 9362 3782 9374 3834
rect 9426 3782 9438 3834
rect 9490 3782 18952 3834
rect 19334 3816 19340 3868
rect 19392 3856 19398 3868
rect 21358 3856 21364 3868
rect 19392 3828 21364 3856
rect 19392 3816 19398 3828
rect 21358 3816 21364 3828
rect 21416 3816 21422 3868
rect 22554 3816 22560 3868
rect 22612 3856 22618 3868
rect 24302 3856 24308 3868
rect 22612 3828 24308 3856
rect 22612 3816 22618 3828
rect 24302 3816 24308 3828
rect 24360 3816 24366 3868
rect 30285 3859 30343 3865
rect 30285 3825 30297 3859
rect 30331 3856 30343 3859
rect 37016 3856 37044 3896
rect 38746 3884 38752 3896
rect 38804 3884 38810 3936
rect 38856 3924 38884 3964
rect 39666 3952 39672 4004
rect 39724 3992 39730 4004
rect 39945 3995 40003 4001
rect 39945 3992 39957 3995
rect 39724 3964 39957 3992
rect 39724 3952 39730 3964
rect 39945 3961 39957 3964
rect 39991 3961 40003 3995
rect 39945 3955 40003 3961
rect 40034 3952 40040 4004
rect 40092 3992 40098 4004
rect 41233 3995 41291 4001
rect 41233 3992 41245 3995
rect 40092 3964 41245 3992
rect 40092 3952 40098 3964
rect 41233 3961 41245 3964
rect 41279 3961 41291 3995
rect 41233 3955 41291 3961
rect 41417 3995 41475 4001
rect 41417 3961 41429 3995
rect 41463 3992 41475 3995
rect 42242 3992 42248 4004
rect 41463 3964 42248 3992
rect 41463 3961 41475 3964
rect 41417 3955 41475 3961
rect 42242 3952 42248 3964
rect 42300 3952 42306 4004
rect 43533 3995 43591 4001
rect 43533 3961 43545 3995
rect 43579 3961 43591 3995
rect 43533 3955 43591 3961
rect 40589 3927 40647 3933
rect 40589 3924 40601 3927
rect 38856 3896 40601 3924
rect 40589 3893 40601 3896
rect 40635 3893 40647 3927
rect 40589 3887 40647 3893
rect 41506 3884 41512 3936
rect 41564 3924 41570 3936
rect 43441 3927 43499 3933
rect 43441 3924 43453 3927
rect 41564 3896 43453 3924
rect 41564 3884 41570 3896
rect 43441 3893 43453 3896
rect 43487 3893 43499 3927
rect 43548 3924 43576 3955
rect 43622 3952 43628 4004
rect 43680 3992 43686 4004
rect 44453 3995 44511 4001
rect 44453 3992 44465 3995
rect 43680 3964 44465 3992
rect 43680 3952 43686 3964
rect 44453 3961 44465 3964
rect 44499 3961 44511 3995
rect 44453 3955 44511 3961
rect 43714 3924 43720 3936
rect 43548 3896 43720 3924
rect 43441 3887 43499 3893
rect 43714 3884 43720 3896
rect 43772 3884 43778 3936
rect 44560 3924 44588 4032
rect 44637 4029 44649 4063
rect 44683 4060 44695 4063
rect 45278 4060 45284 4072
rect 44683 4032 45284 4060
rect 44683 4029 44695 4032
rect 44637 4023 44695 4029
rect 45278 4020 45284 4032
rect 45336 4020 45342 4072
rect 45388 4069 45416 4100
rect 45373 4063 45431 4069
rect 45373 4029 45385 4063
rect 45419 4029 45431 4063
rect 45480 4060 45508 4168
rect 45572 4128 45600 4236
rect 45646 4224 45652 4276
rect 45704 4264 45710 4276
rect 45830 4264 45836 4276
rect 45704 4236 45836 4264
rect 45704 4224 45710 4236
rect 45830 4224 45836 4236
rect 45888 4224 45894 4276
rect 46934 4224 46940 4276
rect 46992 4264 46998 4276
rect 50338 4264 50344 4276
rect 46992 4236 50344 4264
rect 46992 4224 46998 4236
rect 50338 4224 50344 4236
rect 50396 4224 50402 4276
rect 56226 4264 56232 4276
rect 55232 4236 56232 4264
rect 47578 4196 47584 4208
rect 46676 4168 47584 4196
rect 46676 4128 46704 4168
rect 47578 4156 47584 4168
rect 47636 4156 47642 4208
rect 48406 4156 48412 4208
rect 48464 4196 48470 4208
rect 49234 4196 49240 4208
rect 48464 4168 49240 4196
rect 48464 4156 48470 4168
rect 49234 4156 49240 4168
rect 49292 4156 49298 4208
rect 55232 4196 55260 4236
rect 56226 4224 56232 4236
rect 56284 4224 56290 4276
rect 63604 4236 63816 4264
rect 54772 4168 55260 4196
rect 45572 4100 46704 4128
rect 46017 4063 46075 4069
rect 46017 4060 46029 4063
rect 45480 4032 46029 4060
rect 45373 4023 45431 4029
rect 46017 4029 46029 4032
rect 46063 4060 46075 4063
rect 46566 4060 46572 4072
rect 46063 4032 46572 4060
rect 46063 4029 46075 4032
rect 46017 4023 46075 4029
rect 46566 4020 46572 4032
rect 46624 4020 46630 4072
rect 46676 4069 46704 4100
rect 48038 4088 48044 4140
rect 48096 4128 48102 4140
rect 49050 4128 49056 4140
rect 48096 4100 49056 4128
rect 48096 4088 48102 4100
rect 49050 4088 49056 4100
rect 49108 4088 49114 4140
rect 49786 4128 49792 4140
rect 49160 4100 49792 4128
rect 46661 4063 46719 4069
rect 46661 4029 46673 4063
rect 46707 4029 46719 4063
rect 46661 4023 46719 4029
rect 47118 4020 47124 4072
rect 47176 4060 47182 4072
rect 47305 4063 47363 4069
rect 47305 4060 47317 4063
rect 47176 4032 47317 4060
rect 47176 4020 47182 4032
rect 47305 4029 47317 4032
rect 47351 4029 47363 4063
rect 47305 4023 47363 4029
rect 47578 4020 47584 4072
rect 47636 4060 47642 4072
rect 48777 4063 48835 4069
rect 48777 4060 48789 4063
rect 47636 4032 48789 4060
rect 47636 4020 47642 4032
rect 48777 4029 48789 4032
rect 48823 4060 48835 4063
rect 49160 4060 49188 4100
rect 49786 4088 49792 4100
rect 49844 4088 49850 4140
rect 50614 4088 50620 4140
rect 50672 4128 50678 4140
rect 51166 4128 51172 4140
rect 50672 4100 51172 4128
rect 50672 4088 50678 4100
rect 51166 4088 51172 4100
rect 51224 4088 51230 4140
rect 52638 4128 52644 4140
rect 51368 4100 52644 4128
rect 48823 4032 49188 4060
rect 48823 4029 48835 4032
rect 48777 4023 48835 4029
rect 49234 4020 49240 4072
rect 49292 4060 49298 4072
rect 49878 4060 49884 4072
rect 49292 4032 49337 4060
rect 49839 4032 49884 4060
rect 49292 4020 49298 4032
rect 49878 4020 49884 4032
rect 49936 4020 49942 4072
rect 50706 4060 50712 4072
rect 50667 4032 50712 4060
rect 50706 4020 50712 4032
rect 50764 4020 50770 4072
rect 50798 4020 50804 4072
rect 50856 4060 50862 4072
rect 51368 4069 51396 4100
rect 52638 4088 52644 4100
rect 52696 4088 52702 4140
rect 54772 4128 54800 4168
rect 55858 4156 55864 4208
rect 55916 4156 55922 4208
rect 58069 4199 58127 4205
rect 58069 4165 58081 4199
rect 58115 4196 58127 4199
rect 58115 4168 60734 4196
rect 58115 4165 58127 4168
rect 58069 4159 58127 4165
rect 53208 4100 54800 4128
rect 51353 4063 51411 4069
rect 51353 4060 51365 4063
rect 50856 4032 51365 4060
rect 50856 4020 50862 4032
rect 51353 4029 51365 4032
rect 51399 4029 51411 4063
rect 51353 4023 51411 4029
rect 51997 4063 52055 4069
rect 51997 4029 52009 4063
rect 52043 4029 52055 4063
rect 51997 4023 52055 4029
rect 45830 3952 45836 4004
rect 45888 3992 45894 4004
rect 47486 3992 47492 4004
rect 45888 3964 47492 3992
rect 45888 3952 45894 3964
rect 47486 3952 47492 3964
rect 47544 3952 47550 4004
rect 48590 3952 48596 4004
rect 48648 3992 48654 4004
rect 49252 3992 49280 4020
rect 48648 3964 49280 3992
rect 48648 3952 48654 3964
rect 51534 3952 51540 4004
rect 51592 3992 51598 4004
rect 52012 3992 52040 4023
rect 52086 4020 52092 4072
rect 52144 4060 52150 4072
rect 52457 4063 52515 4069
rect 52457 4060 52469 4063
rect 52144 4032 52469 4060
rect 52144 4020 52150 4032
rect 52457 4029 52469 4032
rect 52503 4060 52515 4063
rect 52546 4060 52552 4072
rect 52503 4032 52552 4060
rect 52503 4029 52515 4032
rect 52457 4023 52515 4029
rect 52546 4020 52552 4032
rect 52604 4020 52610 4072
rect 53208 3992 53236 4100
rect 54846 4088 54852 4140
rect 54904 4128 54910 4140
rect 55490 4128 55496 4140
rect 54904 4100 55496 4128
rect 54904 4088 54910 4100
rect 55490 4088 55496 4100
rect 55548 4088 55554 4140
rect 55876 4128 55904 4156
rect 56318 4128 56324 4140
rect 55876 4100 56324 4128
rect 56318 4088 56324 4100
rect 56376 4088 56382 4140
rect 60706 4128 60734 4168
rect 63604 4128 63632 4236
rect 63678 4156 63684 4208
rect 63736 4156 63742 4208
rect 60706 4100 63632 4128
rect 53837 4063 53895 4069
rect 53837 4060 53849 4063
rect 53760 4032 53849 4060
rect 53760 4004 53788 4032
rect 53837 4029 53849 4032
rect 53883 4029 53895 4063
rect 53837 4023 53895 4029
rect 54481 4063 54539 4069
rect 54481 4029 54493 4063
rect 54527 4060 54539 4063
rect 54754 4060 54760 4072
rect 54527 4032 54760 4060
rect 54527 4029 54539 4032
rect 54481 4023 54539 4029
rect 54754 4020 54760 4032
rect 54812 4020 54818 4072
rect 55122 4060 55128 4072
rect 54864 4032 55128 4060
rect 51592 3964 53236 3992
rect 51592 3952 51598 3964
rect 53742 3952 53748 4004
rect 53800 3952 53806 4004
rect 45738 3924 45744 3936
rect 44560 3896 45744 3924
rect 45738 3884 45744 3896
rect 45796 3884 45802 3936
rect 45922 3884 45928 3936
rect 45980 3924 45986 3936
rect 47302 3924 47308 3936
rect 45980 3896 47308 3924
rect 45980 3884 45986 3896
rect 47302 3884 47308 3896
rect 47360 3884 47366 3936
rect 49050 3884 49056 3936
rect 49108 3924 49114 3936
rect 50154 3924 50160 3936
rect 49108 3896 50160 3924
rect 49108 3884 49114 3896
rect 50154 3884 50160 3896
rect 50212 3884 50218 3936
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 52178 3924 52184 3936
rect 51132 3896 52184 3924
rect 51132 3884 51138 3896
rect 52178 3884 52184 3896
rect 52236 3884 52242 3936
rect 53926 3884 53932 3936
rect 53984 3924 53990 3936
rect 54864 3924 54892 4032
rect 55122 4020 55128 4032
rect 55180 4020 55186 4072
rect 55582 4020 55588 4072
rect 55640 4060 55646 4072
rect 55769 4063 55827 4069
rect 55769 4060 55781 4063
rect 55640 4032 55781 4060
rect 55640 4020 55646 4032
rect 55769 4029 55781 4032
rect 55815 4029 55827 4063
rect 55769 4023 55827 4029
rect 55858 4020 55864 4072
rect 55916 4060 55922 4072
rect 56597 4063 56655 4069
rect 56597 4060 56609 4063
rect 55916 4032 56609 4060
rect 55916 4020 55922 4032
rect 56597 4029 56609 4032
rect 56643 4060 56655 4063
rect 56778 4060 56784 4072
rect 56643 4032 56784 4060
rect 56643 4029 56655 4032
rect 56597 4023 56655 4029
rect 56778 4020 56784 4032
rect 56836 4020 56842 4072
rect 57241 4063 57299 4069
rect 57241 4029 57253 4063
rect 57287 4060 57299 4063
rect 57698 4060 57704 4072
rect 57287 4032 57704 4060
rect 57287 4029 57299 4032
rect 57241 4023 57299 4029
rect 54938 3952 54944 4004
rect 54996 3992 55002 4004
rect 55600 3992 55628 4020
rect 54996 3964 55628 3992
rect 54996 3952 55002 3964
rect 56226 3952 56232 4004
rect 56284 3992 56290 4004
rect 57256 3992 57284 4023
rect 57698 4020 57704 4032
rect 57756 4020 57762 4072
rect 58250 4020 58256 4072
rect 58308 4060 58314 4072
rect 58802 4060 58808 4072
rect 58308 4032 58808 4060
rect 58308 4020 58314 4032
rect 58802 4020 58808 4032
rect 58860 4060 58866 4072
rect 59081 4063 59139 4069
rect 59081 4060 59093 4063
rect 58860 4032 59093 4060
rect 58860 4020 58866 4032
rect 59081 4029 59093 4032
rect 59127 4029 59139 4063
rect 59081 4023 59139 4029
rect 59170 4020 59176 4072
rect 59228 4060 59234 4072
rect 59725 4063 59783 4069
rect 59725 4060 59737 4063
rect 59228 4032 59737 4060
rect 59228 4020 59234 4032
rect 59725 4029 59737 4032
rect 59771 4060 59783 4063
rect 59814 4060 59820 4072
rect 59771 4032 59820 4060
rect 59771 4029 59783 4032
rect 59725 4023 59783 4029
rect 59814 4020 59820 4032
rect 59872 4020 59878 4072
rect 60458 4020 60464 4072
rect 60516 4060 60522 4072
rect 60645 4063 60703 4069
rect 60645 4060 60657 4063
rect 60516 4032 60657 4060
rect 60516 4020 60522 4032
rect 60645 4029 60657 4032
rect 60691 4029 60703 4063
rect 60645 4023 60703 4029
rect 61378 4020 61384 4072
rect 61436 4060 61442 4072
rect 61565 4063 61623 4069
rect 61565 4060 61577 4063
rect 61436 4032 61577 4060
rect 61436 4020 61442 4032
rect 61565 4029 61577 4032
rect 61611 4060 61623 4063
rect 61654 4060 61660 4072
rect 61611 4032 61660 4060
rect 61611 4029 61623 4032
rect 61565 4023 61623 4029
rect 61654 4020 61660 4032
rect 61712 4020 61718 4072
rect 62574 4020 62580 4072
rect 62632 4060 62638 4072
rect 62761 4063 62819 4069
rect 62761 4060 62773 4063
rect 62632 4032 62773 4060
rect 62632 4020 62638 4032
rect 62761 4029 62773 4032
rect 62807 4060 62819 4063
rect 62850 4060 62856 4072
rect 62807 4032 62856 4060
rect 62807 4029 62819 4032
rect 62761 4023 62819 4029
rect 62850 4020 62856 4032
rect 62908 4020 62914 4072
rect 63034 4020 63040 4072
rect 63092 4060 63098 4072
rect 63402 4060 63408 4072
rect 63092 4032 63408 4060
rect 63092 4020 63098 4032
rect 63402 4020 63408 4032
rect 63460 4020 63466 4072
rect 63696 4060 63724 4156
rect 63788 4128 63816 4236
rect 63788 4100 66024 4128
rect 65996 4069 66024 4100
rect 66162 4088 66168 4140
rect 66220 4128 66226 4140
rect 68186 4128 68192 4140
rect 66220 4100 68192 4128
rect 66220 4088 66226 4100
rect 68186 4088 68192 4100
rect 68244 4088 68250 4140
rect 64325 4063 64383 4069
rect 64325 4060 64337 4063
rect 63696 4032 64337 4060
rect 56284 3964 57284 3992
rect 56284 3952 56290 3964
rect 53984 3896 54892 3924
rect 53984 3884 53990 3896
rect 55582 3884 55588 3936
rect 55640 3924 55646 3936
rect 55950 3924 55956 3936
rect 55640 3896 55956 3924
rect 55640 3884 55646 3896
rect 55950 3884 55956 3896
rect 56008 3884 56014 3936
rect 58986 3884 58992 3936
rect 59044 3924 59050 3936
rect 62025 3927 62083 3933
rect 62025 3924 62037 3927
rect 59044 3896 62037 3924
rect 59044 3884 59050 3896
rect 62025 3893 62037 3896
rect 62071 3893 62083 3927
rect 62025 3887 62083 3893
rect 63586 3884 63592 3936
rect 63644 3924 63650 3936
rect 63696 3924 63724 4032
rect 64325 4029 64337 4032
rect 64371 4029 64383 4063
rect 64325 4023 64383 4029
rect 65429 4063 65487 4069
rect 65429 4029 65441 4063
rect 65475 4029 65487 4063
rect 65429 4023 65487 4029
rect 65981 4063 66039 4069
rect 65981 4029 65993 4063
rect 66027 4029 66039 4063
rect 65981 4023 66039 4029
rect 63644 3896 63724 3924
rect 65444 3924 65472 4023
rect 66070 4020 66076 4072
rect 66128 4060 66134 4072
rect 66809 4063 66867 4069
rect 66809 4060 66821 4063
rect 66128 4032 66821 4060
rect 66128 4020 66134 4032
rect 66809 4029 66821 4032
rect 66855 4029 66867 4063
rect 66809 4023 66867 4029
rect 66990 4020 66996 4072
rect 67048 4060 67054 4072
rect 68554 4060 68560 4072
rect 67048 4032 68560 4060
rect 67048 4020 67054 4032
rect 68554 4020 68560 4032
rect 68612 4020 68618 4072
rect 66622 3992 66628 4004
rect 66583 3964 66628 3992
rect 66622 3952 66628 3964
rect 66680 3952 66686 4004
rect 67450 3992 67456 4004
rect 67411 3964 67456 3992
rect 67450 3952 67456 3964
rect 67508 3952 67514 4004
rect 67637 3995 67695 4001
rect 67637 3961 67649 3995
rect 67683 3992 67695 3995
rect 68278 3992 68284 4004
rect 67683 3964 68284 3992
rect 67683 3961 67695 3964
rect 67637 3955 67695 3961
rect 68278 3952 68284 3964
rect 68336 3952 68342 4004
rect 65978 3924 65984 3936
rect 65444 3896 65984 3924
rect 63644 3884 63650 3896
rect 65978 3884 65984 3896
rect 66036 3884 66042 3936
rect 66073 3927 66131 3933
rect 66073 3893 66085 3927
rect 66119 3924 66131 3927
rect 69566 3924 69572 3936
rect 66119 3896 69572 3924
rect 66119 3893 66131 3896
rect 66073 3887 66131 3893
rect 69566 3884 69572 3896
rect 69624 3884 69630 3936
rect 30331 3828 37044 3856
rect 37628 3834 68816 3856
rect 30331 3825 30343 3828
rect 30285 3819 30343 3825
rect 1104 3760 18952 3782
rect 19426 3748 19432 3800
rect 19484 3788 19490 3800
rect 23382 3788 23388 3800
rect 19484 3760 23388 3788
rect 19484 3748 19490 3760
rect 23382 3748 23388 3760
rect 23440 3748 23446 3800
rect 23474 3748 23480 3800
rect 23532 3788 23538 3800
rect 23750 3788 23756 3800
rect 23532 3760 23756 3788
rect 23532 3748 23538 3760
rect 23750 3748 23756 3760
rect 23808 3748 23814 3800
rect 23934 3748 23940 3800
rect 23992 3788 23998 3800
rect 26513 3791 26571 3797
rect 26513 3788 26525 3791
rect 23992 3760 26525 3788
rect 23992 3748 23998 3760
rect 26513 3757 26525 3760
rect 26559 3757 26571 3791
rect 26513 3751 26571 3757
rect 31113 3791 31171 3797
rect 31113 3757 31125 3791
rect 31159 3788 31171 3791
rect 32398 3788 32404 3800
rect 31159 3760 32404 3788
rect 31159 3757 31171 3760
rect 31113 3751 31171 3757
rect 32398 3748 32404 3760
rect 32456 3748 32462 3800
rect 33321 3791 33379 3797
rect 33321 3757 33333 3791
rect 33367 3788 33379 3791
rect 35434 3788 35440 3800
rect 33367 3760 35440 3788
rect 33367 3757 33379 3760
rect 33321 3751 33379 3757
rect 35434 3748 35440 3760
rect 35492 3748 35498 3800
rect 37628 3782 39246 3834
rect 39298 3782 39310 3834
rect 39362 3782 39374 3834
rect 39426 3782 39438 3834
rect 39490 3782 49246 3834
rect 49298 3782 49310 3834
rect 49362 3782 49374 3834
rect 49426 3782 49438 3834
rect 49490 3782 59246 3834
rect 59298 3782 59310 3834
rect 59362 3782 59374 3834
rect 59426 3782 59438 3834
rect 59490 3782 68816 3834
rect 37628 3760 68816 3782
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2314 3720 2320 3732
rect 1728 3692 2320 3720
rect 1728 3680 1734 3692
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 4706 3720 4712 3732
rect 4448 3692 4712 3720
rect 3878 3652 3884 3664
rect 1596 3624 3884 3652
rect 1596 3596 1624 3624
rect 3878 3612 3884 3624
rect 3936 3612 3942 3664
rect 4448 3661 4476 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5718 3720 5724 3732
rect 5224 3692 5724 3720
rect 5224 3680 5230 3692
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 7558 3720 7564 3732
rect 6236 3692 7564 3720
rect 6236 3680 6242 3692
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 8386 3720 8392 3732
rect 7800 3692 8392 3720
rect 7800 3680 7806 3692
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 10560 3692 10609 3720
rect 10560 3680 10566 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 10597 3683 10655 3689
rect 14553 3723 14611 3729
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 15378 3720 15384 3732
rect 14599 3692 15384 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 18138 3720 18144 3732
rect 15764 3692 18144 3720
rect 4433 3655 4491 3661
rect 4433 3621 4445 3655
rect 4479 3621 4491 3655
rect 5626 3652 5632 3664
rect 5587 3624 5632 3652
rect 4433 3615 4491 3621
rect 5626 3612 5632 3624
rect 5684 3612 5690 3664
rect 6362 3652 6368 3664
rect 6323 3624 6368 3652
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 9309 3655 9367 3661
rect 9309 3621 9321 3655
rect 9355 3652 9367 3655
rect 11054 3652 11060 3664
rect 9355 3624 11060 3652
rect 9355 3621 9367 3624
rect 9309 3615 9367 3621
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 12621 3655 12679 3661
rect 12621 3621 12633 3655
rect 12667 3652 12679 3655
rect 13078 3652 13084 3664
rect 12667 3624 13084 3652
rect 12667 3621 12679 3624
rect 12621 3615 12679 3621
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 13354 3652 13360 3664
rect 13315 3624 13360 3652
rect 13354 3612 13360 3624
rect 13412 3612 13418 3664
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 15289 3655 15347 3661
rect 13596 3624 15240 3652
rect 13596 3612 13602 3624
rect 1578 3584 1584 3596
rect 1491 3556 1584 3584
rect 1578 3544 1584 3556
rect 1636 3544 1642 3596
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 2590 3584 2596 3596
rect 2271 3556 2596 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 14 3476 20 3528
rect 72 3516 78 3528
rect 1118 3516 1124 3528
rect 72 3488 1124 3516
rect 72 3476 78 3488
rect 1118 3476 1124 3488
rect 1176 3476 1182 3528
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 2240 3516 2268 3547
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2746 3556 2881 3584
rect 1452 3488 2268 3516
rect 1452 3476 1458 3488
rect 658 3408 664 3460
rect 716 3448 722 3460
rect 1762 3448 1768 3460
rect 716 3420 1768 3448
rect 716 3408 722 3420
rect 1762 3408 1768 3420
rect 1820 3408 1826 3460
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2746 3448 2774 3556
rect 2869 3553 2881 3556
rect 2915 3584 2927 3587
rect 3602 3584 3608 3596
rect 2915 3556 3608 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 6730 3584 6736 3596
rect 5644 3556 6736 3584
rect 5644 3528 5672 3556
rect 6730 3544 6736 3556
rect 6788 3584 6794 3596
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6788 3556 6929 3584
rect 6788 3544 6794 3556
rect 6917 3553 6929 3556
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 7650 3584 7656 3596
rect 7607 3556 7656 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 7576 3516 7604 3547
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 8018 3544 8024 3596
rect 8076 3584 8082 3596
rect 8205 3587 8263 3593
rect 8205 3584 8217 3587
rect 8076 3556 8217 3584
rect 8076 3544 8082 3556
rect 8205 3553 8217 3556
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3584 10011 3587
rect 10134 3584 10140 3596
rect 9999 3556 10140 3584
rect 9999 3553 10011 3556
rect 9953 3547 10011 3553
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11710 3587 11768 3593
rect 11710 3584 11722 3587
rect 11204 3556 11722 3584
rect 11204 3544 11210 3556
rect 11710 3553 11722 3556
rect 11756 3553 11768 3587
rect 15102 3584 15108 3596
rect 15063 3556 15108 3584
rect 11710 3547 11768 3553
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 15212 3584 15240 3624
rect 15289 3621 15301 3655
rect 15335 3652 15347 3655
rect 15764 3652 15792 3692
rect 18138 3680 18144 3692
rect 18196 3680 18202 3732
rect 18230 3680 18236 3732
rect 18288 3720 18294 3732
rect 18288 3692 20760 3720
rect 18288 3680 18294 3692
rect 15335 3624 15792 3652
rect 15841 3655 15899 3661
rect 15335 3621 15347 3624
rect 15289 3615 15347 3621
rect 15841 3621 15853 3655
rect 15887 3652 15899 3655
rect 16390 3652 16396 3664
rect 15887 3624 16396 3652
rect 15887 3621 15899 3624
rect 15841 3615 15899 3621
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 16577 3655 16635 3661
rect 16577 3621 16589 3655
rect 16623 3652 16635 3655
rect 17218 3652 17224 3664
rect 16623 3624 17224 3652
rect 16623 3621 16635 3624
rect 16577 3615 16635 3621
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 17954 3612 17960 3664
rect 18012 3652 18018 3664
rect 18049 3655 18107 3661
rect 18049 3652 18061 3655
rect 18012 3624 18061 3652
rect 18012 3612 18018 3624
rect 18049 3621 18061 3624
rect 18095 3621 18107 3655
rect 19702 3652 19708 3664
rect 18049 3615 18107 3621
rect 18156 3624 19708 3652
rect 16666 3584 16672 3596
rect 15212 3556 16672 3584
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 17368 3556 17413 3584
rect 17368 3544 17374 3556
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 18156 3584 18184 3624
rect 19702 3612 19708 3624
rect 19760 3612 19766 3664
rect 17920 3556 18184 3584
rect 18233 3587 18291 3593
rect 17920 3544 17926 3556
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 20622 3584 20628 3596
rect 18279 3556 20628 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 20732 3584 20760 3692
rect 20990 3680 20996 3732
rect 21048 3720 21054 3732
rect 22925 3723 22983 3729
rect 22925 3720 22937 3723
rect 21048 3692 22937 3720
rect 21048 3680 21054 3692
rect 22925 3689 22937 3692
rect 22971 3689 22983 3723
rect 22925 3683 22983 3689
rect 28721 3723 28779 3729
rect 28721 3689 28733 3723
rect 28767 3720 28779 3723
rect 33042 3720 33048 3732
rect 28767 3692 33048 3720
rect 28767 3689 28779 3692
rect 28721 3683 28779 3689
rect 33042 3680 33048 3692
rect 33100 3680 33106 3732
rect 33873 3723 33931 3729
rect 33873 3689 33885 3723
rect 33919 3720 33931 3723
rect 33962 3720 33968 3732
rect 33919 3692 33968 3720
rect 33919 3689 33931 3692
rect 33873 3683 33931 3689
rect 33962 3680 33968 3692
rect 34020 3680 34026 3732
rect 34149 3723 34207 3729
rect 34149 3689 34161 3723
rect 34195 3720 34207 3723
rect 35526 3720 35532 3732
rect 34195 3692 35532 3720
rect 34195 3689 34207 3692
rect 34149 3683 34207 3689
rect 35526 3680 35532 3692
rect 35584 3680 35590 3732
rect 37274 3680 37280 3732
rect 37332 3720 37338 3732
rect 38286 3720 38292 3732
rect 37332 3692 38292 3720
rect 37332 3680 37338 3692
rect 38286 3680 38292 3692
rect 38344 3680 38350 3732
rect 38562 3680 38568 3732
rect 38620 3720 38626 3732
rect 38620 3692 42748 3720
rect 38620 3680 38626 3692
rect 21634 3612 21640 3664
rect 21692 3652 21698 3664
rect 27157 3655 27215 3661
rect 27157 3652 27169 3655
rect 21692 3624 27169 3652
rect 21692 3612 21698 3624
rect 27157 3621 27169 3624
rect 27203 3621 27215 3655
rect 27157 3615 27215 3621
rect 27341 3655 27399 3661
rect 27341 3621 27353 3655
rect 27387 3652 27399 3655
rect 31573 3655 31631 3661
rect 31573 3652 31585 3655
rect 27387 3624 31585 3652
rect 27387 3621 27399 3624
rect 27341 3615 27399 3621
rect 31573 3621 31585 3624
rect 31619 3621 31631 3655
rect 31573 3615 31631 3621
rect 31662 3612 31668 3664
rect 31720 3652 31726 3664
rect 35805 3655 35863 3661
rect 35805 3652 35817 3655
rect 31720 3624 35817 3652
rect 31720 3612 31726 3624
rect 35805 3621 35817 3624
rect 35851 3621 35863 3655
rect 35805 3615 35863 3621
rect 36354 3612 36360 3664
rect 36412 3652 36418 3664
rect 37461 3655 37519 3661
rect 36412 3624 37320 3652
rect 36412 3612 36418 3624
rect 22557 3587 22615 3593
rect 22557 3584 22569 3587
rect 20732 3556 22569 3584
rect 22557 3553 22569 3556
rect 22603 3553 22615 3587
rect 22557 3547 22615 3553
rect 22646 3544 22652 3596
rect 22704 3584 22710 3596
rect 24210 3584 24216 3596
rect 22704 3556 24216 3584
rect 22704 3544 22710 3556
rect 24210 3544 24216 3556
rect 24268 3544 24274 3596
rect 30837 3587 30895 3593
rect 30837 3553 30849 3587
rect 30883 3584 30895 3587
rect 35066 3584 35072 3596
rect 30883 3556 35072 3584
rect 30883 3553 30895 3556
rect 30837 3547 30895 3553
rect 35066 3544 35072 3556
rect 35124 3544 35130 3596
rect 35158 3544 35164 3596
rect 35216 3584 35222 3596
rect 37182 3584 37188 3596
rect 35216 3556 37188 3584
rect 35216 3544 35222 3556
rect 37182 3544 37188 3556
rect 37240 3544 37246 3596
rect 37292 3584 37320 3624
rect 37461 3621 37473 3655
rect 37507 3652 37519 3655
rect 37550 3652 37556 3664
rect 37507 3624 37556 3652
rect 37507 3621 37519 3624
rect 37461 3615 37519 3621
rect 37550 3612 37556 3624
rect 37608 3612 37614 3664
rect 37642 3612 37648 3664
rect 37700 3652 37706 3664
rect 38473 3655 38531 3661
rect 38473 3652 38485 3655
rect 37700 3624 38485 3652
rect 37700 3612 37706 3624
rect 38473 3621 38485 3624
rect 38519 3621 38531 3655
rect 38473 3615 38531 3621
rect 38580 3624 39344 3652
rect 38580 3584 38608 3624
rect 39022 3584 39028 3596
rect 37292 3556 38608 3584
rect 38983 3556 39028 3584
rect 39022 3544 39028 3556
rect 39080 3544 39086 3596
rect 39206 3584 39212 3596
rect 39167 3556 39212 3584
rect 39206 3544 39212 3556
rect 39264 3544 39270 3596
rect 39316 3584 39344 3624
rect 40678 3612 40684 3664
rect 40736 3652 40742 3664
rect 40957 3655 41015 3661
rect 40957 3652 40969 3655
rect 40736 3624 40969 3652
rect 40736 3612 40742 3624
rect 40957 3621 40969 3624
rect 41003 3621 41015 3655
rect 42150 3652 42156 3664
rect 42111 3624 42156 3652
rect 40957 3615 41015 3621
rect 42150 3612 42156 3624
rect 42208 3612 42214 3664
rect 42720 3661 42748 3692
rect 42886 3680 42892 3732
rect 42944 3720 42950 3732
rect 44913 3723 44971 3729
rect 44913 3720 44925 3723
rect 42944 3692 44925 3720
rect 42944 3680 42950 3692
rect 44913 3689 44925 3692
rect 44959 3689 44971 3723
rect 44913 3683 44971 3689
rect 45186 3680 45192 3732
rect 45244 3720 45250 3732
rect 46382 3720 46388 3732
rect 45244 3692 46388 3720
rect 45244 3680 45250 3692
rect 46382 3680 46388 3692
rect 46440 3680 46446 3732
rect 47210 3680 47216 3732
rect 47268 3720 47274 3732
rect 48498 3720 48504 3732
rect 47268 3692 48504 3720
rect 47268 3680 47274 3692
rect 48498 3680 48504 3692
rect 48556 3680 48562 3732
rect 50154 3680 50160 3732
rect 50212 3720 50218 3732
rect 51442 3720 51448 3732
rect 50212 3692 51448 3720
rect 50212 3680 50218 3692
rect 51442 3680 51448 3692
rect 51500 3680 51506 3732
rect 61654 3680 61660 3732
rect 61712 3720 61718 3732
rect 62390 3720 62396 3732
rect 61712 3692 62396 3720
rect 61712 3680 61718 3692
rect 62390 3680 62396 3692
rect 62448 3680 62454 3732
rect 63954 3680 63960 3732
rect 64012 3720 64018 3732
rect 64012 3692 64276 3720
rect 64012 3680 64018 3692
rect 42705 3655 42763 3661
rect 42705 3621 42717 3655
rect 42751 3621 42763 3655
rect 44361 3655 44419 3661
rect 42705 3615 42763 3621
rect 42812 3624 43852 3652
rect 39316 3556 40816 3584
rect 6144 3488 7604 3516
rect 6144 3476 6150 3488
rect 2004 3420 2774 3448
rect 2004 3408 2010 3420
rect 3786 3408 3792 3460
rect 3844 3448 3850 3460
rect 4249 3451 4307 3457
rect 4249 3448 4261 3451
rect 3844 3420 4261 3448
rect 3844 3408 3850 3420
rect 4249 3417 4261 3420
rect 4295 3417 4307 3451
rect 4249 3411 4307 3417
rect 4798 3408 4804 3460
rect 4856 3448 4862 3460
rect 5445 3451 5503 3457
rect 5445 3448 5457 3451
rect 4856 3420 5457 3448
rect 4856 3408 4862 3420
rect 5445 3417 5457 3420
rect 5491 3417 5503 3451
rect 5445 3411 5503 3417
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 8036 3448 8064 3544
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 6972 3420 8064 3448
rect 6972 3408 6978 3420
rect 8938 3408 8944 3460
rect 8996 3448 9002 3460
rect 8996 3420 11100 3448
rect 8996 3408 9002 3420
rect 11072 3392 11100 3420
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 6273 3383 6331 3389
rect 6273 3380 6285 3383
rect 5132 3352 6285 3380
rect 5132 3340 5138 3352
rect 6273 3349 6285 3352
rect 6319 3349 6331 3383
rect 6273 3343 6331 3349
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8846 3380 8852 3392
rect 8076 3352 8852 3380
rect 8076 3340 8082 3352
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 9858 3380 9864 3392
rect 9819 3352 9864 3380
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 10594 3380 10600 3392
rect 10284 3352 10600 3380
rect 10284 3340 10290 3352
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 11054 3340 11060 3392
rect 11112 3340 11118 3392
rect 11992 3380 12020 3479
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12308 3488 12449 3516
rect 12308 3476 12314 3488
rect 12437 3485 12449 3488
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 15378 3476 15384 3528
rect 15436 3516 15442 3528
rect 15930 3516 15936 3528
rect 15436 3488 15936 3516
rect 15436 3476 15442 3488
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3516 16819 3519
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 16807 3488 20729 3516
rect 16807 3485 16819 3488
rect 16761 3479 16819 3485
rect 20717 3485 20729 3488
rect 20763 3485 20775 3519
rect 20717 3479 20775 3485
rect 20898 3476 20904 3528
rect 20956 3516 20962 3528
rect 23474 3516 23480 3528
rect 20956 3488 23480 3516
rect 20956 3476 20962 3488
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3516 30803 3519
rect 32677 3519 32735 3525
rect 32677 3516 32689 3519
rect 30791 3488 32689 3516
rect 30791 3485 30803 3488
rect 30745 3479 30803 3485
rect 32677 3485 32689 3488
rect 32723 3485 32735 3519
rect 32677 3479 32735 3485
rect 32766 3476 32772 3528
rect 32824 3516 32830 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 32824 3488 34897 3516
rect 32824 3476 32830 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 34977 3519 35035 3525
rect 34977 3485 34989 3519
rect 35023 3516 35035 3519
rect 37277 3519 37335 3525
rect 37277 3516 37289 3519
rect 35023 3488 37289 3516
rect 35023 3485 35035 3488
rect 34977 3479 35035 3485
rect 37277 3485 37289 3488
rect 37323 3485 37335 3519
rect 37277 3479 37335 3485
rect 37369 3519 37427 3525
rect 37369 3485 37381 3519
rect 37415 3516 37427 3519
rect 40788 3516 40816 3556
rect 40862 3544 40868 3596
rect 40920 3584 40926 3596
rect 42058 3584 42064 3596
rect 40920 3556 42064 3584
rect 40920 3544 40926 3556
rect 42058 3544 42064 3556
rect 42116 3544 42122 3596
rect 42334 3544 42340 3596
rect 42392 3584 42398 3596
rect 42812 3584 42840 3624
rect 42392 3556 42840 3584
rect 42889 3587 42947 3593
rect 42392 3544 42398 3556
rect 42889 3553 42901 3587
rect 42935 3584 42947 3587
rect 43254 3584 43260 3596
rect 42935 3556 43260 3584
rect 42935 3553 42947 3556
rect 42889 3547 42947 3553
rect 43254 3544 43260 3556
rect 43312 3544 43318 3596
rect 43625 3587 43683 3593
rect 43625 3553 43637 3587
rect 43671 3584 43683 3587
rect 43714 3584 43720 3596
rect 43671 3556 43720 3584
rect 43671 3553 43683 3556
rect 43625 3547 43683 3553
rect 43714 3544 43720 3556
rect 43772 3544 43778 3596
rect 43824 3584 43852 3624
rect 44361 3621 44373 3655
rect 44407 3652 44419 3655
rect 45462 3652 45468 3664
rect 44407 3624 45468 3652
rect 44407 3621 44419 3624
rect 44361 3615 44419 3621
rect 45462 3612 45468 3624
rect 45520 3612 45526 3664
rect 45646 3652 45652 3664
rect 45607 3624 45652 3652
rect 45646 3612 45652 3624
rect 45704 3612 45710 3664
rect 47118 3652 47124 3664
rect 46308 3624 47124 3652
rect 45094 3584 45100 3596
rect 43824 3556 45100 3584
rect 45094 3544 45100 3556
rect 45152 3544 45158 3596
rect 41969 3519 42027 3525
rect 41969 3516 41981 3519
rect 37415 3488 40724 3516
rect 40788 3488 41981 3516
rect 37415 3485 37427 3488
rect 37369 3479 37427 3485
rect 16025 3451 16083 3457
rect 16025 3417 16037 3451
rect 16071 3448 16083 3451
rect 16071 3420 19012 3448
rect 16071 3417 16083 3420
rect 16025 3411 16083 3417
rect 12434 3380 12440 3392
rect 11992 3352 12440 3380
rect 12434 3340 12440 3352
rect 12492 3340 12498 3392
rect 13265 3383 13323 3389
rect 13265 3349 13277 3383
rect 13311 3380 13323 3383
rect 13354 3380 13360 3392
rect 13311 3352 13360 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 17405 3383 17463 3389
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 17954 3380 17960 3392
rect 17451 3352 17960 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18984 3312 19012 3420
rect 19058 3408 19064 3460
rect 19116 3448 19122 3460
rect 22646 3448 22652 3460
rect 19116 3420 22652 3448
rect 19116 3408 19122 3420
rect 22646 3408 22652 3420
rect 22704 3408 22710 3460
rect 23658 3408 23664 3460
rect 23716 3448 23722 3460
rect 25869 3451 25927 3457
rect 25869 3448 25881 3451
rect 23716 3420 25881 3448
rect 23716 3408 23722 3420
rect 25869 3417 25881 3420
rect 25915 3417 25927 3451
rect 25869 3411 25927 3417
rect 30469 3451 30527 3457
rect 30469 3417 30481 3451
rect 30515 3448 30527 3451
rect 39114 3448 39120 3460
rect 30515 3420 39120 3448
rect 30515 3417 30527 3420
rect 30469 3411 30527 3417
rect 39114 3408 39120 3420
rect 39172 3408 39178 3460
rect 39206 3408 39212 3460
rect 39264 3448 39270 3460
rect 39482 3448 39488 3460
rect 39264 3420 39488 3448
rect 39264 3408 39270 3420
rect 39482 3408 39488 3420
rect 39540 3408 39546 3460
rect 40696 3448 40724 3488
rect 41969 3485 41981 3488
rect 42015 3485 42027 3519
rect 41969 3479 42027 3485
rect 42242 3476 42248 3528
rect 42300 3516 42306 3528
rect 42794 3516 42800 3528
rect 42300 3488 42800 3516
rect 42300 3476 42306 3488
rect 42794 3476 42800 3488
rect 42852 3476 42858 3528
rect 44818 3476 44824 3528
rect 44876 3516 44882 3528
rect 45738 3516 45744 3528
rect 44876 3488 45744 3516
rect 44876 3476 44882 3488
rect 45738 3476 45744 3488
rect 45796 3476 45802 3528
rect 40773 3451 40831 3457
rect 40773 3448 40785 3451
rect 40696 3420 40785 3448
rect 40773 3417 40785 3420
rect 40819 3417 40831 3451
rect 43441 3451 43499 3457
rect 43441 3448 43453 3451
rect 40773 3411 40831 3417
rect 40880 3420 43453 3448
rect 19150 3340 19156 3392
rect 19208 3380 19214 3392
rect 20898 3380 20904 3392
rect 19208 3352 20904 3380
rect 19208 3340 19214 3352
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 21450 3340 21456 3392
rect 21508 3380 21514 3392
rect 23934 3380 23940 3392
rect 21508 3352 23940 3380
rect 21508 3340 21514 3352
rect 23934 3340 23940 3352
rect 23992 3340 23998 3392
rect 29181 3383 29239 3389
rect 29181 3349 29193 3383
rect 29227 3380 29239 3383
rect 34977 3383 35035 3389
rect 34977 3380 34989 3383
rect 29227 3352 34989 3380
rect 29227 3349 29239 3352
rect 29181 3343 29239 3349
rect 34977 3349 34989 3352
rect 35023 3349 35035 3383
rect 38381 3383 38439 3389
rect 38381 3380 38393 3383
rect 34977 3343 35035 3349
rect 35084 3352 38393 3380
rect 25777 3315 25835 3321
rect 25777 3312 25789 3315
rect 1104 3290 18952 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 14246 3290
rect 14298 3238 14310 3290
rect 14362 3238 14374 3290
rect 14426 3238 14438 3290
rect 14490 3238 18952 3290
rect 18984 3284 25789 3312
rect 25777 3281 25789 3284
rect 25823 3281 25835 3315
rect 25777 3275 25835 3281
rect 27433 3315 27491 3321
rect 27433 3281 27445 3315
rect 27479 3312 27491 3315
rect 35084 3312 35112 3352
rect 38381 3349 38393 3352
rect 38427 3349 38439 3383
rect 38381 3343 38439 3349
rect 38746 3340 38752 3392
rect 38804 3380 38810 3392
rect 39761 3383 39819 3389
rect 39761 3380 39773 3383
rect 38804 3352 39773 3380
rect 38804 3340 38810 3352
rect 39761 3349 39773 3352
rect 39807 3349 39819 3383
rect 39761 3343 39819 3349
rect 39850 3340 39856 3392
rect 39908 3380 39914 3392
rect 40880 3380 40908 3420
rect 43441 3417 43453 3420
rect 43487 3417 43499 3451
rect 43441 3411 43499 3417
rect 43898 3408 43904 3460
rect 43956 3448 43962 3460
rect 46308 3448 46336 3624
rect 47118 3612 47124 3624
rect 47176 3612 47182 3664
rect 47670 3652 47676 3664
rect 47631 3624 47676 3652
rect 47670 3612 47676 3624
rect 47728 3612 47734 3664
rect 48130 3612 48136 3664
rect 48188 3652 48194 3664
rect 51994 3652 52000 3664
rect 48188 3624 49096 3652
rect 48188 3612 48194 3624
rect 46566 3544 46572 3596
rect 46624 3584 46630 3596
rect 46753 3587 46811 3593
rect 46753 3584 46765 3587
rect 46624 3556 46765 3584
rect 46624 3544 46630 3556
rect 46753 3553 46765 3556
rect 46799 3553 46811 3587
rect 48222 3584 48228 3596
rect 46753 3547 46811 3553
rect 46860 3556 48228 3584
rect 46382 3476 46388 3528
rect 46440 3516 46446 3528
rect 46860 3516 46888 3556
rect 48222 3544 48228 3556
rect 48280 3544 48286 3596
rect 48869 3587 48927 3593
rect 48869 3553 48881 3587
rect 48915 3584 48927 3587
rect 48958 3584 48964 3596
rect 48915 3556 48964 3584
rect 48915 3553 48927 3556
rect 48869 3547 48927 3553
rect 46440 3488 46888 3516
rect 46440 3476 46446 3488
rect 47302 3476 47308 3528
rect 47360 3516 47366 3528
rect 48884 3516 48912 3547
rect 48958 3544 48964 3556
rect 49016 3544 49022 3596
rect 49068 3584 49096 3624
rect 51046 3624 52000 3652
rect 49697 3587 49755 3593
rect 49697 3584 49709 3587
rect 49068 3556 49709 3584
rect 49697 3553 49709 3556
rect 49743 3584 49755 3587
rect 50062 3584 50068 3596
rect 49743 3556 50068 3584
rect 49743 3553 49755 3556
rect 49697 3547 49755 3553
rect 50062 3544 50068 3556
rect 50120 3544 50126 3596
rect 50341 3587 50399 3593
rect 50341 3553 50353 3587
rect 50387 3584 50399 3587
rect 51046 3584 51074 3624
rect 51994 3612 52000 3624
rect 52052 3612 52058 3664
rect 52733 3655 52791 3661
rect 52733 3621 52745 3655
rect 52779 3652 52791 3655
rect 53374 3652 53380 3664
rect 52779 3624 53380 3652
rect 52779 3621 52791 3624
rect 52733 3615 52791 3621
rect 53374 3612 53380 3624
rect 53432 3612 53438 3664
rect 54110 3612 54116 3664
rect 54168 3652 54174 3664
rect 54481 3655 54539 3661
rect 54481 3652 54493 3655
rect 54168 3624 54493 3652
rect 54168 3612 54174 3624
rect 54481 3621 54493 3624
rect 54527 3621 54539 3655
rect 54481 3615 54539 3621
rect 55309 3655 55367 3661
rect 55309 3621 55321 3655
rect 55355 3652 55367 3655
rect 55674 3652 55680 3664
rect 55355 3624 55680 3652
rect 55355 3621 55367 3624
rect 55309 3615 55367 3621
rect 55674 3612 55680 3624
rect 55732 3612 55738 3664
rect 56689 3655 56747 3661
rect 56689 3621 56701 3655
rect 56735 3652 56747 3655
rect 57146 3652 57152 3664
rect 56735 3624 57152 3652
rect 56735 3621 56747 3624
rect 56689 3615 56747 3621
rect 57146 3612 57152 3624
rect 57204 3612 57210 3664
rect 57422 3652 57428 3664
rect 57383 3624 57428 3652
rect 57422 3612 57428 3624
rect 57480 3612 57486 3664
rect 59538 3652 59544 3664
rect 59004 3624 59544 3652
rect 50387 3556 51074 3584
rect 50387 3553 50399 3556
rect 50341 3547 50399 3553
rect 47360 3488 48912 3516
rect 47360 3476 47366 3488
rect 49142 3476 49148 3528
rect 49200 3516 49206 3528
rect 50356 3516 50384 3547
rect 51258 3544 51264 3596
rect 51316 3584 51322 3596
rect 51445 3587 51503 3593
rect 51445 3584 51457 3587
rect 51316 3556 51457 3584
rect 51316 3544 51322 3556
rect 51445 3553 51457 3556
rect 51491 3553 51503 3587
rect 51445 3547 51503 3553
rect 51810 3544 51816 3596
rect 51868 3584 51874 3596
rect 51905 3587 51963 3593
rect 51905 3584 51917 3587
rect 51868 3556 51917 3584
rect 51868 3544 51874 3556
rect 51905 3553 51917 3556
rect 51951 3553 51963 3587
rect 51905 3547 51963 3553
rect 53006 3544 53012 3596
rect 53064 3584 53070 3596
rect 53561 3587 53619 3593
rect 53561 3584 53573 3587
rect 53064 3556 53573 3584
rect 53064 3544 53070 3556
rect 53561 3553 53573 3556
rect 53607 3553 53619 3587
rect 53561 3547 53619 3553
rect 57974 3544 57980 3596
rect 58032 3584 58038 3596
rect 58161 3587 58219 3593
rect 58161 3584 58173 3587
rect 58032 3556 58173 3584
rect 58032 3544 58038 3556
rect 58161 3553 58173 3556
rect 58207 3584 58219 3587
rect 58710 3584 58716 3596
rect 58207 3556 58716 3584
rect 58207 3553 58219 3556
rect 58161 3547 58219 3553
rect 58710 3544 58716 3556
rect 58768 3544 58774 3596
rect 58802 3544 58808 3596
rect 58860 3584 58866 3596
rect 59004 3593 59032 3624
rect 59538 3612 59544 3624
rect 59596 3612 59602 3664
rect 61746 3612 61752 3664
rect 61804 3612 61810 3664
rect 64248 3661 64276 3692
rect 65978 3680 65984 3732
rect 66036 3720 66042 3732
rect 66530 3720 66536 3732
rect 66036 3692 66536 3720
rect 66036 3680 66042 3692
rect 66530 3680 66536 3692
rect 66588 3680 66594 3732
rect 64233 3655 64291 3661
rect 64233 3621 64245 3655
rect 64279 3621 64291 3655
rect 64233 3615 64291 3621
rect 64874 3612 64880 3664
rect 64932 3652 64938 3664
rect 65061 3655 65119 3661
rect 65061 3652 65073 3655
rect 64932 3624 65073 3652
rect 64932 3612 64938 3624
rect 65061 3621 65073 3624
rect 65107 3621 65119 3655
rect 65061 3615 65119 3621
rect 65518 3612 65524 3664
rect 65576 3652 65582 3664
rect 65889 3655 65947 3661
rect 65889 3652 65901 3655
rect 65576 3624 65901 3652
rect 65576 3612 65582 3624
rect 65889 3621 65901 3624
rect 65935 3621 65947 3655
rect 65889 3615 65947 3621
rect 66806 3612 66812 3664
rect 66864 3652 66870 3664
rect 67177 3655 67235 3661
rect 67177 3652 67189 3655
rect 66864 3624 67189 3652
rect 66864 3612 66870 3624
rect 67177 3621 67189 3624
rect 67223 3621 67235 3655
rect 67177 3615 67235 3621
rect 67358 3612 67364 3664
rect 67416 3652 67422 3664
rect 67913 3655 67971 3661
rect 67913 3652 67925 3655
rect 67416 3624 67925 3652
rect 67416 3612 67422 3624
rect 67913 3621 67925 3624
rect 67959 3621 67971 3655
rect 67913 3615 67971 3621
rect 58989 3587 59047 3593
rect 58989 3584 59001 3587
rect 58860 3556 59001 3584
rect 58860 3544 58866 3556
rect 58989 3553 59001 3556
rect 59035 3553 59047 3587
rect 58989 3547 59047 3553
rect 59449 3587 59507 3593
rect 59449 3553 59461 3587
rect 59495 3584 59507 3587
rect 59998 3584 60004 3596
rect 59495 3556 60004 3584
rect 59495 3553 59507 3556
rect 59449 3547 59507 3553
rect 49200 3488 50384 3516
rect 49200 3476 49206 3488
rect 46566 3448 46572 3460
rect 43956 3420 46336 3448
rect 46527 3420 46572 3448
rect 43956 3408 43962 3420
rect 46566 3408 46572 3420
rect 46624 3408 46630 3460
rect 47486 3448 47492 3460
rect 47447 3420 47492 3448
rect 47486 3408 47492 3420
rect 47544 3408 47550 3460
rect 47670 3408 47676 3460
rect 47728 3448 47734 3460
rect 47728 3420 50292 3448
rect 47728 3408 47734 3420
rect 39908 3352 40908 3380
rect 39908 3340 39914 3352
rect 41322 3340 41328 3392
rect 41380 3380 41386 3392
rect 42702 3380 42708 3392
rect 41380 3352 42708 3380
rect 41380 3340 41386 3352
rect 42702 3340 42708 3352
rect 42760 3340 42766 3392
rect 42794 3340 42800 3392
rect 42852 3380 42858 3392
rect 44269 3383 44327 3389
rect 44269 3380 44281 3383
rect 42852 3352 44281 3380
rect 42852 3340 42858 3352
rect 44269 3349 44281 3352
rect 44315 3349 44327 3383
rect 44269 3343 44327 3349
rect 45738 3340 45744 3392
rect 45796 3380 45802 3392
rect 50062 3380 50068 3392
rect 45796 3352 50068 3380
rect 45796 3340 45802 3352
rect 50062 3340 50068 3352
rect 50120 3340 50126 3392
rect 50264 3380 50292 3420
rect 50338 3408 50344 3460
rect 50396 3448 50402 3460
rect 51276 3448 51304 3544
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 52270 3516 52276 3528
rect 51408 3488 52276 3516
rect 51408 3476 51414 3488
rect 52270 3476 52276 3488
rect 52328 3476 52334 3528
rect 53282 3476 53288 3528
rect 53340 3516 53346 3528
rect 54754 3516 54760 3528
rect 53340 3488 54760 3516
rect 53340 3476 53346 3488
rect 54754 3476 54760 3488
rect 54812 3476 54818 3528
rect 57790 3476 57796 3528
rect 57848 3516 57854 3528
rect 59464 3516 59492 3547
rect 59998 3544 60004 3556
rect 60056 3544 60062 3596
rect 60090 3544 60096 3596
rect 60148 3584 60154 3596
rect 60277 3587 60335 3593
rect 60277 3584 60289 3587
rect 60148 3556 60289 3584
rect 60148 3544 60154 3556
rect 60277 3553 60289 3556
rect 60323 3584 60335 3587
rect 60550 3584 60556 3596
rect 60323 3556 60556 3584
rect 60323 3553 60335 3556
rect 60277 3547 60335 3553
rect 60550 3544 60556 3556
rect 60608 3544 60614 3596
rect 60918 3544 60924 3596
rect 60976 3584 60982 3596
rect 61764 3584 61792 3612
rect 61933 3587 61991 3593
rect 61933 3584 61945 3587
rect 60976 3556 61945 3584
rect 60976 3544 60982 3556
rect 61933 3553 61945 3556
rect 61979 3553 61991 3587
rect 61933 3547 61991 3553
rect 62298 3544 62304 3596
rect 62356 3584 62362 3596
rect 62393 3587 62451 3593
rect 62393 3584 62405 3587
rect 62356 3556 62405 3584
rect 62356 3544 62362 3556
rect 62393 3553 62405 3556
rect 62439 3553 62451 3587
rect 62393 3547 62451 3553
rect 62666 3544 62672 3596
rect 62724 3584 62730 3596
rect 63037 3587 63095 3593
rect 63037 3584 63049 3587
rect 62724 3556 63049 3584
rect 62724 3544 62730 3556
rect 63037 3553 63049 3556
rect 63083 3584 63095 3587
rect 63218 3584 63224 3596
rect 63083 3556 63224 3584
rect 63083 3553 63095 3556
rect 63037 3547 63095 3553
rect 63218 3544 63224 3556
rect 63276 3544 63282 3596
rect 66073 3587 66131 3593
rect 66073 3553 66085 3587
rect 66119 3584 66131 3587
rect 66119 3556 67864 3584
rect 66119 3553 66131 3556
rect 66073 3547 66131 3553
rect 57848 3488 59492 3516
rect 57848 3476 57854 3488
rect 61746 3476 61752 3528
rect 61804 3516 61810 3528
rect 62316 3516 62344 3544
rect 61804 3488 62344 3516
rect 61804 3476 61810 3488
rect 66806 3476 66812 3528
rect 66864 3516 66870 3528
rect 67266 3516 67272 3528
rect 66864 3488 67272 3516
rect 66864 3476 66870 3488
rect 67266 3476 67272 3488
rect 67324 3476 67330 3528
rect 67836 3516 67864 3556
rect 68278 3516 68284 3528
rect 67836 3488 68284 3516
rect 68278 3476 68284 3488
rect 68336 3476 68342 3528
rect 50396 3420 51304 3448
rect 50396 3408 50402 3420
rect 51442 3408 51448 3460
rect 51500 3448 51506 3460
rect 51718 3448 51724 3460
rect 51500 3420 51724 3448
rect 51500 3408 51506 3420
rect 51718 3408 51724 3420
rect 51776 3408 51782 3460
rect 52546 3448 52552 3460
rect 52507 3420 52552 3448
rect 52546 3408 52552 3420
rect 52604 3408 52610 3460
rect 53374 3448 53380 3460
rect 53335 3420 53380 3448
rect 53374 3408 53380 3420
rect 53432 3408 53438 3460
rect 54110 3408 54116 3460
rect 54168 3448 54174 3460
rect 54297 3451 54355 3457
rect 54297 3448 54309 3451
rect 54168 3420 54309 3448
rect 54168 3408 54174 3420
rect 54297 3417 54309 3420
rect 54343 3417 54355 3451
rect 55122 3448 55128 3460
rect 55083 3420 55128 3448
rect 54297 3411 54355 3417
rect 55122 3408 55128 3420
rect 55180 3408 55186 3460
rect 56410 3408 56416 3460
rect 56468 3448 56474 3460
rect 56505 3451 56563 3457
rect 56505 3448 56517 3451
rect 56468 3420 56517 3448
rect 56468 3408 56474 3420
rect 56505 3417 56517 3420
rect 56551 3417 56563 3451
rect 57238 3448 57244 3460
rect 57199 3420 57244 3448
rect 56505 3411 56563 3417
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 64046 3448 64052 3460
rect 64007 3420 64052 3448
rect 64046 3408 64052 3420
rect 64104 3408 64110 3460
rect 64874 3448 64880 3460
rect 64835 3420 64880 3448
rect 64874 3408 64880 3420
rect 64932 3408 64938 3460
rect 65794 3408 65800 3460
rect 65852 3448 65858 3460
rect 66346 3448 66352 3460
rect 65852 3420 66352 3448
rect 65852 3408 65858 3420
rect 66346 3408 66352 3420
rect 66404 3408 66410 3460
rect 66990 3408 66996 3460
rect 67048 3448 67054 3460
rect 67729 3451 67787 3457
rect 67729 3448 67741 3451
rect 67048 3420 67741 3448
rect 67048 3408 67054 3420
rect 67729 3417 67741 3420
rect 67775 3417 67787 3451
rect 67729 3411 67787 3417
rect 50522 3380 50528 3392
rect 50264 3352 50528 3380
rect 50522 3340 50528 3352
rect 50580 3340 50586 3392
rect 50798 3340 50804 3392
rect 50856 3380 50862 3392
rect 51074 3380 51080 3392
rect 50856 3352 51080 3380
rect 50856 3340 50862 3352
rect 51074 3340 51080 3352
rect 51132 3340 51138 3392
rect 51166 3340 51172 3392
rect 51224 3380 51230 3392
rect 51810 3380 51816 3392
rect 51224 3352 51816 3380
rect 51224 3340 51230 3352
rect 51810 3340 51816 3352
rect 51868 3340 51874 3392
rect 52362 3340 52368 3392
rect 52420 3380 52426 3392
rect 53190 3380 53196 3392
rect 52420 3352 53196 3380
rect 52420 3340 52426 3352
rect 53190 3340 53196 3352
rect 53248 3380 53254 3392
rect 53742 3380 53748 3392
rect 53248 3352 53748 3380
rect 53248 3340 53254 3352
rect 53742 3340 53748 3352
rect 53800 3340 53806 3392
rect 58526 3340 58532 3392
rect 58584 3380 58590 3392
rect 60737 3383 60795 3389
rect 60737 3380 60749 3383
rect 58584 3352 60749 3380
rect 58584 3340 58590 3352
rect 60737 3349 60749 3352
rect 60783 3349 60795 3383
rect 60737 3343 60795 3349
rect 66162 3340 66168 3392
rect 66220 3380 66226 3392
rect 67085 3383 67143 3389
rect 67085 3380 67097 3383
rect 66220 3352 67097 3380
rect 66220 3340 66226 3352
rect 67085 3349 67097 3352
rect 67131 3349 67143 3383
rect 67085 3343 67143 3349
rect 27479 3284 35112 3312
rect 27479 3281 27491 3284
rect 27433 3275 27491 3281
rect 35526 3272 35532 3324
rect 35584 3312 35590 3324
rect 37369 3315 37427 3321
rect 37369 3312 37381 3315
rect 35584 3284 37381 3312
rect 35584 3272 35590 3284
rect 37369 3281 37381 3284
rect 37415 3281 37427 3315
rect 37369 3275 37427 3281
rect 37628 3290 68816 3312
rect 1104 3216 18952 3238
rect 19058 3204 19064 3256
rect 19116 3244 19122 3256
rect 21634 3244 21640 3256
rect 19116 3216 21640 3244
rect 19116 3204 19122 3216
rect 21634 3204 21640 3216
rect 21692 3204 21698 3256
rect 21729 3247 21787 3253
rect 21729 3213 21741 3247
rect 21775 3244 21787 3247
rect 22097 3247 22155 3253
rect 22097 3244 22109 3247
rect 21775 3216 22109 3244
rect 21775 3213 21787 3216
rect 21729 3207 21787 3213
rect 22097 3213 22109 3216
rect 22143 3213 22155 3247
rect 22097 3207 22155 3213
rect 31573 3247 31631 3253
rect 31573 3213 31585 3247
rect 31619 3244 31631 3247
rect 33870 3244 33876 3256
rect 31619 3216 33876 3244
rect 31619 3213 31631 3216
rect 31573 3207 31631 3213
rect 33870 3204 33876 3216
rect 33928 3204 33934 3256
rect 33965 3247 34023 3253
rect 33965 3213 33977 3247
rect 34011 3244 34023 3247
rect 35342 3244 35348 3256
rect 34011 3216 35348 3244
rect 34011 3213 34023 3216
rect 33965 3207 34023 3213
rect 35342 3204 35348 3216
rect 35400 3204 35406 3256
rect 35434 3204 35440 3256
rect 35492 3244 35498 3256
rect 37090 3244 37096 3256
rect 35492 3216 37096 3244
rect 35492 3204 35498 3216
rect 37090 3204 37096 3216
rect 37148 3204 37154 3256
rect 37628 3238 44246 3290
rect 44298 3238 44310 3290
rect 44362 3238 44374 3290
rect 44426 3238 44438 3290
rect 44490 3238 54246 3290
rect 54298 3238 54310 3290
rect 54362 3238 54374 3290
rect 54426 3238 54438 3290
rect 54490 3238 64246 3290
rect 64298 3238 64310 3290
rect 64362 3238 64374 3290
rect 64426 3238 64438 3290
rect 64490 3238 68816 3290
rect 37628 3216 68816 3238
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 2866 3176 2872 3188
rect 2547 3148 2872 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 3384 3148 5641 3176
rect 3384 3136 3390 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 5629 3139 5687 3145
rect 10686 3136 10692 3188
rect 10744 3136 10750 3188
rect 13538 3176 13544 3188
rect 12176 3148 13544 3176
rect 2774 3068 2780 3120
rect 2832 3108 2838 3120
rect 4801 3111 4859 3117
rect 4801 3108 4813 3111
rect 2832 3080 4813 3108
rect 2832 3068 2838 3080
rect 4801 3077 4813 3080
rect 4847 3077 4859 3111
rect 4801 3071 4859 3077
rect 8110 3068 8116 3120
rect 8168 3108 8174 3120
rect 10704 3108 10732 3136
rect 8168 3080 10088 3108
rect 10704 3080 11468 3108
rect 8168 3068 8174 3080
rect 2222 3000 2228 3052
rect 2280 3040 2286 3052
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 2280 3012 4077 3040
rect 2280 3000 2286 3012
rect 4065 3009 4077 3012
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4706 3040 4712 3052
rect 4212 3012 4712 3040
rect 4212 3000 4218 3012
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5810 3040 5816 3052
rect 5000 3012 5816 3040
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 1728 2944 3341 2972
rect 1728 2932 1734 2944
rect 3329 2941 3341 2944
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 3694 2972 3700 2984
rect 3559 2944 3700 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 5000 2981 5028 3012
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8536 3012 8800 3040
rect 8536 3000 8542 3012
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2941 5043 2975
rect 4985 2935 5043 2941
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 5592 2944 6837 2972
rect 5592 2932 5598 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7190 2972 7196 2984
rect 7055 2944 7196 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8110 2972 8116 2984
rect 8067 2944 8116 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8662 2972 8668 2984
rect 8623 2944 8668 2972
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 1949 2907 2007 2913
rect 1949 2873 1961 2907
rect 1995 2904 2007 2907
rect 2314 2904 2320 2916
rect 1995 2876 2320 2904
rect 1995 2873 2007 2876
rect 1949 2867 2007 2873
rect 2314 2864 2320 2876
rect 2372 2864 2378 2916
rect 2501 2907 2559 2913
rect 2501 2873 2513 2907
rect 2547 2904 2559 2907
rect 2777 2907 2835 2913
rect 2777 2904 2789 2907
rect 2547 2876 2789 2904
rect 2547 2873 2559 2876
rect 2501 2867 2559 2873
rect 2777 2873 2789 2876
rect 2823 2873 2835 2907
rect 4062 2904 4068 2916
rect 2777 2867 2835 2873
rect 3712 2876 4068 2904
rect 3712 2848 3740 2876
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 4249 2907 4307 2913
rect 4249 2873 4261 2907
rect 4295 2904 4307 2907
rect 5258 2904 5264 2916
rect 4295 2876 5264 2904
rect 4295 2873 4307 2876
rect 4249 2867 4307 2873
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 5721 2907 5779 2913
rect 5721 2873 5733 2907
rect 5767 2904 5779 2907
rect 6546 2904 6552 2916
rect 5767 2876 6552 2904
rect 5767 2873 5779 2876
rect 5721 2867 5779 2873
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 8478 2904 8484 2916
rect 8439 2876 8484 2904
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 106 2796 112 2848
rect 164 2836 170 2848
rect 1578 2836 1584 2848
rect 164 2808 1584 2836
rect 164 2796 170 2808
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 2866 2836 2872 2848
rect 2731 2808 2872 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 3694 2796 3700 2848
rect 3752 2796 3758 2848
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 7006 2836 7012 2848
rect 5868 2808 7012 2836
rect 5868 2796 5874 2808
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 8772 2836 8800 3012
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 8904 2944 9965 2972
rect 8904 2932 8910 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 10060 2972 10088 3080
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10192 3012 10701 3040
rect 10192 3000 10198 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 11440 3040 11468 3080
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 12176 3108 12204 3148
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 19153 3179 19211 3185
rect 19153 3176 19165 3179
rect 14108 3148 19165 3176
rect 14108 3108 14136 3148
rect 19153 3145 19165 3148
rect 19199 3145 19211 3179
rect 19153 3139 19211 3145
rect 20717 3179 20775 3185
rect 20717 3145 20729 3179
rect 20763 3176 20775 3179
rect 23658 3176 23664 3188
rect 20763 3148 23664 3176
rect 20763 3145 20775 3148
rect 20717 3139 20775 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 24486 3136 24492 3188
rect 24544 3176 24550 3188
rect 26329 3179 26387 3185
rect 26329 3176 26341 3179
rect 24544 3148 26341 3176
rect 24544 3136 24550 3148
rect 26329 3145 26341 3148
rect 26375 3145 26387 3179
rect 26329 3139 26387 3145
rect 29457 3179 29515 3185
rect 29457 3145 29469 3179
rect 29503 3176 29515 3179
rect 34698 3176 34704 3188
rect 29503 3148 34008 3176
rect 29503 3145 29515 3148
rect 29457 3139 29515 3145
rect 11572 3080 12204 3108
rect 12268 3080 14136 3108
rect 14185 3111 14243 3117
rect 11572 3068 11578 3080
rect 12268 3040 12296 3080
rect 14185 3077 14197 3111
rect 14231 3108 14243 3111
rect 16393 3111 16451 3117
rect 14231 3080 16344 3108
rect 14231 3077 14243 3080
rect 14185 3071 14243 3077
rect 11440 3012 12296 3040
rect 16316 3040 16344 3080
rect 16393 3077 16405 3111
rect 16439 3108 16451 3111
rect 19061 3111 19119 3117
rect 19061 3108 19073 3111
rect 16439 3080 19073 3108
rect 16439 3077 16451 3080
rect 16393 3071 16451 3077
rect 19061 3077 19073 3080
rect 19107 3077 19119 3111
rect 19061 3071 19119 3077
rect 21082 3068 21088 3120
rect 21140 3108 21146 3120
rect 22465 3111 22523 3117
rect 22465 3108 22477 3111
rect 21140 3080 22477 3108
rect 21140 3068 21146 3080
rect 22465 3077 22477 3080
rect 22511 3077 22523 3111
rect 22465 3071 22523 3077
rect 24394 3068 24400 3120
rect 24452 3108 24458 3120
rect 26053 3111 26111 3117
rect 26053 3108 26065 3111
rect 24452 3080 26065 3108
rect 24452 3068 24458 3080
rect 26053 3077 26065 3080
rect 26099 3077 26111 3111
rect 26053 3071 26111 3077
rect 29549 3111 29607 3117
rect 29549 3077 29561 3111
rect 29595 3108 29607 3111
rect 33873 3111 33931 3117
rect 33873 3108 33885 3111
rect 29595 3080 33885 3108
rect 29595 3077 29607 3080
rect 29549 3071 29607 3077
rect 33873 3077 33885 3080
rect 33919 3077 33931 3111
rect 33980 3108 34008 3148
rect 34624 3148 34704 3176
rect 34624 3108 34652 3148
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 34885 3179 34943 3185
rect 34885 3145 34897 3179
rect 34931 3176 34943 3179
rect 35621 3179 35679 3185
rect 35621 3176 35633 3179
rect 34931 3148 35633 3176
rect 34931 3145 34943 3148
rect 34885 3139 34943 3145
rect 35621 3145 35633 3148
rect 35667 3145 35679 3179
rect 35621 3139 35679 3145
rect 35713 3179 35771 3185
rect 35713 3145 35725 3179
rect 35759 3176 35771 3179
rect 39117 3179 39175 3185
rect 39117 3176 39129 3179
rect 35759 3148 39129 3176
rect 35759 3145 35771 3148
rect 35713 3139 35771 3145
rect 39117 3145 39129 3148
rect 39163 3145 39175 3179
rect 40034 3176 40040 3188
rect 39117 3139 39175 3145
rect 39224 3148 40040 3176
rect 33980 3080 34652 3108
rect 34716 3080 34928 3108
rect 33873 3071 33931 3077
rect 18506 3040 18512 3052
rect 16316 3012 18512 3040
rect 10689 3003 10747 3009
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 24946 3040 24952 3052
rect 18656 3012 24952 3040
rect 18656 3000 18662 3012
rect 24946 3000 24952 3012
rect 25004 3000 25010 3052
rect 26605 3043 26663 3049
rect 26605 3009 26617 3043
rect 26651 3040 26663 3043
rect 34716 3040 34744 3080
rect 26651 3012 34744 3040
rect 34900 3040 34928 3080
rect 35066 3068 35072 3120
rect 35124 3108 35130 3120
rect 39224 3108 39252 3148
rect 40034 3136 40040 3148
rect 40092 3136 40098 3188
rect 40310 3136 40316 3188
rect 40368 3176 40374 3188
rect 41414 3176 41420 3188
rect 40368 3148 41420 3176
rect 40368 3136 40374 3148
rect 41414 3136 41420 3148
rect 41472 3136 41478 3188
rect 41874 3136 41880 3188
rect 41932 3176 41938 3188
rect 44177 3179 44235 3185
rect 44177 3176 44189 3179
rect 41932 3148 44189 3176
rect 41932 3136 41938 3148
rect 44177 3145 44189 3148
rect 44223 3145 44235 3179
rect 44177 3139 44235 3145
rect 45646 3136 45652 3188
rect 45704 3176 45710 3188
rect 47394 3176 47400 3188
rect 45704 3148 47400 3176
rect 45704 3136 45710 3148
rect 47394 3136 47400 3148
rect 47452 3136 47458 3188
rect 48286 3148 48636 3176
rect 39758 3108 39764 3120
rect 35124 3080 39252 3108
rect 39719 3080 39764 3108
rect 35124 3068 35130 3080
rect 39758 3068 39764 3080
rect 39816 3068 39822 3120
rect 41233 3111 41291 3117
rect 41233 3108 41245 3111
rect 40236 3080 41245 3108
rect 38289 3043 38347 3049
rect 38289 3040 38301 3043
rect 34900 3012 38301 3040
rect 26651 3009 26663 3012
rect 26605 3003 26663 3009
rect 38289 3009 38301 3012
rect 38335 3009 38347 3043
rect 38289 3003 38347 3009
rect 39114 3000 39120 3052
rect 39172 3040 39178 3052
rect 40126 3040 40132 3052
rect 39172 3012 40132 3040
rect 39172 3000 39178 3012
rect 40126 3000 40132 3012
rect 40184 3000 40190 3052
rect 10502 2972 10508 2984
rect 10060 2944 10508 2972
rect 9953 2935 10011 2941
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 10594 2932 10600 2984
rect 10652 2972 10658 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 10652 2944 12081 2972
rect 10652 2932 10658 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12860 2944 13001 2972
rect 12860 2932 12866 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 13998 2972 14004 2984
rect 13959 2944 14004 2972
rect 12989 2935 13047 2941
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 15010 2972 15016 2984
rect 14783 2944 15016 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 15565 2975 15623 2981
rect 15565 2941 15577 2975
rect 15611 2972 15623 2975
rect 15930 2972 15936 2984
rect 15611 2944 15936 2972
rect 15611 2941 15623 2944
rect 15565 2935 15623 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16206 2972 16212 2984
rect 16167 2944 16212 2972
rect 16206 2932 16212 2944
rect 16264 2932 16270 2984
rect 16298 2932 16304 2984
rect 16356 2972 16362 2984
rect 17494 2972 17500 2984
rect 16356 2944 16528 2972
rect 17455 2944 17500 2972
rect 16356 2932 16362 2944
rect 8938 2864 8944 2916
rect 8996 2904 9002 2916
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 8996 2876 9229 2904
rect 8996 2864 9002 2876
rect 9217 2873 9229 2876
rect 9263 2873 9275 2907
rect 9217 2867 9275 2873
rect 9401 2907 9459 2913
rect 9401 2873 9413 2907
rect 9447 2873 9459 2907
rect 9401 2867 9459 2873
rect 9416 2836 9444 2867
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 10137 2907 10195 2913
rect 10137 2904 10149 2907
rect 9824 2876 10149 2904
rect 9824 2864 9830 2876
rect 10137 2873 10149 2876
rect 10183 2873 10195 2907
rect 10870 2904 10876 2916
rect 10831 2876 10876 2904
rect 10137 2867 10195 2873
rect 10870 2864 10876 2876
rect 10928 2864 10934 2916
rect 11790 2864 11796 2916
rect 11848 2904 11854 2916
rect 12253 2907 12311 2913
rect 12253 2904 12265 2907
rect 11848 2876 12265 2904
rect 11848 2864 11854 2876
rect 12253 2873 12265 2876
rect 12299 2873 12311 2907
rect 12253 2867 12311 2873
rect 14921 2907 14979 2913
rect 14921 2873 14933 2907
rect 14967 2904 14979 2907
rect 16390 2904 16396 2916
rect 14967 2876 16396 2904
rect 14967 2873 14979 2876
rect 14921 2867 14979 2873
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 16500 2904 16528 2944
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 22554 2972 22560 2984
rect 18012 2944 22560 2972
rect 18012 2932 18018 2944
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 25317 2975 25375 2981
rect 25317 2941 25329 2975
rect 25363 2972 25375 2975
rect 31846 2972 31852 2984
rect 25363 2944 31852 2972
rect 25363 2941 25375 2944
rect 25317 2935 25375 2941
rect 31846 2932 31852 2944
rect 31904 2932 31910 2984
rect 32950 2972 32956 2984
rect 32140 2944 32956 2972
rect 17862 2904 17868 2916
rect 16500 2876 17868 2904
rect 17862 2864 17868 2876
rect 17920 2864 17926 2916
rect 18049 2907 18107 2913
rect 18049 2873 18061 2907
rect 18095 2873 18107 2907
rect 18049 2867 18107 2873
rect 18233 2907 18291 2913
rect 18233 2873 18245 2907
rect 18279 2904 18291 2907
rect 20254 2904 20260 2916
rect 18279 2876 20260 2904
rect 18279 2873 18291 2876
rect 18233 2867 18291 2873
rect 8772 2808 9444 2836
rect 12802 2796 12808 2848
rect 12860 2836 12866 2848
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12860 2808 12909 2836
rect 12860 2796 12866 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 15470 2836 15476 2848
rect 15431 2808 15476 2836
rect 12897 2799 12955 2805
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 17494 2836 17500 2848
rect 16172 2808 17500 2836
rect 16172 2796 16178 2808
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 18064 2836 18092 2867
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 20346 2864 20352 2916
rect 20404 2904 20410 2916
rect 21729 2907 21787 2913
rect 21729 2904 21741 2907
rect 20404 2876 21741 2904
rect 20404 2864 20410 2876
rect 21729 2873 21741 2876
rect 21775 2873 21787 2907
rect 21729 2867 21787 2873
rect 23566 2864 23572 2916
rect 23624 2904 23630 2916
rect 26789 2907 26847 2913
rect 26789 2904 26801 2907
rect 23624 2876 26801 2904
rect 23624 2864 23630 2876
rect 26789 2873 26801 2876
rect 26835 2873 26847 2907
rect 26789 2867 26847 2873
rect 31297 2907 31355 2913
rect 31297 2873 31309 2907
rect 31343 2904 31355 2907
rect 31662 2904 31668 2916
rect 31343 2876 31668 2904
rect 31343 2873 31355 2876
rect 31297 2867 31355 2873
rect 31662 2864 31668 2876
rect 31720 2864 31726 2916
rect 32140 2904 32168 2944
rect 32950 2932 32956 2944
rect 33008 2932 33014 2984
rect 37458 2932 37464 2984
rect 37516 2972 37522 2984
rect 38473 2975 38531 2981
rect 38473 2972 38485 2975
rect 37516 2944 38485 2972
rect 37516 2932 37522 2944
rect 38473 2941 38485 2944
rect 38519 2941 38531 2975
rect 39206 2972 39212 2984
rect 39167 2944 39212 2972
rect 38473 2935 38531 2941
rect 39206 2932 39212 2944
rect 39264 2932 39270 2984
rect 39942 2972 39948 2984
rect 39903 2944 39948 2972
rect 39942 2932 39948 2944
rect 40000 2932 40006 2984
rect 32582 2904 32588 2916
rect 31864 2876 32168 2904
rect 32232 2876 32588 2904
rect 18690 2836 18696 2848
rect 18064 2808 18696 2836
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 19794 2836 19800 2848
rect 18984 2808 19800 2836
rect 1104 2746 18952 2768
rect 1104 2694 9246 2746
rect 9298 2694 9310 2746
rect 9362 2694 9374 2746
rect 9426 2694 9438 2746
rect 9490 2694 18952 2746
rect 1104 2672 18952 2694
rect 15933 2635 15991 2641
rect 15933 2601 15945 2635
rect 15979 2632 15991 2635
rect 16298 2632 16304 2644
rect 15979 2604 16304 2632
rect 15979 2601 15991 2604
rect 15933 2595 15991 2601
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 16577 2635 16635 2641
rect 16577 2601 16589 2635
rect 16623 2632 16635 2635
rect 18984 2632 19012 2808
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 21174 2796 21180 2848
rect 21232 2836 21238 2848
rect 23382 2836 23388 2848
rect 21232 2808 23152 2836
rect 23343 2808 23388 2836
rect 21232 2796 21238 2808
rect 23124 2712 23152 2808
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 24118 2796 24124 2848
rect 24176 2836 24182 2848
rect 25593 2839 25651 2845
rect 25593 2836 25605 2839
rect 24176 2808 25605 2836
rect 24176 2796 24182 2808
rect 25593 2805 25605 2808
rect 25639 2805 25651 2839
rect 25593 2799 25651 2805
rect 27617 2839 27675 2845
rect 27617 2805 27629 2839
rect 27663 2836 27675 2839
rect 31864 2836 31892 2876
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 27663 2808 31892 2836
rect 31956 2808 32137 2836
rect 27663 2805 27675 2808
rect 27617 2799 27675 2805
rect 22557 2703 22615 2709
rect 22557 2669 22569 2703
rect 22603 2700 22615 2703
rect 22738 2700 22744 2712
rect 22603 2672 22744 2700
rect 22603 2669 22615 2672
rect 22557 2663 22615 2669
rect 22738 2660 22744 2672
rect 22796 2660 22802 2712
rect 23106 2660 23112 2712
rect 23164 2660 23170 2712
rect 23382 2700 23388 2712
rect 23343 2672 23388 2700
rect 23382 2660 23388 2672
rect 23440 2660 23446 2712
rect 31846 2660 31852 2712
rect 31904 2700 31910 2712
rect 31956 2700 31984 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 32030 2728 32036 2780
rect 32088 2728 32094 2780
rect 31904 2672 31984 2700
rect 31904 2660 31910 2672
rect 16623 2604 19012 2632
rect 19153 2635 19211 2641
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 19153 2601 19165 2635
rect 19199 2632 19211 2635
rect 24026 2632 24032 2644
rect 19199 2604 24032 2632
rect 19199 2601 19211 2604
rect 19153 2595 19211 2601
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 32048 2576 32076 2728
rect 1118 2524 1124 2576
rect 1176 2564 1182 2576
rect 4985 2567 5043 2573
rect 4985 2564 4997 2567
rect 1176 2536 4997 2564
rect 1176 2524 1182 2536
rect 4985 2533 4997 2536
rect 5031 2533 5043 2567
rect 4985 2527 5043 2533
rect 5169 2567 5227 2573
rect 5169 2533 5181 2567
rect 5215 2564 5227 2567
rect 5350 2564 5356 2576
rect 5215 2536 5356 2564
rect 5215 2533 5227 2536
rect 5169 2527 5227 2533
rect 5350 2524 5356 2536
rect 5408 2524 5414 2576
rect 5902 2564 5908 2576
rect 5863 2536 5908 2564
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 7098 2564 7104 2576
rect 7059 2536 7104 2564
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 7834 2564 7840 2576
rect 7795 2536 7840 2564
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8570 2564 8576 2576
rect 8531 2536 8576 2564
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 9766 2564 9772 2576
rect 9727 2536 9772 2564
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 10686 2564 10692 2576
rect 10551 2536 10692 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 10686 2524 10692 2536
rect 10744 2524 10750 2576
rect 12342 2564 12348 2576
rect 12303 2536 12348 2564
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 13078 2564 13084 2576
rect 13039 2536 13084 2564
rect 13078 2524 13084 2536
rect 13136 2524 13142 2576
rect 13814 2564 13820 2576
rect 13775 2536 13820 2564
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 15289 2567 15347 2573
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 15378 2564 15384 2576
rect 15335 2536 15384 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 15378 2524 15384 2536
rect 15436 2524 15442 2576
rect 16485 2567 16543 2573
rect 16485 2533 16497 2567
rect 16531 2564 16543 2567
rect 16758 2564 16764 2576
rect 16531 2536 16764 2564
rect 16531 2533 16543 2536
rect 16485 2527 16543 2533
rect 16758 2524 16764 2536
rect 16816 2524 16822 2576
rect 18049 2567 18107 2573
rect 18049 2533 18061 2567
rect 18095 2564 18107 2567
rect 18414 2564 18420 2576
rect 18095 2536 18420 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 18414 2524 18420 2536
rect 18472 2524 18478 2576
rect 18782 2524 18788 2576
rect 18840 2564 18846 2576
rect 19245 2567 19303 2573
rect 19245 2564 19257 2567
rect 18840 2536 19257 2564
rect 18840 2524 18846 2536
rect 19245 2533 19257 2536
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 32030 2524 32036 2576
rect 32088 2524 32094 2576
rect 32122 2524 32128 2576
rect 32180 2564 32186 2576
rect 32232 2564 32260 2876
rect 32582 2864 32588 2876
rect 32640 2864 32646 2916
rect 35713 2907 35771 2913
rect 35713 2873 35725 2907
rect 35759 2904 35771 2907
rect 40236 2904 40264 3080
rect 41233 3077 41245 3080
rect 41279 3077 41291 3111
rect 41233 3071 41291 3077
rect 42886 3068 42892 3120
rect 42944 3108 42950 3120
rect 44910 3108 44916 3120
rect 42944 3080 44916 3108
rect 42944 3068 42950 3080
rect 44910 3068 44916 3080
rect 44968 3068 44974 3120
rect 45278 3068 45284 3120
rect 45336 3108 45342 3120
rect 45336 3080 47900 3108
rect 45336 3068 45342 3080
rect 40494 3040 40500 3052
rect 40455 3012 40500 3040
rect 40494 3000 40500 3012
rect 40552 3000 40558 3052
rect 40770 3000 40776 3052
rect 40828 3040 40834 3052
rect 43349 3043 43407 3049
rect 43349 3040 43361 3043
rect 40828 3012 43361 3040
rect 40828 3000 40834 3012
rect 43349 3009 43361 3012
rect 43395 3009 43407 3043
rect 43349 3003 43407 3009
rect 44082 3000 44088 3052
rect 44140 3040 44146 3052
rect 45557 3043 45615 3049
rect 45557 3040 45569 3043
rect 44140 3012 45569 3040
rect 44140 3000 44146 3012
rect 45557 3009 45569 3012
rect 45603 3009 45615 3043
rect 45557 3003 45615 3009
rect 46106 3000 46112 3052
rect 46164 3040 46170 3052
rect 47029 3043 47087 3049
rect 47029 3040 47041 3043
rect 46164 3012 47041 3040
rect 46164 3000 46170 3012
rect 47029 3009 47041 3012
rect 47075 3009 47087 3043
rect 47762 3040 47768 3052
rect 47029 3003 47087 3009
rect 47228 3012 47768 3040
rect 40678 2972 40684 2984
rect 40639 2944 40684 2972
rect 40678 2932 40684 2944
rect 40736 2932 40742 2984
rect 41414 2972 41420 2984
rect 41375 2944 41420 2972
rect 41414 2932 41420 2944
rect 41472 2932 41478 2984
rect 41966 2972 41972 2984
rect 41927 2944 41972 2972
rect 41966 2932 41972 2944
rect 42024 2932 42030 2984
rect 43162 2972 43168 2984
rect 42076 2944 43168 2972
rect 35759 2876 40264 2904
rect 35759 2873 35771 2876
rect 35713 2867 35771 2873
rect 40494 2864 40500 2916
rect 40552 2904 40558 2916
rect 42076 2904 42104 2944
rect 43162 2932 43168 2944
rect 43220 2932 43226 2984
rect 43533 2975 43591 2981
rect 43533 2941 43545 2975
rect 43579 2972 43591 2975
rect 43714 2972 43720 2984
rect 43579 2944 43720 2972
rect 43579 2941 43591 2944
rect 43533 2935 43591 2941
rect 43714 2932 43720 2944
rect 43772 2932 43778 2984
rect 44269 2975 44327 2981
rect 44269 2941 44281 2975
rect 44315 2972 44327 2975
rect 44634 2972 44640 2984
rect 44315 2944 44640 2972
rect 44315 2941 44327 2944
rect 44269 2935 44327 2941
rect 44634 2932 44640 2944
rect 44692 2932 44698 2984
rect 46474 2932 46480 2984
rect 46532 2972 46538 2984
rect 47228 2981 47256 3012
rect 47762 3000 47768 3012
rect 47820 3000 47826 3052
rect 47213 2975 47271 2981
rect 46532 2944 46577 2972
rect 46532 2932 46538 2944
rect 47213 2941 47225 2975
rect 47259 2941 47271 2975
rect 47872 2972 47900 3080
rect 48286 3052 48314 3148
rect 48222 3000 48228 3052
rect 48280 3012 48314 3052
rect 48280 3000 48286 3012
rect 48498 3000 48504 3052
rect 48556 3000 48562 3052
rect 48516 2972 48544 3000
rect 47872 2944 48544 2972
rect 48608 2972 48636 3148
rect 62850 3136 62856 3188
rect 62908 3176 62914 3188
rect 62908 3148 65932 3176
rect 62908 3136 62914 3148
rect 48774 3068 48780 3120
rect 48832 3068 48838 3120
rect 49786 3108 49792 3120
rect 48884 3080 49792 3108
rect 48682 2972 48688 2984
rect 48608 2944 48688 2972
rect 47213 2935 47271 2941
rect 48682 2932 48688 2944
rect 48740 2932 48746 2984
rect 48792 2981 48820 3068
rect 48777 2975 48835 2981
rect 48777 2941 48789 2975
rect 48823 2941 48835 2975
rect 48777 2935 48835 2941
rect 40552 2876 42104 2904
rect 42153 2907 42211 2913
rect 40552 2864 40558 2876
rect 42153 2873 42165 2907
rect 42199 2904 42211 2907
rect 42426 2904 42432 2916
rect 42199 2876 42432 2904
rect 42199 2873 42211 2876
rect 42153 2867 42211 2873
rect 42426 2864 42432 2876
rect 42484 2864 42490 2916
rect 44821 2907 44879 2913
rect 44821 2904 44833 2907
rect 43640 2876 44833 2904
rect 32309 2839 32367 2845
rect 32309 2805 32321 2839
rect 32355 2836 32367 2839
rect 32766 2836 32772 2848
rect 32355 2808 32772 2836
rect 32355 2805 32367 2808
rect 32309 2799 32367 2805
rect 32766 2796 32772 2808
rect 32824 2796 32830 2848
rect 32950 2836 32956 2848
rect 32911 2808 32956 2836
rect 32950 2796 32956 2808
rect 33008 2796 33014 2848
rect 35989 2839 36047 2845
rect 35989 2805 36001 2839
rect 36035 2836 36047 2839
rect 40126 2836 40132 2848
rect 36035 2808 40132 2836
rect 36035 2805 36047 2808
rect 35989 2799 36047 2805
rect 40126 2796 40132 2808
rect 40184 2796 40190 2848
rect 41782 2796 41788 2848
rect 41840 2836 41846 2848
rect 42978 2836 42984 2848
rect 41840 2808 42984 2836
rect 41840 2796 41846 2808
rect 42978 2796 42984 2808
rect 43036 2796 43042 2848
rect 43254 2796 43260 2848
rect 43312 2836 43318 2848
rect 43640 2836 43668 2876
rect 44821 2873 44833 2876
rect 44867 2873 44879 2907
rect 45002 2904 45008 2916
rect 44963 2876 45008 2904
rect 44821 2867 44879 2873
rect 45002 2864 45008 2876
rect 45060 2864 45066 2916
rect 45462 2864 45468 2916
rect 45520 2904 45526 2916
rect 45741 2907 45799 2913
rect 45741 2904 45753 2907
rect 45520 2876 45753 2904
rect 45520 2864 45526 2876
rect 45741 2873 45753 2876
rect 45787 2873 45799 2907
rect 45741 2867 45799 2873
rect 47854 2864 47860 2916
rect 47912 2904 47918 2916
rect 48593 2907 48651 2913
rect 48593 2904 48605 2907
rect 47912 2876 48605 2904
rect 47912 2864 47918 2876
rect 48593 2873 48605 2876
rect 48639 2873 48651 2907
rect 48593 2867 48651 2873
rect 43312 2808 43668 2836
rect 43312 2796 43318 2808
rect 44910 2796 44916 2848
rect 44968 2836 44974 2848
rect 46385 2839 46443 2845
rect 46385 2836 46397 2839
rect 44968 2808 46397 2836
rect 44968 2796 44974 2808
rect 46385 2805 46397 2808
rect 46431 2805 46443 2839
rect 46385 2799 46443 2805
rect 47026 2796 47032 2848
rect 47084 2836 47090 2848
rect 48884 2836 48912 3080
rect 49786 3068 49792 3080
rect 49844 3068 49850 3120
rect 50522 3068 50528 3120
rect 50580 3108 50586 3120
rect 54202 3108 54208 3120
rect 50580 3080 54208 3108
rect 50580 3068 50586 3080
rect 54202 3068 54208 3080
rect 54260 3068 54266 3120
rect 62758 3068 62764 3120
rect 62816 3108 62822 3120
rect 65794 3108 65800 3120
rect 62816 3080 65800 3108
rect 62816 3068 62822 3080
rect 65794 3068 65800 3080
rect 65852 3068 65858 3120
rect 65904 3108 65932 3148
rect 66070 3136 66076 3188
rect 66128 3176 66134 3188
rect 67269 3179 67327 3185
rect 67269 3176 67281 3179
rect 66128 3148 67281 3176
rect 66128 3136 66134 3148
rect 67269 3145 67281 3148
rect 67315 3145 67327 3179
rect 69382 3176 69388 3188
rect 67269 3139 67327 3145
rect 67376 3148 69388 3176
rect 67376 3108 67404 3148
rect 69382 3136 69388 3148
rect 69440 3136 69446 3188
rect 68094 3108 68100 3120
rect 65904 3080 67404 3108
rect 68055 3080 68100 3108
rect 68094 3068 68100 3080
rect 68152 3068 68158 3120
rect 50890 3000 50896 3052
rect 50948 3040 50954 3052
rect 51537 3043 51595 3049
rect 51537 3040 51549 3043
rect 50948 3012 51549 3040
rect 50948 3000 50954 3012
rect 51537 3009 51549 3012
rect 51583 3009 51595 3043
rect 51537 3003 51595 3009
rect 51718 3000 51724 3052
rect 51776 3040 51782 3052
rect 52273 3043 52331 3049
rect 52273 3040 52285 3043
rect 51776 3012 52285 3040
rect 51776 3000 51782 3012
rect 52273 3009 52285 3012
rect 52319 3009 52331 3043
rect 52273 3003 52331 3009
rect 53834 3000 53840 3052
rect 53892 3040 53898 3052
rect 54573 3043 54631 3049
rect 54573 3040 54585 3043
rect 53892 3012 54585 3040
rect 53892 3000 53898 3012
rect 54573 3009 54585 3012
rect 54619 3009 54631 3043
rect 54573 3003 54631 3009
rect 55490 3000 55496 3052
rect 55548 3040 55554 3052
rect 56045 3043 56103 3049
rect 56045 3040 56057 3043
rect 55548 3012 56057 3040
rect 55548 3000 55554 3012
rect 56045 3009 56057 3012
rect 56091 3009 56103 3043
rect 61749 3043 61807 3049
rect 61749 3040 61761 3043
rect 56045 3003 56103 3009
rect 59280 3012 61761 3040
rect 49329 2975 49387 2981
rect 49329 2972 49341 2975
rect 48976 2944 49341 2972
rect 48976 2848 49004 2944
rect 49329 2941 49341 2944
rect 49375 2941 49387 2975
rect 50246 2972 50252 2984
rect 50207 2944 50252 2972
rect 49329 2935 49387 2941
rect 50246 2932 50252 2944
rect 50304 2932 50310 2984
rect 50985 2975 51043 2981
rect 50985 2941 50997 2975
rect 51031 2972 51043 2975
rect 51350 2972 51356 2984
rect 51031 2944 51356 2972
rect 51031 2941 51043 2944
rect 50985 2935 51043 2941
rect 51350 2932 51356 2944
rect 51408 2932 51414 2984
rect 51902 2972 51908 2984
rect 51736 2944 51908 2972
rect 49234 2864 49240 2916
rect 49292 2904 49298 2916
rect 49513 2907 49571 2913
rect 49513 2904 49525 2907
rect 49292 2876 49525 2904
rect 49292 2864 49298 2876
rect 49513 2873 49525 2876
rect 49559 2873 49571 2907
rect 49513 2867 49571 2873
rect 49602 2864 49608 2916
rect 49660 2904 49666 2916
rect 51736 2913 51764 2944
rect 51902 2932 51908 2944
rect 51960 2932 51966 2984
rect 52454 2972 52460 2984
rect 52415 2944 52460 2972
rect 52454 2932 52460 2944
rect 52512 2932 52518 2984
rect 54018 2972 54024 2984
rect 53979 2944 54024 2972
rect 54018 2932 54024 2944
rect 54076 2932 54082 2984
rect 54662 2932 54668 2984
rect 54720 2972 54726 2984
rect 54757 2975 54815 2981
rect 54757 2972 54769 2975
rect 54720 2944 54769 2972
rect 54720 2932 54726 2944
rect 54757 2941 54769 2944
rect 54803 2941 54815 2975
rect 54757 2935 54815 2941
rect 56778 2932 56784 2984
rect 56836 2972 56842 2984
rect 57517 2975 57575 2981
rect 57517 2972 57529 2975
rect 56836 2944 57529 2972
rect 56836 2932 56842 2944
rect 57517 2941 57529 2944
rect 57563 2941 57575 2975
rect 57517 2935 57575 2941
rect 58342 2932 58348 2984
rect 58400 2972 58406 2984
rect 59280 2981 59308 3012
rect 61749 3009 61761 3012
rect 61795 3009 61807 3043
rect 61749 3003 61807 3009
rect 63218 3000 63224 3052
rect 63276 3040 63282 3052
rect 63405 3043 63463 3049
rect 63405 3040 63417 3043
rect 63276 3012 63417 3040
rect 63276 3000 63282 3012
rect 63405 3009 63417 3012
rect 63451 3009 63463 3043
rect 63405 3003 63463 3009
rect 67910 3000 67916 3052
rect 67968 3000 67974 3052
rect 59265 2975 59323 2981
rect 59265 2972 59277 2975
rect 58400 2944 59277 2972
rect 58400 2932 58406 2944
rect 59265 2941 59277 2944
rect 59311 2941 59323 2975
rect 59909 2975 59967 2981
rect 59909 2972 59921 2975
rect 59265 2935 59323 2941
rect 59740 2944 59921 2972
rect 50065 2907 50123 2913
rect 50065 2904 50077 2907
rect 49660 2876 50077 2904
rect 49660 2864 49666 2876
rect 50065 2873 50077 2876
rect 50111 2873 50123 2907
rect 50065 2867 50123 2873
rect 51721 2907 51779 2913
rect 51721 2873 51733 2907
rect 51767 2873 51779 2907
rect 51721 2867 51779 2873
rect 51810 2864 51816 2916
rect 51868 2904 51874 2916
rect 52914 2904 52920 2916
rect 51868 2876 52920 2904
rect 51868 2864 51874 2876
rect 52914 2864 52920 2876
rect 52972 2864 52978 2916
rect 53006 2864 53012 2916
rect 53064 2904 53070 2916
rect 53837 2907 53895 2913
rect 53837 2904 53849 2907
rect 53064 2876 53849 2904
rect 53064 2864 53070 2876
rect 53837 2873 53849 2876
rect 53883 2873 53895 2907
rect 53837 2867 53895 2873
rect 55214 2864 55220 2916
rect 55272 2904 55278 2916
rect 55493 2907 55551 2913
rect 55493 2904 55505 2907
rect 55272 2876 55505 2904
rect 55272 2864 55278 2876
rect 55493 2873 55505 2876
rect 55539 2873 55551 2907
rect 55493 2867 55551 2873
rect 56042 2864 56048 2916
rect 56100 2904 56106 2916
rect 56229 2907 56287 2913
rect 56229 2904 56241 2907
rect 56100 2876 56241 2904
rect 56100 2864 56106 2876
rect 56229 2873 56241 2876
rect 56275 2873 56287 2907
rect 56229 2867 56287 2873
rect 56318 2864 56324 2916
rect 56376 2904 56382 2916
rect 56965 2907 57023 2913
rect 56965 2904 56977 2907
rect 56376 2876 56977 2904
rect 56376 2864 56382 2876
rect 56965 2873 56977 2876
rect 57011 2873 57023 2907
rect 56965 2867 57023 2873
rect 57330 2864 57336 2916
rect 57388 2904 57394 2916
rect 57701 2907 57759 2913
rect 57701 2904 57713 2907
rect 57388 2876 57713 2904
rect 57388 2864 57394 2876
rect 57701 2873 57713 2876
rect 57747 2873 57759 2907
rect 57701 2867 57759 2873
rect 58986 2864 58992 2916
rect 59044 2904 59050 2916
rect 59740 2904 59768 2944
rect 59909 2941 59921 2944
rect 59955 2941 59967 2975
rect 59909 2935 59967 2941
rect 60274 2932 60280 2984
rect 60332 2972 60338 2984
rect 60369 2975 60427 2981
rect 60369 2972 60381 2975
rect 60332 2944 60381 2972
rect 60332 2932 60338 2944
rect 60369 2941 60381 2944
rect 60415 2941 60427 2975
rect 61194 2972 61200 2984
rect 61155 2944 61200 2972
rect 60369 2935 60427 2941
rect 61194 2932 61200 2944
rect 61252 2932 61258 2984
rect 62206 2932 62212 2984
rect 62264 2972 62270 2984
rect 62485 2975 62543 2981
rect 62485 2972 62497 2975
rect 62264 2944 62497 2972
rect 62264 2932 62270 2944
rect 62485 2941 62497 2944
rect 62531 2941 62543 2975
rect 62485 2935 62543 2941
rect 63954 2932 63960 2984
rect 64012 2972 64018 2984
rect 64509 2975 64567 2981
rect 64509 2972 64521 2975
rect 64012 2944 64521 2972
rect 64012 2932 64018 2944
rect 64509 2941 64521 2944
rect 64555 2941 64567 2975
rect 64509 2935 64567 2941
rect 64966 2932 64972 2984
rect 65024 2972 65030 2984
rect 65245 2975 65303 2981
rect 65245 2972 65257 2975
rect 65024 2944 65257 2972
rect 65024 2932 65030 2944
rect 65245 2941 65257 2944
rect 65291 2941 65303 2975
rect 65245 2935 65303 2941
rect 65702 2932 65708 2984
rect 65760 2972 65766 2984
rect 65981 2975 66039 2981
rect 65981 2972 65993 2975
rect 65760 2944 65993 2972
rect 65760 2932 65766 2944
rect 65981 2941 65993 2944
rect 66027 2941 66039 2975
rect 65981 2935 66039 2941
rect 66717 2975 66775 2981
rect 66717 2941 66729 2975
rect 66763 2972 66775 2975
rect 67928 2972 67956 3000
rect 66763 2944 67956 2972
rect 66763 2941 66775 2944
rect 66717 2935 66775 2941
rect 59044 2876 59768 2904
rect 59044 2864 59050 2876
rect 59814 2864 59820 2916
rect 59872 2904 59878 2916
rect 60292 2904 60320 2932
rect 61010 2904 61016 2916
rect 59872 2876 60320 2904
rect 60971 2876 61016 2904
rect 59872 2864 59878 2876
rect 61010 2864 61016 2876
rect 61068 2864 61074 2916
rect 62298 2904 62304 2916
rect 62259 2876 62304 2904
rect 62298 2864 62304 2876
rect 62356 2864 62362 2916
rect 63126 2864 63132 2916
rect 63184 2904 63190 2916
rect 63221 2907 63279 2913
rect 63221 2904 63233 2907
rect 63184 2876 63233 2904
rect 63184 2864 63190 2876
rect 63221 2873 63233 2876
rect 63267 2873 63279 2907
rect 63221 2867 63279 2873
rect 63586 2864 63592 2916
rect 63644 2904 63650 2916
rect 64325 2907 64383 2913
rect 64325 2904 64337 2907
rect 63644 2876 64337 2904
rect 63644 2864 63650 2876
rect 64325 2873 64337 2876
rect 64371 2873 64383 2907
rect 64325 2867 64383 2873
rect 64690 2864 64696 2916
rect 64748 2904 64754 2916
rect 65061 2907 65119 2913
rect 65061 2904 65073 2907
rect 64748 2876 65073 2904
rect 64748 2864 64754 2876
rect 65061 2873 65073 2876
rect 65107 2873 65119 2907
rect 65061 2867 65119 2873
rect 65334 2864 65340 2916
rect 65392 2904 65398 2916
rect 65797 2907 65855 2913
rect 65797 2904 65809 2907
rect 65392 2876 65809 2904
rect 65392 2864 65398 2876
rect 65797 2873 65809 2876
rect 65843 2873 65855 2907
rect 65797 2867 65855 2873
rect 67082 2864 67088 2916
rect 67140 2904 67146 2916
rect 67913 2907 67971 2913
rect 67913 2904 67925 2907
rect 67140 2876 67925 2904
rect 67140 2864 67146 2876
rect 67913 2873 67925 2876
rect 67959 2873 67971 2907
rect 67913 2867 67971 2873
rect 47084 2808 48912 2836
rect 47084 2796 47090 2808
rect 48958 2796 48964 2848
rect 49016 2796 49022 2848
rect 49970 2796 49976 2848
rect 50028 2836 50034 2848
rect 50893 2839 50951 2845
rect 50893 2836 50905 2839
rect 50028 2808 50905 2836
rect 50028 2796 50034 2808
rect 50893 2805 50905 2808
rect 50939 2805 50951 2839
rect 50893 2799 50951 2805
rect 51258 2796 51264 2848
rect 51316 2836 51322 2848
rect 54478 2836 54484 2848
rect 51316 2808 54484 2836
rect 51316 2796 51322 2808
rect 54478 2796 54484 2808
rect 54536 2796 54542 2848
rect 54754 2796 54760 2848
rect 54812 2836 54818 2848
rect 55401 2839 55459 2845
rect 55401 2836 55413 2839
rect 54812 2808 55413 2836
rect 54812 2796 54818 2808
rect 55401 2805 55413 2808
rect 55447 2805 55459 2839
rect 55401 2799 55459 2805
rect 55950 2796 55956 2848
rect 56008 2836 56014 2848
rect 56873 2839 56931 2845
rect 56873 2836 56885 2839
rect 56008 2808 56885 2836
rect 56008 2796 56014 2808
rect 56873 2805 56885 2808
rect 56919 2805 56931 2839
rect 56873 2799 56931 2805
rect 62206 2796 62212 2848
rect 62264 2836 62270 2848
rect 62666 2836 62672 2848
rect 62264 2808 62672 2836
rect 62264 2796 62270 2808
rect 62666 2796 62672 2808
rect 62724 2796 62730 2848
rect 65702 2796 65708 2848
rect 65760 2836 65766 2848
rect 66625 2839 66683 2845
rect 66625 2836 66637 2839
rect 65760 2808 66637 2836
rect 65760 2796 65766 2808
rect 66625 2805 66637 2808
rect 66671 2805 66683 2839
rect 66625 2799 66683 2805
rect 32180 2536 32260 2564
rect 32324 2740 33732 2768
rect 32180 2524 32186 2536
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2496 1547 2499
rect 1578 2496 1584 2508
rect 1535 2468 1584 2496
rect 1535 2465 1547 2468
rect 1489 2459 1547 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 6362 2496 6368 2508
rect 4479 2468 6368 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 7708 2468 9597 2496
rect 7708 2456 7714 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 10226 2456 10232 2508
rect 10284 2496 10290 2508
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 10284 2468 11161 2496
rect 10284 2456 10290 2468
rect 11149 2465 11161 2468
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2496 11391 2499
rect 13906 2496 13912 2508
rect 11379 2468 13912 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14148 2468 14657 2496
rect 14148 2456 14154 2468
rect 14645 2465 14657 2468
rect 14691 2496 14703 2499
rect 18598 2496 18604 2508
rect 14691 2468 18604 2496
rect 14691 2465 14703 2468
rect 14645 2459 14703 2465
rect 18598 2456 18604 2468
rect 18656 2456 18662 2508
rect 31662 2456 31668 2508
rect 31720 2496 31726 2508
rect 32324 2496 32352 2740
rect 33318 2700 33324 2712
rect 33279 2672 33324 2700
rect 33318 2660 33324 2672
rect 33376 2660 33382 2712
rect 33704 2700 33732 2740
rect 37628 2746 68816 2768
rect 36722 2700 36728 2712
rect 33704 2672 36728 2700
rect 36722 2660 36728 2672
rect 36780 2660 36786 2712
rect 37628 2694 39246 2746
rect 39298 2694 39310 2746
rect 39362 2694 39374 2746
rect 39426 2694 39438 2746
rect 39490 2694 49246 2746
rect 49298 2694 49310 2746
rect 49362 2694 49374 2746
rect 49426 2694 49438 2746
rect 49490 2694 59246 2746
rect 59298 2694 59310 2746
rect 59362 2694 59374 2746
rect 59426 2694 59438 2746
rect 59490 2694 68816 2746
rect 37628 2672 68816 2694
rect 32766 2592 32772 2644
rect 32824 2632 32830 2644
rect 44269 2635 44327 2641
rect 44269 2632 44281 2635
rect 32824 2604 44281 2632
rect 32824 2592 32830 2604
rect 44269 2601 44281 2604
rect 44315 2601 44327 2635
rect 44269 2595 44327 2601
rect 48498 2592 48504 2644
rect 48556 2632 48562 2644
rect 49605 2635 49663 2641
rect 49605 2632 49617 2635
rect 48556 2604 49617 2632
rect 48556 2592 48562 2604
rect 49605 2601 49617 2604
rect 49651 2601 49663 2635
rect 49605 2595 49663 2601
rect 49786 2592 49792 2644
rect 49844 2632 49850 2644
rect 51537 2635 51595 2641
rect 51537 2632 51549 2635
rect 49844 2604 51549 2632
rect 49844 2592 49850 2604
rect 51537 2601 51549 2604
rect 51583 2601 51595 2635
rect 54202 2632 54208 2644
rect 54163 2604 54208 2632
rect 51537 2595 51595 2601
rect 54202 2592 54208 2604
rect 54260 2592 54266 2644
rect 57514 2592 57520 2644
rect 57572 2632 57578 2644
rect 58526 2632 58532 2644
rect 57572 2604 58532 2632
rect 57572 2592 57578 2604
rect 58526 2592 58532 2604
rect 58584 2592 58590 2644
rect 60642 2592 60648 2644
rect 60700 2632 60706 2644
rect 63681 2635 63739 2641
rect 63681 2632 63693 2635
rect 60700 2604 63693 2632
rect 60700 2592 60706 2604
rect 63681 2601 63693 2604
rect 63727 2601 63739 2635
rect 63681 2595 63739 2601
rect 66346 2592 66352 2644
rect 66404 2632 66410 2644
rect 66404 2604 67956 2632
rect 66404 2592 66410 2604
rect 33410 2564 33416 2576
rect 33371 2536 33416 2564
rect 33410 2524 33416 2536
rect 33468 2524 33474 2576
rect 33686 2524 33692 2576
rect 33744 2564 33750 2576
rect 33965 2567 34023 2573
rect 33965 2564 33977 2567
rect 33744 2536 33977 2564
rect 33744 2524 33750 2536
rect 33965 2533 33977 2536
rect 34011 2533 34023 2567
rect 33965 2527 34023 2533
rect 38930 2524 38936 2576
rect 38988 2564 38994 2576
rect 39209 2567 39267 2573
rect 39209 2564 39221 2567
rect 38988 2536 39221 2564
rect 38988 2524 38994 2536
rect 39209 2533 39221 2536
rect 39255 2533 39267 2567
rect 39209 2527 39267 2533
rect 39850 2524 39856 2576
rect 39908 2564 39914 2576
rect 40310 2564 40316 2576
rect 39908 2536 40316 2564
rect 39908 2524 39914 2536
rect 40310 2524 40316 2536
rect 40368 2524 40374 2576
rect 40954 2564 40960 2576
rect 40915 2536 40960 2564
rect 40954 2524 40960 2536
rect 41012 2524 41018 2576
rect 42426 2564 42432 2576
rect 42387 2536 42432 2564
rect 42426 2524 42432 2536
rect 42484 2524 42490 2576
rect 43162 2524 43168 2576
rect 43220 2564 43226 2576
rect 43625 2567 43683 2573
rect 43625 2564 43637 2567
rect 43220 2536 43637 2564
rect 43220 2524 43226 2536
rect 43625 2533 43637 2536
rect 43671 2533 43683 2567
rect 43625 2527 43683 2533
rect 44361 2567 44419 2573
rect 44361 2533 44373 2567
rect 44407 2564 44419 2567
rect 44542 2564 44548 2576
rect 44407 2536 44548 2564
rect 44407 2533 44419 2536
rect 44361 2527 44419 2533
rect 44542 2524 44548 2536
rect 44600 2524 44606 2576
rect 45097 2567 45155 2573
rect 45097 2533 45109 2567
rect 45143 2564 45155 2567
rect 46014 2564 46020 2576
rect 45143 2536 46020 2564
rect 45143 2533 45155 2536
rect 45097 2527 45155 2533
rect 46014 2524 46020 2536
rect 46072 2524 46078 2576
rect 46290 2564 46296 2576
rect 46251 2536 46296 2564
rect 46290 2524 46296 2536
rect 46348 2524 46354 2576
rect 46658 2524 46664 2576
rect 46716 2564 46722 2576
rect 47029 2567 47087 2573
rect 47029 2564 47041 2567
rect 46716 2536 47041 2564
rect 46716 2524 46722 2536
rect 47029 2533 47041 2536
rect 47075 2533 47087 2567
rect 47029 2527 47087 2533
rect 47765 2567 47823 2573
rect 47765 2533 47777 2567
rect 47811 2564 47823 2567
rect 48314 2564 48320 2576
rect 47811 2536 48320 2564
rect 47811 2533 47823 2536
rect 47765 2527 47823 2533
rect 48314 2524 48320 2536
rect 48372 2524 48378 2576
rect 48682 2524 48688 2576
rect 48740 2564 48746 2576
rect 48777 2567 48835 2573
rect 48777 2564 48789 2567
rect 48740 2536 48789 2564
rect 48740 2524 48746 2536
rect 48777 2533 48789 2536
rect 48823 2533 48835 2567
rect 48777 2527 48835 2533
rect 48866 2524 48872 2576
rect 48924 2564 48930 2576
rect 48961 2567 49019 2573
rect 48961 2564 48973 2567
rect 48924 2536 48973 2564
rect 48924 2524 48930 2536
rect 48961 2533 48973 2536
rect 49007 2533 49019 2567
rect 49694 2564 49700 2576
rect 49655 2536 49700 2564
rect 48961 2527 49019 2533
rect 49694 2524 49700 2536
rect 49752 2524 49758 2576
rect 50062 2524 50068 2576
rect 50120 2564 50126 2576
rect 50249 2567 50307 2573
rect 50249 2564 50261 2567
rect 50120 2536 50261 2564
rect 50120 2524 50126 2536
rect 50249 2533 50261 2536
rect 50295 2533 50307 2567
rect 50430 2564 50436 2576
rect 50391 2536 50436 2564
rect 50249 2527 50307 2533
rect 50430 2524 50436 2536
rect 50488 2524 50494 2576
rect 51626 2564 51632 2576
rect 51587 2536 51632 2564
rect 51626 2524 51632 2536
rect 51684 2524 51690 2576
rect 52917 2567 52975 2573
rect 52917 2564 52929 2567
rect 52012 2536 52929 2564
rect 31720 2468 32352 2496
rect 38473 2499 38531 2505
rect 31720 2456 31726 2468
rect 38473 2465 38485 2499
rect 38519 2496 38531 2499
rect 41693 2499 41751 2505
rect 38519 2468 39896 2496
rect 38519 2465 38531 2468
rect 38473 2459 38531 2465
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2087 2400 2605 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2593 2397 2605 2400
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 32858 2428 32864 2440
rect 3283 2400 32864 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 32858 2388 32864 2400
rect 32916 2388 32922 2440
rect 39868 2437 39896 2468
rect 41693 2465 41705 2499
rect 41739 2496 41751 2499
rect 42702 2496 42708 2508
rect 41739 2468 42708 2496
rect 41739 2465 41751 2468
rect 41693 2459 41751 2465
rect 42702 2456 42708 2468
rect 42760 2456 42766 2508
rect 49234 2456 49240 2508
rect 49292 2496 49298 2508
rect 52012 2496 52040 2536
rect 52917 2533 52929 2536
rect 52963 2533 52975 2567
rect 52917 2527 52975 2533
rect 53101 2567 53159 2573
rect 53101 2533 53113 2567
rect 53147 2564 53159 2567
rect 53466 2564 53472 2576
rect 53147 2536 53472 2564
rect 53147 2533 53159 2536
rect 53101 2527 53159 2533
rect 53466 2524 53472 2536
rect 53524 2524 53530 2576
rect 53742 2524 53748 2576
rect 53800 2564 53806 2576
rect 54297 2567 54355 2573
rect 54297 2564 54309 2567
rect 53800 2536 54309 2564
rect 53800 2524 53806 2536
rect 54297 2533 54309 2536
rect 54343 2533 54355 2567
rect 54297 2527 54355 2533
rect 54478 2524 54484 2576
rect 54536 2564 54542 2576
rect 54849 2567 54907 2573
rect 54849 2564 54861 2567
rect 54536 2536 54861 2564
rect 54536 2524 54542 2536
rect 54849 2533 54861 2536
rect 54895 2533 54907 2567
rect 54849 2527 54907 2533
rect 55033 2567 55091 2573
rect 55033 2533 55045 2567
rect 55079 2564 55091 2567
rect 55306 2564 55312 2576
rect 55079 2536 55312 2564
rect 55079 2533 55091 2536
rect 55033 2527 55091 2533
rect 55306 2524 55312 2536
rect 55364 2524 55370 2576
rect 55769 2567 55827 2573
rect 55769 2533 55781 2567
rect 55815 2564 55827 2567
rect 55858 2564 55864 2576
rect 55815 2536 55864 2564
rect 55815 2533 55827 2536
rect 55769 2527 55827 2533
rect 55858 2524 55864 2536
rect 55916 2524 55922 2576
rect 56962 2564 56968 2576
rect 56923 2536 56968 2564
rect 56962 2524 56968 2536
rect 57020 2524 57026 2576
rect 57793 2567 57851 2573
rect 57793 2533 57805 2567
rect 57839 2564 57851 2567
rect 58158 2564 58164 2576
rect 57839 2536 58164 2564
rect 57839 2533 57851 2536
rect 57793 2527 57851 2533
rect 58158 2524 58164 2536
rect 58216 2524 58222 2576
rect 59354 2564 59360 2576
rect 58452 2536 59360 2564
rect 52178 2496 52184 2508
rect 49292 2468 52040 2496
rect 52139 2468 52184 2496
rect 49292 2456 49298 2468
rect 52178 2456 52184 2468
rect 52236 2456 52242 2508
rect 52365 2499 52423 2505
rect 52365 2465 52377 2499
rect 52411 2465 52423 2499
rect 52365 2459 52423 2465
rect 57149 2499 57207 2505
rect 57149 2465 57161 2499
rect 57195 2496 57207 2499
rect 58452 2496 58480 2536
rect 59354 2524 59360 2536
rect 59412 2524 59418 2576
rect 59630 2564 59636 2576
rect 59591 2536 59636 2564
rect 59630 2524 59636 2536
rect 59688 2524 59694 2576
rect 60369 2567 60427 2573
rect 60369 2533 60381 2567
rect 60415 2564 60427 2567
rect 60550 2564 60556 2576
rect 60415 2536 60556 2564
rect 60415 2533 60427 2536
rect 60369 2527 60427 2533
rect 60550 2524 60556 2536
rect 60608 2524 60614 2576
rect 61102 2564 61108 2576
rect 61063 2536 61108 2564
rect 61102 2524 61108 2536
rect 61160 2524 61166 2576
rect 61838 2524 61844 2576
rect 61896 2564 61902 2576
rect 62301 2567 62359 2573
rect 62301 2564 62313 2567
rect 61896 2536 62313 2564
rect 61896 2524 61902 2536
rect 62301 2533 62313 2536
rect 62347 2533 62359 2567
rect 63770 2564 63776 2576
rect 63731 2536 63776 2564
rect 62301 2527 62359 2533
rect 63770 2524 63776 2536
rect 63828 2524 63834 2576
rect 64969 2567 65027 2573
rect 64969 2533 64981 2567
rect 65015 2564 65027 2567
rect 65242 2564 65248 2576
rect 65015 2536 65248 2564
rect 65015 2533 65027 2536
rect 64969 2527 65027 2533
rect 65242 2524 65248 2536
rect 65300 2524 65306 2576
rect 65518 2524 65524 2576
rect 65576 2564 65582 2576
rect 65705 2567 65763 2573
rect 65705 2564 65717 2567
rect 65576 2536 65717 2564
rect 65576 2524 65582 2536
rect 65705 2533 65717 2536
rect 65751 2533 65763 2567
rect 65705 2527 65763 2533
rect 65794 2524 65800 2576
rect 65852 2564 65858 2576
rect 66257 2567 66315 2573
rect 66257 2564 66269 2567
rect 65852 2536 66269 2564
rect 65852 2524 65858 2536
rect 66257 2533 66269 2536
rect 66303 2533 66315 2567
rect 66257 2527 66315 2533
rect 66441 2567 66499 2573
rect 66441 2533 66453 2567
rect 66487 2564 66499 2567
rect 67358 2564 67364 2576
rect 66487 2536 67364 2564
rect 66487 2533 66499 2536
rect 66441 2527 66499 2533
rect 67358 2524 67364 2536
rect 67416 2524 67422 2576
rect 67928 2573 67956 2604
rect 67913 2567 67971 2573
rect 67913 2533 67925 2567
rect 67959 2533 67971 2567
rect 67913 2527 67971 2533
rect 57195 2468 58480 2496
rect 57195 2465 57207 2468
rect 57149 2459 57207 2465
rect 35437 2431 35495 2437
rect 35437 2397 35449 2431
rect 35483 2428 35495 2431
rect 39025 2431 39083 2437
rect 39025 2428 39037 2431
rect 35483 2400 39037 2428
rect 35483 2397 35495 2400
rect 35437 2391 35495 2397
rect 39025 2397 39037 2400
rect 39071 2397 39083 2431
rect 39025 2391 39083 2397
rect 39853 2431 39911 2437
rect 39853 2397 39865 2431
rect 39899 2428 39911 2431
rect 39899 2400 46980 2428
rect 39899 2397 39911 2400
rect 39853 2391 39911 2397
rect 290 2320 296 2372
rect 348 2360 354 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 348 2332 4261 2360
rect 348 2320 354 2332
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 6362 2320 6368 2372
rect 6420 2360 6426 2372
rect 6917 2363 6975 2369
rect 6917 2360 6929 2363
rect 6420 2332 6929 2360
rect 6420 2320 6426 2332
rect 6917 2329 6929 2332
rect 6963 2329 6975 2363
rect 6917 2323 6975 2329
rect 7282 2320 7288 2372
rect 7340 2360 7346 2372
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 7340 2332 8401 2360
rect 7340 2320 7346 2332
rect 8389 2329 8401 2332
rect 8435 2329 8447 2363
rect 8389 2323 8447 2329
rect 12529 2363 12587 2369
rect 12529 2329 12541 2363
rect 12575 2360 12587 2363
rect 15102 2360 15108 2372
rect 12575 2332 14964 2360
rect 15063 2332 15108 2360
rect 12575 2329 12587 2332
rect 12529 2323 12587 2329
rect 5813 2295 5871 2301
rect 5813 2261 5825 2295
rect 5859 2292 5871 2295
rect 5902 2292 5908 2304
rect 5859 2264 5908 2292
rect 5859 2261 5871 2264
rect 5813 2255 5871 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 7745 2295 7803 2301
rect 7745 2292 7757 2295
rect 6788 2264 7757 2292
rect 6788 2252 6794 2264
rect 7745 2261 7757 2264
rect 7791 2261 7803 2295
rect 7745 2255 7803 2261
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 8168 2264 10425 2292
rect 8168 2252 8174 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 13173 2295 13231 2301
rect 13173 2261 13185 2295
rect 13219 2292 13231 2295
rect 13722 2292 13728 2304
rect 13219 2264 13728 2292
rect 13219 2261 13231 2264
rect 13173 2255 13231 2261
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 14090 2292 14096 2304
rect 13955 2264 14096 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 14936 2292 14964 2332
rect 15102 2320 15108 2332
rect 15160 2320 15166 2372
rect 33594 2360 33600 2372
rect 16500 2332 22094 2360
rect 33555 2332 33600 2360
rect 16500 2292 16528 2332
rect 14936 2264 16528 2292
rect 17497 2295 17555 2301
rect 17497 2261 17509 2295
rect 17543 2292 17555 2295
rect 17586 2292 17592 2304
rect 17543 2264 17592 2292
rect 17543 2261 17555 2264
rect 17497 2255 17555 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 18141 2295 18199 2301
rect 18141 2261 18153 2295
rect 18187 2292 18199 2295
rect 19426 2292 19432 2304
rect 18187 2264 19432 2292
rect 18187 2261 18199 2264
rect 18141 2255 18199 2261
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 1104 2202 18952 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 14246 2202
rect 14298 2150 14310 2202
rect 14362 2150 14374 2202
rect 14426 2150 14438 2202
rect 14490 2150 18952 2202
rect 1104 2128 18952 2150
rect 13906 2048 13912 2100
rect 13964 2088 13970 2100
rect 17218 2088 17224 2100
rect 13964 2060 17224 2088
rect 13964 2048 13970 2060
rect 17218 2048 17224 2060
rect 17276 2048 17282 2100
rect 22066 2088 22094 2332
rect 33594 2320 33600 2332
rect 33652 2320 33658 2372
rect 37277 2363 37335 2369
rect 37277 2329 37289 2363
rect 37323 2360 37335 2363
rect 38289 2363 38347 2369
rect 38289 2360 38301 2363
rect 37323 2332 38301 2360
rect 37323 2329 37335 2332
rect 37277 2323 37335 2329
rect 38289 2329 38301 2332
rect 38335 2329 38347 2363
rect 40773 2363 40831 2369
rect 40773 2360 40785 2363
rect 38289 2323 38347 2329
rect 38396 2332 40785 2360
rect 38396 2292 38424 2332
rect 40773 2329 40785 2332
rect 40819 2329 40831 2363
rect 40773 2323 40831 2329
rect 42426 2320 42432 2372
rect 42484 2360 42490 2372
rect 46842 2360 46848 2372
rect 42484 2332 46336 2360
rect 46803 2332 46848 2360
rect 42484 2320 42490 2332
rect 41598 2292 41604 2304
rect 31726 2264 38424 2292
rect 41559 2264 41604 2292
rect 22922 2156 22928 2168
rect 22883 2128 22928 2156
rect 22922 2116 22928 2128
rect 22980 2116 22986 2168
rect 23198 2088 23204 2100
rect 22066 2060 23204 2088
rect 23198 2048 23204 2060
rect 23256 2048 23262 2100
rect 31726 2088 31754 2264
rect 41598 2252 41604 2264
rect 41656 2252 41662 2304
rect 42334 2292 42340 2304
rect 42295 2264 42340 2292
rect 42334 2252 42340 2264
rect 42392 2252 42398 2304
rect 43530 2292 43536 2304
rect 43491 2264 43536 2292
rect 43530 2252 43536 2264
rect 43588 2252 43594 2304
rect 43714 2252 43720 2304
rect 43772 2292 43778 2304
rect 45005 2295 45063 2301
rect 45005 2292 45017 2295
rect 43772 2264 45017 2292
rect 43772 2252 43778 2264
rect 45005 2261 45017 2264
rect 45051 2261 45063 2295
rect 45005 2255 45063 2261
rect 45094 2252 45100 2304
rect 45152 2292 45158 2304
rect 46201 2295 46259 2301
rect 46201 2292 46213 2295
rect 45152 2264 46213 2292
rect 45152 2252 45158 2264
rect 46201 2261 46213 2264
rect 46247 2261 46259 2295
rect 46308 2292 46336 2332
rect 46842 2320 46848 2332
rect 46900 2320 46906 2372
rect 46952 2360 46980 2400
rect 49786 2388 49792 2440
rect 49844 2428 49850 2440
rect 52380 2428 52408 2459
rect 58526 2456 58532 2508
rect 58584 2505 58590 2508
rect 58584 2496 58595 2505
rect 58584 2468 58629 2496
rect 58584 2459 58595 2468
rect 58584 2456 58590 2459
rect 61930 2456 61936 2508
rect 61988 2496 61994 2508
rect 63037 2499 63095 2505
rect 63037 2496 63049 2499
rect 61988 2468 63049 2496
rect 61988 2456 61994 2468
rect 63037 2465 63049 2468
rect 63083 2465 63095 2499
rect 63037 2459 63095 2465
rect 65150 2456 65156 2508
rect 65208 2496 65214 2508
rect 67085 2499 67143 2505
rect 67085 2496 67097 2499
rect 65208 2468 67097 2496
rect 65208 2456 65214 2468
rect 67085 2465 67097 2468
rect 67131 2465 67143 2499
rect 67085 2459 67143 2465
rect 49844 2400 52408 2428
rect 49844 2388 49850 2400
rect 58894 2388 58900 2440
rect 58952 2428 58958 2440
rect 60921 2431 60979 2437
rect 60921 2428 60933 2431
rect 58952 2400 60933 2428
rect 58952 2388 58958 2400
rect 60921 2397 60933 2400
rect 60967 2397 60979 2431
rect 62853 2431 62911 2437
rect 62853 2428 62865 2431
rect 60921 2391 60979 2397
rect 61396 2400 62865 2428
rect 46952 2332 51074 2360
rect 47673 2295 47731 2301
rect 47673 2292 47685 2295
rect 46308 2264 47685 2292
rect 46201 2255 46259 2261
rect 47673 2261 47685 2264
rect 47719 2261 47731 2295
rect 51046 2292 51074 2332
rect 52086 2320 52092 2372
rect 52144 2360 52150 2372
rect 55585 2363 55643 2369
rect 55585 2360 55597 2363
rect 52144 2332 55597 2360
rect 52144 2320 52150 2332
rect 55585 2329 55597 2332
rect 55631 2329 55643 2363
rect 57606 2360 57612 2372
rect 57567 2332 57612 2360
rect 55585 2323 55643 2329
rect 57606 2320 57612 2332
rect 57664 2320 57670 2372
rect 58066 2320 58072 2372
rect 58124 2360 58130 2372
rect 59449 2363 59507 2369
rect 59449 2360 59461 2363
rect 58124 2332 59461 2360
rect 58124 2320 58130 2332
rect 59449 2329 59461 2332
rect 59495 2329 59507 2363
rect 59449 2323 59507 2329
rect 60182 2320 60188 2372
rect 60240 2360 60246 2372
rect 61396 2360 61424 2400
rect 62853 2397 62865 2400
rect 62899 2397 62911 2431
rect 62853 2391 62911 2397
rect 63402 2388 63408 2440
rect 63460 2428 63466 2440
rect 65521 2431 65579 2437
rect 65521 2428 65533 2431
rect 63460 2400 65533 2428
rect 63460 2388 63466 2400
rect 65521 2397 65533 2400
rect 65567 2397 65579 2431
rect 65521 2391 65579 2397
rect 60240 2332 61424 2360
rect 60240 2320 60246 2332
rect 61470 2320 61476 2372
rect 61528 2360 61534 2372
rect 62117 2363 62175 2369
rect 62117 2360 62129 2363
rect 61528 2332 62129 2360
rect 61528 2320 61534 2332
rect 62117 2329 62129 2332
rect 62163 2329 62175 2363
rect 62117 2323 62175 2329
rect 64785 2363 64843 2369
rect 64785 2329 64797 2363
rect 64831 2329 64843 2363
rect 64785 2323 64843 2329
rect 68097 2363 68155 2369
rect 68097 2329 68109 2363
rect 68143 2360 68155 2363
rect 68186 2360 68192 2372
rect 68143 2332 68192 2360
rect 68143 2329 68155 2332
rect 68097 2323 68155 2329
rect 58434 2292 58440 2304
rect 51046 2264 58440 2292
rect 47673 2255 47731 2261
rect 58434 2252 58440 2264
rect 58492 2252 58498 2304
rect 58526 2252 58532 2304
rect 58584 2292 58590 2304
rect 60277 2295 60335 2301
rect 60277 2292 60289 2295
rect 58584 2264 60289 2292
rect 58584 2252 58590 2264
rect 60277 2261 60289 2264
rect 60323 2261 60335 2295
rect 60277 2255 60335 2261
rect 61562 2252 61568 2304
rect 61620 2292 61626 2304
rect 64800 2292 64828 2323
rect 68186 2320 68192 2332
rect 68244 2320 68250 2372
rect 61620 2264 64828 2292
rect 61620 2252 61626 2264
rect 37628 2202 68816 2224
rect 37628 2150 44246 2202
rect 44298 2150 44310 2202
rect 44362 2150 44374 2202
rect 44426 2150 44438 2202
rect 44490 2150 54246 2202
rect 54298 2150 54310 2202
rect 54362 2150 54374 2202
rect 54426 2150 54438 2202
rect 54490 2150 64246 2202
rect 64298 2150 64310 2202
rect 64362 2150 64374 2202
rect 64426 2150 64438 2202
rect 64490 2150 68816 2202
rect 37628 2128 68816 2150
rect 26160 2060 31754 2088
rect 14090 1980 14096 2032
rect 14148 2020 14154 2032
rect 21082 2020 21088 2032
rect 14148 1992 21088 2020
rect 14148 1980 14154 1992
rect 21082 1980 21088 1992
rect 21140 1980 21146 2032
rect 22830 1980 22836 2032
rect 22888 2020 22894 2032
rect 23290 2020 23296 2032
rect 22888 1992 23296 2020
rect 22888 1980 22894 1992
rect 23290 1980 23296 1992
rect 23348 1980 23354 2032
rect 13722 1912 13728 1964
rect 13780 1952 13786 1964
rect 21910 1952 21916 1964
rect 13780 1924 21916 1952
rect 13780 1912 13786 1924
rect 21910 1912 21916 1924
rect 21968 1912 21974 1964
rect 22094 1952 22100 1964
rect 22055 1924 22100 1952
rect 22094 1912 22100 1924
rect 22152 1912 22158 1964
rect 26160 1896 26188 2060
rect 32214 2048 32220 2100
rect 32272 2088 32278 2100
rect 39666 2088 39672 2100
rect 32272 2060 39672 2088
rect 32272 2048 32278 2060
rect 39666 2048 39672 2060
rect 39724 2048 39730 2100
rect 39761 2091 39819 2097
rect 39761 2057 39773 2091
rect 39807 2088 39819 2091
rect 39942 2088 39948 2100
rect 39807 2060 39948 2088
rect 39807 2057 39819 2060
rect 39761 2051 39819 2057
rect 39942 2048 39948 2060
rect 40000 2048 40006 2100
rect 41046 2048 41052 2100
rect 41104 2088 41110 2100
rect 46842 2088 46848 2100
rect 41104 2060 46848 2088
rect 41104 2048 41110 2060
rect 46842 2048 46848 2060
rect 46900 2048 46906 2100
rect 49326 2048 49332 2100
rect 49384 2088 49390 2100
rect 51074 2088 51080 2100
rect 49384 2060 51080 2088
rect 49384 2048 49390 2060
rect 51074 2048 51080 2060
rect 51132 2048 51138 2100
rect 30929 2023 30987 2029
rect 30929 1989 30941 2023
rect 30975 2020 30987 2023
rect 37277 2023 37335 2029
rect 37277 2020 37289 2023
rect 30975 1992 37289 2020
rect 30975 1989 30987 1992
rect 30929 1983 30987 1989
rect 37277 1989 37289 1992
rect 37323 1989 37335 2023
rect 37277 1983 37335 1989
rect 38562 1980 38568 2032
rect 38620 2020 38626 2032
rect 45094 2020 45100 2032
rect 38620 1992 45100 2020
rect 38620 1980 38626 1992
rect 45094 1980 45100 1992
rect 45152 1980 45158 2032
rect 26326 1952 26332 1964
rect 26287 1924 26332 1952
rect 26326 1912 26332 1924
rect 26384 1912 26390 1964
rect 26510 1952 26516 1964
rect 26471 1924 26516 1952
rect 26510 1912 26516 1924
rect 26568 1912 26574 1964
rect 26602 1912 26608 1964
rect 26660 1952 26666 1964
rect 26878 1952 26884 1964
rect 26660 1924 26705 1952
rect 26839 1924 26884 1952
rect 26660 1912 26666 1924
rect 26878 1912 26884 1924
rect 26936 1912 26942 1964
rect 27154 1952 27160 1964
rect 27115 1924 27160 1952
rect 27154 1912 27160 1924
rect 27212 1912 27218 1964
rect 27430 1952 27436 1964
rect 27391 1924 27436 1952
rect 27430 1912 27436 1924
rect 27488 1912 27494 1964
rect 27614 1952 27620 1964
rect 27575 1924 27620 1952
rect 27614 1912 27620 1924
rect 27672 1912 27678 1964
rect 27890 1952 27896 1964
rect 27851 1924 27896 1952
rect 27890 1912 27896 1924
rect 27948 1912 27954 1964
rect 28718 1952 28724 1964
rect 28679 1924 28724 1952
rect 28718 1912 28724 1924
rect 28776 1912 28782 1964
rect 28994 1952 29000 1964
rect 28955 1924 29000 1952
rect 28994 1912 29000 1924
rect 29052 1912 29058 1964
rect 29178 1952 29184 1964
rect 29139 1924 29184 1952
rect 29178 1912 29184 1924
rect 29236 1912 29242 1964
rect 29270 1912 29276 1964
rect 29328 1952 29334 1964
rect 31754 1952 31760 1964
rect 29328 1924 31760 1952
rect 29328 1912 29334 1924
rect 31754 1912 31760 1924
rect 31812 1912 31818 1964
rect 34146 1952 34152 1964
rect 34107 1924 34152 1952
rect 34146 1912 34152 1924
rect 34204 1912 34210 1964
rect 34422 1952 34428 1964
rect 34383 1924 34428 1952
rect 34422 1912 34428 1924
rect 34480 1912 34486 1964
rect 36449 1955 36507 1961
rect 36449 1921 36461 1955
rect 36495 1952 36507 1955
rect 41598 1952 41604 1964
rect 36495 1924 41604 1952
rect 36495 1921 36507 1924
rect 36449 1915 36507 1921
rect 41598 1912 41604 1924
rect 41656 1912 41662 1964
rect 46842 1912 46848 1964
rect 46900 1952 46906 1964
rect 47946 1952 47952 1964
rect 46900 1924 47952 1952
rect 46900 1912 46906 1924
rect 47946 1912 47952 1924
rect 48004 1912 48010 1964
rect 16574 1844 16580 1896
rect 16632 1884 16638 1896
rect 19058 1884 19064 1896
rect 16632 1856 19064 1884
rect 16632 1844 16638 1856
rect 19058 1844 19064 1856
rect 19116 1844 19122 1896
rect 25314 1884 25320 1896
rect 25275 1856 25320 1884
rect 25314 1844 25320 1856
rect 25372 1844 25378 1896
rect 25590 1884 25596 1896
rect 25551 1856 25596 1884
rect 25590 1844 25596 1856
rect 25648 1844 25654 1896
rect 25774 1884 25780 1896
rect 25735 1856 25780 1884
rect 25774 1844 25780 1856
rect 25832 1844 25838 1896
rect 25866 1844 25872 1896
rect 25924 1884 25930 1896
rect 26050 1884 26056 1896
rect 25924 1856 25969 1884
rect 26011 1856 26056 1884
rect 25924 1844 25930 1856
rect 26050 1844 26056 1856
rect 26108 1844 26114 1896
rect 26142 1844 26148 1896
rect 26200 1844 26206 1896
rect 26786 1884 26792 1896
rect 26747 1856 26792 1884
rect 26786 1844 26792 1856
rect 26844 1844 26850 1896
rect 27338 1884 27344 1896
rect 27299 1856 27344 1884
rect 27338 1844 27344 1856
rect 27396 1844 27402 1896
rect 28442 1844 28448 1896
rect 28500 1884 28506 1896
rect 31938 1884 31944 1896
rect 28500 1856 31944 1884
rect 28500 1844 28506 1856
rect 31938 1844 31944 1856
rect 31996 1844 32002 1896
rect 36541 1887 36599 1893
rect 36541 1853 36553 1887
rect 36587 1884 36599 1887
rect 42334 1884 42340 1896
rect 36587 1856 42340 1884
rect 36587 1853 36599 1856
rect 36541 1847 36599 1853
rect 42334 1844 42340 1856
rect 42392 1844 42398 1896
rect 44174 1844 44180 1896
rect 44232 1884 44238 1896
rect 46934 1884 46940 1896
rect 44232 1856 46940 1884
rect 44232 1844 44238 1856
rect 46934 1844 46940 1856
rect 46992 1844 46998 1896
rect 12342 1776 12348 1828
rect 12400 1816 12406 1828
rect 19153 1819 19211 1825
rect 19153 1816 19165 1819
rect 12400 1788 19165 1816
rect 12400 1776 12406 1788
rect 19153 1785 19165 1788
rect 19199 1785 19211 1819
rect 19153 1779 19211 1785
rect 25225 1819 25283 1825
rect 25225 1785 25237 1819
rect 25271 1816 25283 1819
rect 25498 1816 25504 1828
rect 25271 1788 25504 1816
rect 25271 1785 25283 1788
rect 25225 1779 25283 1785
rect 25498 1776 25504 1788
rect 25556 1776 25562 1828
rect 35437 1819 35495 1825
rect 35437 1816 35449 1819
rect 26206 1788 35449 1816
rect 13906 1708 13912 1760
rect 13964 1748 13970 1760
rect 14642 1748 14648 1760
rect 13964 1720 14648 1748
rect 13964 1708 13970 1720
rect 14642 1708 14648 1720
rect 14700 1708 14706 1760
rect 17586 1708 17592 1760
rect 17644 1748 17650 1760
rect 19242 1748 19248 1760
rect 17644 1720 19248 1748
rect 17644 1708 17650 1720
rect 19242 1708 19248 1720
rect 19300 1708 19306 1760
rect 22186 1708 22192 1760
rect 22244 1748 22250 1760
rect 22646 1748 22652 1760
rect 22244 1720 22652 1748
rect 22244 1708 22250 1720
rect 22646 1708 22652 1720
rect 22704 1708 22710 1760
rect 25682 1708 25688 1760
rect 25740 1748 25746 1760
rect 26206 1748 26234 1788
rect 35437 1785 35449 1788
rect 35483 1785 35495 1819
rect 35437 1779 35495 1785
rect 39942 1776 39948 1828
rect 40000 1816 40006 1828
rect 43990 1816 43996 1828
rect 40000 1788 43996 1816
rect 40000 1776 40006 1788
rect 43990 1776 43996 1788
rect 44048 1776 44054 1828
rect 28626 1748 28632 1760
rect 25740 1720 26234 1748
rect 28587 1720 28632 1748
rect 25740 1708 25746 1720
rect 28626 1708 28632 1720
rect 28684 1708 28690 1760
rect 29546 1748 29552 1760
rect 29507 1720 29552 1748
rect 29546 1708 29552 1720
rect 29604 1708 29610 1760
rect 30006 1708 30012 1760
rect 30064 1748 30070 1760
rect 43530 1748 43536 1760
rect 30064 1720 43536 1748
rect 30064 1708 30070 1720
rect 43530 1708 43536 1720
rect 43588 1708 43594 1760
rect 12342 1640 12348 1692
rect 12400 1680 12406 1692
rect 13354 1680 13360 1692
rect 12400 1652 13360 1680
rect 12400 1640 12406 1652
rect 13354 1640 13360 1652
rect 13412 1640 13418 1692
rect 14274 1640 14280 1692
rect 14332 1680 14338 1692
rect 14734 1680 14740 1692
rect 14332 1652 14740 1680
rect 14332 1640 14338 1652
rect 14734 1640 14740 1652
rect 14792 1640 14798 1692
rect 24486 1640 24492 1692
rect 24544 1680 24550 1692
rect 30929 1683 30987 1689
rect 30929 1680 30941 1683
rect 24544 1652 30941 1680
rect 24544 1640 24550 1652
rect 30929 1649 30941 1652
rect 30975 1649 30987 1683
rect 31110 1680 31116 1692
rect 31071 1652 31116 1680
rect 30929 1643 30987 1649
rect 31110 1640 31116 1652
rect 31168 1640 31174 1692
rect 31294 1680 31300 1692
rect 31255 1652 31300 1680
rect 31294 1640 31300 1652
rect 31352 1640 31358 1692
rect 31570 1680 31576 1692
rect 31531 1652 31576 1680
rect 31570 1640 31576 1652
rect 31628 1640 31634 1692
rect 34238 1640 34244 1692
rect 34296 1680 34302 1692
rect 43714 1680 43720 1692
rect 34296 1652 43720 1680
rect 34296 1640 34302 1652
rect 43714 1640 43720 1652
rect 43772 1640 43778 1692
rect 28350 1572 28356 1624
rect 28408 1612 28414 1624
rect 36541 1615 36599 1621
rect 36541 1612 36553 1615
rect 28408 1584 36553 1612
rect 28408 1572 28414 1584
rect 36541 1581 36553 1584
rect 36587 1581 36599 1615
rect 36541 1575 36599 1581
rect 8846 1504 8852 1556
rect 8904 1544 8910 1556
rect 9306 1544 9312 1556
rect 8904 1516 9312 1544
rect 8904 1504 8910 1516
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 13538 1504 13544 1556
rect 13596 1544 13602 1556
rect 13722 1544 13728 1556
rect 13596 1516 13728 1544
rect 13596 1504 13602 1516
rect 13722 1504 13728 1516
rect 13780 1504 13786 1556
rect 29454 1544 29460 1556
rect 29415 1516 29460 1544
rect 29454 1504 29460 1516
rect 29512 1504 29518 1556
rect 30282 1544 30288 1556
rect 30243 1516 30288 1544
rect 30282 1504 30288 1516
rect 30340 1504 30346 1556
rect 30558 1544 30564 1556
rect 30519 1516 30564 1544
rect 30558 1504 30564 1516
rect 30616 1504 30622 1556
rect 30834 1544 30840 1556
rect 30795 1516 30840 1544
rect 30834 1504 30840 1516
rect 30892 1504 30898 1556
rect 31386 1504 31392 1556
rect 31444 1544 31450 1556
rect 31481 1547 31539 1553
rect 31481 1544 31493 1547
rect 31444 1516 31493 1544
rect 31444 1504 31450 1516
rect 31481 1513 31493 1516
rect 31527 1513 31539 1547
rect 31481 1507 31539 1513
rect 4338 1436 4344 1488
rect 4396 1476 4402 1488
rect 4982 1476 4988 1488
rect 4396 1448 4988 1476
rect 4396 1436 4402 1448
rect 4982 1436 4988 1448
rect 5040 1436 5046 1488
rect 14734 1436 14740 1488
rect 14792 1476 14798 1488
rect 15746 1476 15752 1488
rect 14792 1448 15752 1476
rect 14792 1436 14798 1448
rect 15746 1436 15752 1448
rect 15804 1436 15810 1488
rect 22462 1476 22468 1488
rect 22423 1448 22468 1476
rect 22462 1436 22468 1448
rect 22520 1436 22526 1488
rect 24946 1436 24952 1488
rect 25004 1476 25010 1488
rect 25222 1476 25228 1488
rect 25004 1448 25228 1476
rect 25004 1436 25010 1448
rect 25222 1436 25228 1448
rect 25280 1436 25286 1488
rect 27062 1436 27068 1488
rect 27120 1476 27126 1488
rect 36449 1479 36507 1485
rect 36449 1476 36461 1479
rect 27120 1448 36461 1476
rect 27120 1436 27126 1448
rect 36449 1445 36461 1448
rect 36495 1445 36507 1479
rect 36449 1439 36507 1445
rect 4246 1368 4252 1420
rect 4304 1408 4310 1420
rect 4798 1408 4804 1420
rect 4304 1380 4804 1408
rect 4304 1368 4310 1380
rect 4798 1368 4804 1380
rect 4856 1368 4862 1420
rect 8386 1368 8392 1420
rect 8444 1408 8450 1420
rect 8754 1408 8760 1420
rect 8444 1380 8760 1408
rect 8444 1368 8450 1380
rect 8754 1368 8760 1380
rect 8812 1368 8818 1420
rect 10502 1368 10508 1420
rect 10560 1408 10566 1420
rect 16114 1408 16120 1420
rect 10560 1380 16120 1408
rect 10560 1368 10566 1380
rect 16114 1368 16120 1380
rect 16172 1368 16178 1420
rect 16574 1368 16580 1420
rect 16632 1408 16638 1420
rect 17034 1408 17040 1420
rect 16632 1380 17040 1408
rect 16632 1368 16638 1380
rect 17034 1368 17040 1380
rect 17092 1368 17098 1420
rect 18230 1368 18236 1420
rect 18288 1408 18294 1420
rect 19150 1408 19156 1420
rect 18288 1380 19156 1408
rect 18288 1368 18294 1380
rect 19150 1368 19156 1380
rect 19208 1368 19214 1420
rect 19886 1368 19892 1420
rect 19944 1408 19950 1420
rect 20530 1408 20536 1420
rect 19944 1380 20536 1408
rect 19944 1368 19950 1380
rect 20530 1368 20536 1380
rect 20588 1368 20594 1420
rect 25682 1408 25688 1420
rect 24964 1380 25688 1408
rect 24964 1352 24992 1380
rect 25682 1368 25688 1380
rect 25740 1368 25746 1420
rect 29730 1368 29736 1420
rect 29788 1408 29794 1420
rect 31662 1408 31668 1420
rect 29788 1380 31668 1408
rect 29788 1368 29794 1380
rect 31662 1368 31668 1380
rect 31720 1368 31726 1420
rect 32766 1408 32772 1420
rect 32600 1380 32772 1408
rect 32600 1352 32628 1380
rect 32766 1368 32772 1380
rect 32824 1368 32830 1420
rect 38102 1368 38108 1420
rect 38160 1408 38166 1420
rect 38470 1408 38476 1420
rect 38160 1380 38476 1408
rect 38160 1368 38166 1380
rect 38470 1368 38476 1380
rect 38528 1368 38534 1420
rect 40034 1368 40040 1420
rect 40092 1408 40098 1420
rect 41138 1408 41144 1420
rect 40092 1380 41144 1408
rect 40092 1368 40098 1380
rect 41138 1368 41144 1380
rect 41196 1368 41202 1420
rect 44450 1368 44456 1420
rect 44508 1408 44514 1420
rect 48222 1408 48228 1420
rect 44508 1380 48228 1408
rect 44508 1368 44514 1380
rect 48222 1368 48228 1380
rect 48280 1368 48286 1420
rect 49694 1368 49700 1420
rect 49752 1408 49758 1420
rect 50154 1408 50160 1420
rect 49752 1380 50160 1408
rect 49752 1368 49758 1380
rect 50154 1368 50160 1380
rect 50212 1368 50218 1420
rect 55214 1368 55220 1420
rect 55272 1408 55278 1420
rect 55582 1408 55588 1420
rect 55272 1380 55588 1408
rect 55272 1368 55278 1380
rect 55582 1368 55588 1380
rect 55640 1368 55646 1420
rect 61470 1408 61476 1420
rect 59832 1380 61476 1408
rect 15010 1300 15016 1352
rect 15068 1340 15074 1352
rect 15654 1340 15660 1352
rect 15068 1312 15660 1340
rect 15068 1300 15074 1312
rect 15654 1300 15660 1312
rect 15712 1300 15718 1352
rect 24946 1300 24952 1352
rect 25004 1300 25010 1352
rect 30466 1340 30472 1352
rect 30427 1312 30472 1340
rect 30466 1300 30472 1312
rect 30524 1300 30530 1352
rect 30742 1340 30748 1352
rect 30703 1312 30748 1340
rect 30742 1300 30748 1312
rect 30800 1300 30806 1352
rect 32582 1300 32588 1352
rect 32640 1300 32646 1352
rect 32950 1300 32956 1352
rect 33008 1340 33014 1352
rect 35989 1343 36047 1349
rect 35989 1340 36001 1343
rect 33008 1312 36001 1340
rect 33008 1300 33014 1312
rect 35989 1309 36001 1312
rect 36035 1309 36047 1343
rect 35989 1303 36047 1309
rect 58986 1300 58992 1352
rect 59044 1340 59050 1352
rect 59170 1340 59176 1352
rect 59044 1312 59176 1340
rect 59044 1300 59050 1312
rect 59170 1300 59176 1312
rect 59228 1300 59234 1352
rect 4798 1232 4804 1284
rect 4856 1272 4862 1284
rect 5166 1272 5172 1284
rect 4856 1244 5172 1272
rect 4856 1232 4862 1244
rect 5166 1232 5172 1244
rect 5224 1232 5230 1284
rect 33870 1232 33876 1284
rect 33928 1272 33934 1284
rect 34333 1275 34391 1281
rect 34333 1272 34345 1275
rect 33928 1244 34345 1272
rect 33928 1232 33934 1244
rect 34333 1241 34345 1244
rect 34379 1241 34391 1275
rect 34333 1235 34391 1241
rect 40586 1232 40592 1284
rect 40644 1272 40650 1284
rect 40770 1272 40776 1284
rect 40644 1244 40776 1272
rect 40644 1232 40650 1244
rect 40770 1232 40776 1244
rect 40828 1232 40834 1284
rect 50154 1232 50160 1284
rect 50212 1272 50218 1284
rect 50798 1272 50804 1284
rect 50212 1244 50804 1272
rect 50212 1232 50218 1244
rect 50798 1232 50804 1244
rect 50856 1232 50862 1284
rect 11422 1164 11428 1216
rect 11480 1204 11486 1216
rect 12250 1204 12256 1216
rect 11480 1176 12256 1204
rect 11480 1164 11486 1176
rect 12250 1164 12256 1176
rect 12308 1164 12314 1216
rect 15654 1164 15660 1216
rect 15712 1204 15718 1216
rect 16482 1204 16488 1216
rect 15712 1176 16488 1204
rect 15712 1164 15718 1176
rect 16482 1164 16488 1176
rect 16540 1164 16546 1216
rect 44634 1164 44640 1216
rect 44692 1204 44698 1216
rect 45370 1204 45376 1216
rect 44692 1176 45376 1204
rect 44692 1164 44698 1176
rect 45370 1164 45376 1176
rect 45428 1164 45434 1216
rect 48314 1164 48320 1216
rect 48372 1204 48378 1216
rect 52178 1204 52184 1216
rect 48372 1176 52184 1204
rect 48372 1164 48378 1176
rect 52178 1164 52184 1176
rect 52236 1164 52242 1216
rect 11054 1096 11060 1148
rect 11112 1136 11118 1148
rect 12802 1136 12808 1148
rect 11112 1108 12808 1136
rect 11112 1096 11118 1108
rect 12802 1096 12808 1108
rect 12860 1096 12866 1148
rect 36078 1096 36084 1148
rect 36136 1096 36142 1148
rect 33962 960 33968 1012
rect 34020 1000 34026 1012
rect 34057 1003 34115 1009
rect 34057 1000 34069 1003
rect 34020 972 34069 1000
rect 34020 960 34026 972
rect 34057 969 34069 972
rect 34103 969 34115 1003
rect 34057 963 34115 969
rect 36096 944 36124 1096
rect 59832 1080 59860 1380
rect 61470 1368 61476 1380
rect 61528 1368 61534 1420
rect 61930 1368 61936 1420
rect 61988 1408 61994 1420
rect 63402 1408 63408 1420
rect 61988 1380 63408 1408
rect 61988 1368 61994 1380
rect 63402 1368 63408 1380
rect 63460 1368 63466 1420
rect 66806 1368 66812 1420
rect 66864 1408 66870 1420
rect 67266 1408 67272 1420
rect 66864 1380 67272 1408
rect 66864 1368 66870 1380
rect 67266 1368 67272 1380
rect 67324 1368 67330 1420
rect 64414 1232 64420 1284
rect 64472 1272 64478 1284
rect 64690 1272 64696 1284
rect 64472 1244 64696 1272
rect 64472 1232 64478 1244
rect 64690 1232 64696 1244
rect 64748 1232 64754 1284
rect 39758 1068 39764 1080
rect 39719 1040 39764 1068
rect 39758 1028 39764 1040
rect 39816 1028 39822 1080
rect 59814 1028 59820 1080
rect 59872 1028 59878 1080
rect 48682 960 48688 1012
rect 48740 1000 48746 1012
rect 48958 1000 48964 1012
rect 48740 972 48964 1000
rect 48740 960 48746 972
rect 48958 960 48964 972
rect 49016 960 49022 1012
rect 36078 892 36084 944
rect 36136 892 36142 944
rect 53926 892 53932 944
rect 53984 932 53990 944
rect 55030 932 55036 944
rect 53984 904 55036 932
rect 53984 892 53990 904
rect 55030 892 55036 904
rect 55088 892 55094 944
<< via1 >>
rect 4246 67430 4298 67482
rect 4310 67430 4362 67482
rect 4374 67430 4426 67482
rect 4438 67430 4490 67482
rect 14246 67430 14298 67482
rect 14310 67430 14362 67482
rect 14374 67430 14426 67482
rect 14438 67430 14490 67482
rect 24246 67430 24298 67482
rect 24310 67430 24362 67482
rect 24374 67430 24426 67482
rect 24438 67430 24490 67482
rect 34246 67430 34298 67482
rect 34310 67430 34362 67482
rect 34374 67430 34426 67482
rect 34438 67430 34490 67482
rect 44246 67430 44298 67482
rect 44310 67430 44362 67482
rect 44374 67430 44426 67482
rect 44438 67430 44490 67482
rect 54246 67430 54298 67482
rect 54310 67430 54362 67482
rect 54374 67430 54426 67482
rect 54438 67430 54490 67482
rect 64246 67430 64298 67482
rect 64310 67430 64362 67482
rect 64374 67430 64426 67482
rect 64438 67430 64490 67482
rect 16488 67371 16540 67380
rect 16488 67337 16497 67371
rect 16497 67337 16531 67371
rect 16531 67337 16540 67371
rect 16488 67328 16540 67337
rect 940 67260 992 67312
rect 2872 67303 2924 67312
rect 2872 67269 2881 67303
rect 2881 67269 2915 67303
rect 2915 67269 2924 67303
rect 2872 67260 2924 67269
rect 8668 67303 8720 67312
rect 8668 67269 8677 67303
rect 8677 67269 8711 67303
rect 8711 67269 8720 67303
rect 8668 67260 8720 67269
rect 10600 67303 10652 67312
rect 10600 67269 10609 67303
rect 10609 67269 10643 67303
rect 10643 67269 10652 67303
rect 10600 67260 10652 67269
rect 18420 67303 18472 67312
rect 18420 67269 18429 67303
rect 18429 67269 18463 67303
rect 18463 67269 18472 67303
rect 18420 67260 18472 67269
rect 24124 67260 24176 67312
rect 26148 67303 26200 67312
rect 26148 67269 26157 67303
rect 26157 67269 26191 67303
rect 26191 67269 26200 67303
rect 26148 67260 26200 67269
rect 32036 67303 32088 67312
rect 32036 67269 32045 67303
rect 32045 67269 32079 67303
rect 32079 67269 32088 67303
rect 32036 67260 32088 67269
rect 33968 67303 34020 67312
rect 33968 67269 33977 67303
rect 33977 67269 34011 67303
rect 34011 67269 34020 67303
rect 33968 67260 34020 67269
rect 39764 67303 39816 67312
rect 39764 67269 39773 67303
rect 39773 67269 39807 67303
rect 39807 67269 39816 67303
rect 39764 67260 39816 67269
rect 41696 67303 41748 67312
rect 41696 67269 41705 67303
rect 41705 67269 41739 67303
rect 41739 67269 41748 67303
rect 41696 67260 41748 67269
rect 47584 67303 47636 67312
rect 47584 67269 47593 67303
rect 47593 67269 47627 67303
rect 47627 67269 47636 67303
rect 47584 67260 47636 67269
rect 49516 67260 49568 67312
rect 55312 67303 55364 67312
rect 55312 67269 55321 67303
rect 55321 67269 55355 67303
rect 55355 67269 55364 67303
rect 55312 67260 55364 67269
rect 57336 67260 57388 67312
rect 63132 67303 63184 67312
rect 63132 67269 63141 67303
rect 63141 67269 63175 67303
rect 63175 67269 63184 67303
rect 63132 67260 63184 67269
rect 65064 67260 65116 67312
rect 67364 67303 67416 67312
rect 67364 67269 67373 67303
rect 67373 67269 67407 67303
rect 67407 67269 67416 67303
rect 67364 67260 67416 67269
rect 4804 67124 4856 67176
rect 12532 67124 12584 67176
rect 20352 67124 20404 67176
rect 26976 67124 27028 67176
rect 28080 67124 28132 67176
rect 35900 67124 35952 67176
rect 43720 67124 43772 67176
rect 51448 67124 51500 67176
rect 59360 67167 59412 67176
rect 59360 67133 59369 67167
rect 59369 67133 59403 67167
rect 59403 67133 59412 67167
rect 59360 67124 59412 67133
rect 64788 67124 64840 67176
rect 3976 67056 4028 67108
rect 3884 67031 3936 67040
rect 3884 66997 3893 67031
rect 3893 66997 3927 67031
rect 3927 66997 3936 67031
rect 3884 66988 3936 66997
rect 11060 67056 11112 67108
rect 16580 67099 16632 67108
rect 16580 67065 16589 67099
rect 16589 67065 16623 67099
rect 16623 67065 16632 67099
rect 16580 67056 16632 67065
rect 11704 66988 11756 67040
rect 19064 66988 19116 67040
rect 25596 67031 25648 67040
rect 25596 66997 25605 67031
rect 25605 66997 25639 67031
rect 25639 66997 25648 67031
rect 34152 67099 34204 67108
rect 34152 67065 34161 67099
rect 34161 67065 34195 67099
rect 34195 67065 34204 67099
rect 34152 67056 34204 67065
rect 33232 67031 33284 67040
rect 25596 66988 25648 66997
rect 33232 66997 33241 67031
rect 33241 66997 33275 67031
rect 33275 66997 33284 67031
rect 33232 66988 33284 66997
rect 36544 66988 36596 67040
rect 41512 67056 41564 67108
rect 47768 67099 47820 67108
rect 47768 67065 47777 67099
rect 47777 67065 47811 67099
rect 47811 67065 47820 67099
rect 47768 67056 47820 67065
rect 50804 66988 50856 67040
rect 54760 67031 54812 67040
rect 54760 66997 54769 67031
rect 54769 66997 54803 67031
rect 54803 66997 54812 67031
rect 57796 67099 57848 67108
rect 57796 67065 57805 67099
rect 57805 67065 57839 67099
rect 57839 67065 57848 67099
rect 57796 67056 57848 67065
rect 62580 67031 62632 67040
rect 54760 66988 54812 66997
rect 62580 66997 62589 67031
rect 62589 66997 62623 67031
rect 62623 66997 62632 67031
rect 62580 66988 62632 66997
rect 64604 66988 64656 67040
rect 66996 67124 67048 67176
rect 9246 66886 9298 66938
rect 9310 66886 9362 66938
rect 9374 66886 9426 66938
rect 9438 66886 9490 66938
rect 19246 66886 19298 66938
rect 19310 66886 19362 66938
rect 19374 66886 19426 66938
rect 19438 66886 19490 66938
rect 29246 66886 29298 66938
rect 29310 66886 29362 66938
rect 29374 66886 29426 66938
rect 29438 66886 29490 66938
rect 39246 66886 39298 66938
rect 39310 66886 39362 66938
rect 39374 66886 39426 66938
rect 39438 66886 39490 66938
rect 49246 66886 49298 66938
rect 49310 66886 49362 66938
rect 49374 66886 49426 66938
rect 49438 66886 49490 66938
rect 59246 66886 59298 66938
rect 59310 66886 59362 66938
rect 59374 66886 59426 66938
rect 59438 66886 59490 66938
rect 13544 66784 13596 66836
rect 34152 66784 34204 66836
rect 47768 66784 47820 66836
rect 56508 66784 56560 66836
rect 66996 66784 67048 66836
rect 67548 66784 67600 66836
rect 1768 66759 1820 66768
rect 1768 66725 1777 66759
rect 1777 66725 1811 66759
rect 1811 66725 1820 66759
rect 1768 66716 1820 66725
rect 1952 66691 2004 66700
rect 1952 66657 1961 66691
rect 1961 66657 1995 66691
rect 1995 66657 2004 66691
rect 1952 66648 2004 66657
rect 2780 66648 2832 66700
rect 10140 66648 10192 66700
rect 57796 66648 57848 66700
rect 66352 66648 66404 66700
rect 3884 66580 3936 66632
rect 18052 66580 18104 66632
rect 26884 66580 26936 66632
rect 62580 66580 62632 66632
rect 3976 66487 4028 66496
rect 3976 66453 3985 66487
rect 3985 66453 4019 66487
rect 4019 66453 4028 66487
rect 3976 66444 4028 66453
rect 11060 66487 11112 66496
rect 11060 66453 11069 66487
rect 11069 66453 11103 66487
rect 11103 66453 11112 66487
rect 11060 66444 11112 66453
rect 30472 66487 30524 66496
rect 30472 66453 30481 66487
rect 30481 66453 30515 66487
rect 30515 66453 30524 66487
rect 30472 66444 30524 66453
rect 41512 66487 41564 66496
rect 41512 66453 41521 66487
rect 41521 66453 41555 66487
rect 41555 66453 41564 66487
rect 41512 66444 41564 66453
rect 65708 66444 65760 66496
rect 66076 66444 66128 66496
rect 4246 66342 4298 66394
rect 4310 66342 4362 66394
rect 4374 66342 4426 66394
rect 4438 66342 4490 66394
rect 14246 66342 14298 66394
rect 14310 66342 14362 66394
rect 14374 66342 14426 66394
rect 14438 66342 14490 66394
rect 24246 66342 24298 66394
rect 24310 66342 24362 66394
rect 24374 66342 24426 66394
rect 24438 66342 24490 66394
rect 34246 66342 34298 66394
rect 34310 66342 34362 66394
rect 34374 66342 34426 66394
rect 34438 66342 34490 66394
rect 44246 66342 44298 66394
rect 44310 66342 44362 66394
rect 44374 66342 44426 66394
rect 44438 66342 44490 66394
rect 54246 66342 54298 66394
rect 54310 66342 54362 66394
rect 54374 66342 54426 66394
rect 54438 66342 54490 66394
rect 64246 66342 64298 66394
rect 64310 66342 64362 66394
rect 64374 66342 64426 66394
rect 64438 66342 64490 66394
rect 11060 66240 11112 66292
rect 61476 66240 61528 66292
rect 1952 66104 2004 66156
rect 4252 66036 4304 66088
rect 14556 66036 14608 66088
rect 30288 66036 30340 66088
rect 30196 65900 30248 65952
rect 65524 66104 65576 66156
rect 36176 66079 36228 66088
rect 36176 66045 36185 66079
rect 36185 66045 36219 66079
rect 36219 66045 36228 66079
rect 36176 66036 36228 66045
rect 36452 66079 36504 66088
rect 36452 66045 36461 66079
rect 36461 66045 36495 66079
rect 36495 66045 36504 66079
rect 36452 66036 36504 66045
rect 65800 66079 65852 66088
rect 65800 66045 65809 66079
rect 65809 66045 65843 66079
rect 65843 66045 65852 66079
rect 65800 66036 65852 66045
rect 64696 66011 64748 66020
rect 64696 65977 64705 66011
rect 64705 65977 64739 66011
rect 64739 65977 64748 66011
rect 66076 66036 66128 66088
rect 68100 66079 68152 66088
rect 68100 66045 68109 66079
rect 68109 66045 68143 66079
rect 68143 66045 68152 66079
rect 68100 66036 68152 66045
rect 64696 65968 64748 65977
rect 34888 65943 34940 65952
rect 34888 65909 34897 65943
rect 34897 65909 34931 65943
rect 34931 65909 34940 65943
rect 34888 65900 34940 65909
rect 36176 65900 36228 65952
rect 36912 65943 36964 65952
rect 36912 65909 36921 65943
rect 36921 65909 36955 65943
rect 36955 65909 36964 65943
rect 36912 65900 36964 65909
rect 66720 65943 66772 65952
rect 66720 65909 66729 65943
rect 66729 65909 66763 65943
rect 66763 65909 66772 65943
rect 66720 65900 66772 65909
rect 9246 65798 9298 65850
rect 9310 65798 9362 65850
rect 9374 65798 9426 65850
rect 9438 65798 9490 65850
rect 19246 65798 19298 65850
rect 19310 65798 19362 65850
rect 19374 65798 19426 65850
rect 19438 65798 19490 65850
rect 29246 65798 29298 65850
rect 29310 65798 29362 65850
rect 29374 65798 29426 65850
rect 29438 65798 29490 65850
rect 39246 65798 39298 65850
rect 39310 65798 39362 65850
rect 39374 65798 39426 65850
rect 39438 65798 39490 65850
rect 49246 65798 49298 65850
rect 49310 65798 49362 65850
rect 49374 65798 49426 65850
rect 49438 65798 49490 65850
rect 59246 65798 59298 65850
rect 59310 65798 59362 65850
rect 59374 65798 59426 65850
rect 59438 65798 59490 65850
rect 16672 65696 16724 65748
rect 30196 65696 30248 65748
rect 30288 65696 30340 65748
rect 37924 65696 37976 65748
rect 65524 65739 65576 65748
rect 65524 65705 65533 65739
rect 65533 65705 65567 65739
rect 65567 65705 65576 65739
rect 65524 65696 65576 65705
rect 68100 65739 68152 65748
rect 68100 65705 68109 65739
rect 68109 65705 68143 65739
rect 68143 65705 68152 65739
rect 68100 65696 68152 65705
rect 1860 65399 1912 65408
rect 1860 65365 1869 65399
rect 1869 65365 1903 65399
rect 1903 65365 1912 65399
rect 1860 65356 1912 65365
rect 4620 65560 4672 65612
rect 66720 65560 66772 65612
rect 4252 65492 4304 65544
rect 67640 65492 67692 65544
rect 19064 65424 19116 65476
rect 2688 65356 2740 65408
rect 23020 65399 23072 65408
rect 23020 65365 23029 65399
rect 23029 65365 23063 65399
rect 23063 65365 23072 65399
rect 23020 65356 23072 65365
rect 56784 65356 56836 65408
rect 65432 65356 65484 65408
rect 66168 65356 66220 65408
rect 4246 65254 4298 65306
rect 4310 65254 4362 65306
rect 4374 65254 4426 65306
rect 4438 65254 4490 65306
rect 14246 65254 14298 65306
rect 14310 65254 14362 65306
rect 14374 65254 14426 65306
rect 14438 65254 14490 65306
rect 24246 65254 24298 65306
rect 24310 65254 24362 65306
rect 24374 65254 24426 65306
rect 24438 65254 24490 65306
rect 34246 65254 34298 65306
rect 34310 65254 34362 65306
rect 34374 65254 34426 65306
rect 34438 65254 34490 65306
rect 44246 65254 44298 65306
rect 44310 65254 44362 65306
rect 44374 65254 44426 65306
rect 44438 65254 44490 65306
rect 54246 65254 54298 65306
rect 54310 65254 54362 65306
rect 54374 65254 54426 65306
rect 54438 65254 54490 65306
rect 64246 65254 64298 65306
rect 64310 65254 64362 65306
rect 64374 65254 64426 65306
rect 64438 65254 64490 65306
rect 23020 65084 23072 65136
rect 67180 65084 67232 65136
rect 66168 65016 66220 65068
rect 17132 64948 17184 65000
rect 55220 64948 55272 65000
rect 66812 64948 66864 65000
rect 66260 64880 66312 64932
rect 67824 64880 67876 64932
rect 67640 64855 67692 64864
rect 67640 64821 67649 64855
rect 67649 64821 67683 64855
rect 67683 64821 67692 64855
rect 67640 64812 67692 64821
rect 9246 64710 9298 64762
rect 9310 64710 9362 64762
rect 9374 64710 9426 64762
rect 9438 64710 9490 64762
rect 19246 64710 19298 64762
rect 19310 64710 19362 64762
rect 19374 64710 19426 64762
rect 19438 64710 19490 64762
rect 29246 64710 29298 64762
rect 29310 64710 29362 64762
rect 29374 64710 29426 64762
rect 29438 64710 29490 64762
rect 39246 64710 39298 64762
rect 39310 64710 39362 64762
rect 39374 64710 39426 64762
rect 39438 64710 39490 64762
rect 49246 64710 49298 64762
rect 49310 64710 49362 64762
rect 49374 64710 49426 64762
rect 49438 64710 49490 64762
rect 59246 64710 59298 64762
rect 59310 64710 59362 64762
rect 59374 64710 59426 64762
rect 59438 64710 59490 64762
rect 27528 64336 27580 64388
rect 64696 64336 64748 64388
rect 2228 64311 2280 64320
rect 2228 64277 2237 64311
rect 2237 64277 2271 64311
rect 2271 64277 2280 64311
rect 2228 64268 2280 64277
rect 6736 64268 6788 64320
rect 66168 64268 66220 64320
rect 67640 64268 67692 64320
rect 4246 64166 4298 64218
rect 4310 64166 4362 64218
rect 4374 64166 4426 64218
rect 4438 64166 4490 64218
rect 14246 64166 14298 64218
rect 14310 64166 14362 64218
rect 14374 64166 14426 64218
rect 14438 64166 14490 64218
rect 24246 64166 24298 64218
rect 24310 64166 24362 64218
rect 24374 64166 24426 64218
rect 24438 64166 24490 64218
rect 34246 64166 34298 64218
rect 34310 64166 34362 64218
rect 34374 64166 34426 64218
rect 34438 64166 34490 64218
rect 44246 64166 44298 64218
rect 44310 64166 44362 64218
rect 44374 64166 44426 64218
rect 44438 64166 44490 64218
rect 54246 64166 54298 64218
rect 54310 64166 54362 64218
rect 54374 64166 54426 64218
rect 54438 64166 54490 64218
rect 64246 64166 64298 64218
rect 64310 64166 64362 64218
rect 64374 64166 64426 64218
rect 64438 64166 64490 64218
rect 2228 64064 2280 64116
rect 38108 64064 38160 64116
rect 16672 63996 16724 64048
rect 68100 63971 68152 63980
rect 68100 63937 68109 63971
rect 68109 63937 68143 63971
rect 68143 63937 68152 63971
rect 68100 63928 68152 63937
rect 14004 63903 14056 63912
rect 14004 63869 14013 63903
rect 14013 63869 14047 63903
rect 14047 63869 14056 63903
rect 14004 63860 14056 63869
rect 12900 63767 12952 63776
rect 12900 63733 12909 63767
rect 12909 63733 12943 63767
rect 12943 63733 12952 63767
rect 12900 63724 12952 63733
rect 67272 63767 67324 63776
rect 67272 63733 67281 63767
rect 67281 63733 67315 63767
rect 67315 63733 67324 63767
rect 67272 63724 67324 63733
rect 9246 63622 9298 63674
rect 9310 63622 9362 63674
rect 9374 63622 9426 63674
rect 9438 63622 9490 63674
rect 19246 63622 19298 63674
rect 19310 63622 19362 63674
rect 19374 63622 19426 63674
rect 19438 63622 19490 63674
rect 29246 63622 29298 63674
rect 29310 63622 29362 63674
rect 29374 63622 29426 63674
rect 29438 63622 29490 63674
rect 39246 63622 39298 63674
rect 39310 63622 39362 63674
rect 39374 63622 39426 63674
rect 39438 63622 39490 63674
rect 49246 63622 49298 63674
rect 49310 63622 49362 63674
rect 49374 63622 49426 63674
rect 49438 63622 49490 63674
rect 59246 63622 59298 63674
rect 59310 63622 59362 63674
rect 59374 63622 59426 63674
rect 59438 63622 59490 63674
rect 12900 63520 12952 63572
rect 27528 63520 27580 63572
rect 12716 63384 12768 63436
rect 13176 63316 13228 63368
rect 12716 63223 12768 63232
rect 12716 63189 12725 63223
rect 12725 63189 12759 63223
rect 12759 63189 12768 63223
rect 12716 63180 12768 63189
rect 13176 63223 13228 63232
rect 13176 63189 13185 63223
rect 13185 63189 13219 63223
rect 13219 63189 13228 63223
rect 13176 63180 13228 63189
rect 32404 63180 32456 63232
rect 50068 63180 50120 63232
rect 66628 63180 66680 63232
rect 68100 63291 68152 63300
rect 68100 63257 68109 63291
rect 68109 63257 68143 63291
rect 68143 63257 68152 63291
rect 68100 63248 68152 63257
rect 4246 63078 4298 63130
rect 4310 63078 4362 63130
rect 4374 63078 4426 63130
rect 4438 63078 4490 63130
rect 14246 63078 14298 63130
rect 14310 63078 14362 63130
rect 14374 63078 14426 63130
rect 14438 63078 14490 63130
rect 24246 63078 24298 63130
rect 24310 63078 24362 63130
rect 24374 63078 24426 63130
rect 24438 63078 24490 63130
rect 34246 63078 34298 63130
rect 34310 63078 34362 63130
rect 34374 63078 34426 63130
rect 34438 63078 34490 63130
rect 44246 63078 44298 63130
rect 44310 63078 44362 63130
rect 44374 63078 44426 63130
rect 44438 63078 44490 63130
rect 54246 63078 54298 63130
rect 54310 63078 54362 63130
rect 54374 63078 54426 63130
rect 54438 63078 54490 63130
rect 64246 63078 64298 63130
rect 64310 63078 64362 63130
rect 64374 63078 64426 63130
rect 64438 63078 64490 63130
rect 12716 62976 12768 63028
rect 19984 62976 20036 63028
rect 62764 62976 62816 63028
rect 2044 62908 2096 62960
rect 36452 62908 36504 62960
rect 48964 62908 49016 62960
rect 3976 62840 4028 62892
rect 1584 62815 1636 62824
rect 1584 62781 1593 62815
rect 1593 62781 1627 62815
rect 1627 62781 1636 62815
rect 1584 62772 1636 62781
rect 9772 62815 9824 62824
rect 9772 62781 9781 62815
rect 9781 62781 9815 62815
rect 9815 62781 9824 62815
rect 9772 62772 9824 62781
rect 49148 62772 49200 62824
rect 66904 62772 66956 62824
rect 17776 62636 17828 62688
rect 50068 62704 50120 62756
rect 51448 62636 51500 62688
rect 66536 62679 66588 62688
rect 66536 62645 66545 62679
rect 66545 62645 66579 62679
rect 66579 62645 66588 62679
rect 66536 62636 66588 62645
rect 9246 62534 9298 62586
rect 9310 62534 9362 62586
rect 9374 62534 9426 62586
rect 9438 62534 9490 62586
rect 19246 62534 19298 62586
rect 19310 62534 19362 62586
rect 19374 62534 19426 62586
rect 19438 62534 19490 62586
rect 29246 62534 29298 62586
rect 29310 62534 29362 62586
rect 29374 62534 29426 62586
rect 29438 62534 29490 62586
rect 39246 62534 39298 62586
rect 39310 62534 39362 62586
rect 39374 62534 39426 62586
rect 39438 62534 39490 62586
rect 49246 62534 49298 62586
rect 49310 62534 49362 62586
rect 49374 62534 49426 62586
rect 49438 62534 49490 62586
rect 59246 62534 59298 62586
rect 59310 62534 59362 62586
rect 59374 62534 59426 62586
rect 59438 62534 59490 62586
rect 9772 62432 9824 62484
rect 64696 62432 64748 62484
rect 65064 62432 65116 62484
rect 66904 62475 66956 62484
rect 66904 62441 66913 62475
rect 66913 62441 66947 62475
rect 66947 62441 66956 62475
rect 66904 62432 66956 62441
rect 48964 62407 49016 62416
rect 48964 62373 48973 62407
rect 48973 62373 49007 62407
rect 49007 62373 49016 62407
rect 48964 62364 49016 62373
rect 49608 62364 49660 62416
rect 66536 62364 66588 62416
rect 32496 62228 32548 62280
rect 33140 62160 33192 62212
rect 55036 62092 55088 62144
rect 4246 61990 4298 62042
rect 4310 61990 4362 62042
rect 4374 61990 4426 62042
rect 4438 61990 4490 62042
rect 14246 61990 14298 62042
rect 14310 61990 14362 62042
rect 14374 61990 14426 62042
rect 14438 61990 14490 62042
rect 24246 61990 24298 62042
rect 24310 61990 24362 62042
rect 24374 61990 24426 62042
rect 24438 61990 24490 62042
rect 34246 61990 34298 62042
rect 34310 61990 34362 62042
rect 34374 61990 34426 62042
rect 34438 61990 34490 62042
rect 44246 61990 44298 62042
rect 44310 61990 44362 62042
rect 44374 61990 44426 62042
rect 44438 61990 44490 62042
rect 54246 61990 54298 62042
rect 54310 61990 54362 62042
rect 54374 61990 54426 62042
rect 54438 61990 54490 62042
rect 64246 61990 64298 62042
rect 64310 61990 64362 62042
rect 64374 61990 64426 62042
rect 64438 61990 64490 62042
rect 67272 61820 67324 61872
rect 67272 61684 67324 61736
rect 1860 61591 1912 61600
rect 1860 61557 1869 61591
rect 1869 61557 1903 61591
rect 1903 61557 1912 61591
rect 1860 61548 1912 61557
rect 2320 61548 2372 61600
rect 9246 61446 9298 61498
rect 9310 61446 9362 61498
rect 9374 61446 9426 61498
rect 9438 61446 9490 61498
rect 19246 61446 19298 61498
rect 19310 61446 19362 61498
rect 19374 61446 19426 61498
rect 19438 61446 19490 61498
rect 29246 61446 29298 61498
rect 29310 61446 29362 61498
rect 29374 61446 29426 61498
rect 29438 61446 29490 61498
rect 39246 61446 39298 61498
rect 39310 61446 39362 61498
rect 39374 61446 39426 61498
rect 39438 61446 39490 61498
rect 49246 61446 49298 61498
rect 49310 61446 49362 61498
rect 49374 61446 49426 61498
rect 49438 61446 49490 61498
rect 59246 61446 59298 61498
rect 59310 61446 59362 61498
rect 59374 61446 59426 61498
rect 59438 61446 59490 61498
rect 68100 61251 68152 61260
rect 68100 61217 68109 61251
rect 68109 61217 68143 61251
rect 68143 61217 68152 61251
rect 68100 61208 68152 61217
rect 4246 60902 4298 60954
rect 4310 60902 4362 60954
rect 4374 60902 4426 60954
rect 4438 60902 4490 60954
rect 14246 60902 14298 60954
rect 14310 60902 14362 60954
rect 14374 60902 14426 60954
rect 14438 60902 14490 60954
rect 24246 60902 24298 60954
rect 24310 60902 24362 60954
rect 24374 60902 24426 60954
rect 24438 60902 24490 60954
rect 34246 60902 34298 60954
rect 34310 60902 34362 60954
rect 34374 60902 34426 60954
rect 34438 60902 34490 60954
rect 44246 60902 44298 60954
rect 44310 60902 44362 60954
rect 44374 60902 44426 60954
rect 44438 60902 44490 60954
rect 54246 60902 54298 60954
rect 54310 60902 54362 60954
rect 54374 60902 54426 60954
rect 54438 60902 54490 60954
rect 64246 60902 64298 60954
rect 64310 60902 64362 60954
rect 64374 60902 64426 60954
rect 64438 60902 64490 60954
rect 51448 60707 51500 60716
rect 51448 60673 51457 60707
rect 51457 60673 51491 60707
rect 51491 60673 51500 60707
rect 51448 60664 51500 60673
rect 9246 60358 9298 60410
rect 9310 60358 9362 60410
rect 9374 60358 9426 60410
rect 9438 60358 9490 60410
rect 19246 60358 19298 60410
rect 19310 60358 19362 60410
rect 19374 60358 19426 60410
rect 19438 60358 19490 60410
rect 29246 60358 29298 60410
rect 29310 60358 29362 60410
rect 29374 60358 29426 60410
rect 29438 60358 29490 60410
rect 39246 60358 39298 60410
rect 39310 60358 39362 60410
rect 39374 60358 39426 60410
rect 39438 60358 39490 60410
rect 49246 60358 49298 60410
rect 49310 60358 49362 60410
rect 49374 60358 49426 60410
rect 49438 60358 49490 60410
rect 59246 60358 59298 60410
rect 59310 60358 59362 60410
rect 59374 60358 59426 60410
rect 59438 60358 59490 60410
rect 51448 60188 51500 60240
rect 1768 60163 1820 60172
rect 1768 60129 1777 60163
rect 1777 60129 1811 60163
rect 1811 60129 1820 60163
rect 1768 60120 1820 60129
rect 1860 60120 1912 60172
rect 50988 60120 51040 60172
rect 52368 60163 52420 60172
rect 52368 60129 52377 60163
rect 52377 60129 52411 60163
rect 52411 60129 52420 60163
rect 52368 60120 52420 60129
rect 2136 60052 2188 60104
rect 44088 60052 44140 60104
rect 49608 60052 49660 60104
rect 51632 60052 51684 60104
rect 56508 60120 56560 60172
rect 58624 60052 58676 60104
rect 30288 59984 30340 60036
rect 66812 59984 66864 60036
rect 2596 59916 2648 59968
rect 47400 59959 47452 59968
rect 47400 59925 47409 59959
rect 47409 59925 47443 59959
rect 47443 59925 47452 59959
rect 47400 59916 47452 59925
rect 50436 59916 50488 59968
rect 50988 59916 51040 59968
rect 52092 59959 52144 59968
rect 52092 59925 52101 59959
rect 52101 59925 52135 59959
rect 52135 59925 52144 59959
rect 52092 59916 52144 59925
rect 53196 59959 53248 59968
rect 53196 59925 53205 59959
rect 53205 59925 53239 59959
rect 53239 59925 53248 59959
rect 53196 59916 53248 59925
rect 4246 59814 4298 59866
rect 4310 59814 4362 59866
rect 4374 59814 4426 59866
rect 4438 59814 4490 59866
rect 14246 59814 14298 59866
rect 14310 59814 14362 59866
rect 14374 59814 14426 59866
rect 14438 59814 14490 59866
rect 24246 59814 24298 59866
rect 24310 59814 24362 59866
rect 24374 59814 24426 59866
rect 24438 59814 24490 59866
rect 34246 59814 34298 59866
rect 34310 59814 34362 59866
rect 34374 59814 34426 59866
rect 34438 59814 34490 59866
rect 44246 59814 44298 59866
rect 44310 59814 44362 59866
rect 44374 59814 44426 59866
rect 44438 59814 44490 59866
rect 54246 59814 54298 59866
rect 54310 59814 54362 59866
rect 54374 59814 54426 59866
rect 54438 59814 54490 59866
rect 64246 59814 64298 59866
rect 64310 59814 64362 59866
rect 64374 59814 64426 59866
rect 64438 59814 64490 59866
rect 14832 59576 14884 59628
rect 66260 59576 66312 59628
rect 16672 59508 16724 59560
rect 17224 59508 17276 59560
rect 66720 59508 66772 59560
rect 33508 59440 33560 59492
rect 14832 59415 14884 59424
rect 14832 59381 14841 59415
rect 14841 59381 14875 59415
rect 14875 59381 14884 59415
rect 14832 59372 14884 59381
rect 17224 59372 17276 59424
rect 51632 59415 51684 59424
rect 51632 59381 51641 59415
rect 51641 59381 51675 59415
rect 51675 59381 51684 59415
rect 51632 59372 51684 59381
rect 52368 59372 52420 59424
rect 58716 59372 58768 59424
rect 9246 59270 9298 59322
rect 9310 59270 9362 59322
rect 9374 59270 9426 59322
rect 9438 59270 9490 59322
rect 19246 59270 19298 59322
rect 19310 59270 19362 59322
rect 19374 59270 19426 59322
rect 19438 59270 19490 59322
rect 29246 59270 29298 59322
rect 29310 59270 29362 59322
rect 29374 59270 29426 59322
rect 29438 59270 29490 59322
rect 39246 59270 39298 59322
rect 39310 59270 39362 59322
rect 39374 59270 39426 59322
rect 39438 59270 39490 59322
rect 49246 59270 49298 59322
rect 49310 59270 49362 59322
rect 49374 59270 49426 59322
rect 49438 59270 49490 59322
rect 59246 59270 59298 59322
rect 59310 59270 59362 59322
rect 59374 59270 59426 59322
rect 59438 59270 59490 59322
rect 66628 58964 66680 59016
rect 33140 58896 33192 58948
rect 33416 58896 33468 58948
rect 43996 58896 44048 58948
rect 13452 58871 13504 58880
rect 13452 58837 13461 58871
rect 13461 58837 13495 58871
rect 13495 58837 13504 58871
rect 13452 58828 13504 58837
rect 64144 58828 64196 58880
rect 4246 58726 4298 58778
rect 4310 58726 4362 58778
rect 4374 58726 4426 58778
rect 4438 58726 4490 58778
rect 14246 58726 14298 58778
rect 14310 58726 14362 58778
rect 14374 58726 14426 58778
rect 14438 58726 14490 58778
rect 24246 58726 24298 58778
rect 24310 58726 24362 58778
rect 24374 58726 24426 58778
rect 24438 58726 24490 58778
rect 34246 58726 34298 58778
rect 34310 58726 34362 58778
rect 34374 58726 34426 58778
rect 34438 58726 34490 58778
rect 44246 58726 44298 58778
rect 44310 58726 44362 58778
rect 44374 58726 44426 58778
rect 44438 58726 44490 58778
rect 54246 58726 54298 58778
rect 54310 58726 54362 58778
rect 54374 58726 54426 58778
rect 54438 58726 54490 58778
rect 64246 58726 64298 58778
rect 64310 58726 64362 58778
rect 64374 58726 64426 58778
rect 64438 58726 64490 58778
rect 8208 58624 8260 58676
rect 29092 58624 29144 58676
rect 30288 58624 30340 58676
rect 42524 58624 42576 58676
rect 3884 58556 3936 58608
rect 44180 58556 44232 58608
rect 2688 58488 2740 58540
rect 43996 58531 44048 58540
rect 43996 58497 44005 58531
rect 44005 58497 44039 58531
rect 44039 58497 44048 58531
rect 43996 58488 44048 58497
rect 44088 58531 44140 58540
rect 44088 58497 44097 58531
rect 44097 58497 44131 58531
rect 44131 58497 44140 58531
rect 44456 58556 44508 58608
rect 68100 58599 68152 58608
rect 68100 58565 68109 58599
rect 68109 58565 68143 58599
rect 68143 58565 68152 58599
rect 68100 58556 68152 58565
rect 44088 58488 44140 58497
rect 27988 58463 28040 58472
rect 27988 58429 27997 58463
rect 27997 58429 28031 58463
rect 28031 58429 28040 58463
rect 27988 58420 28040 58429
rect 34520 58463 34572 58472
rect 34520 58429 34529 58463
rect 34529 58429 34563 58463
rect 34563 58429 34572 58463
rect 34520 58420 34572 58429
rect 43260 58420 43312 58472
rect 67364 58352 67416 58404
rect 42524 58327 42576 58336
rect 42524 58293 42533 58327
rect 42533 58293 42567 58327
rect 42567 58293 42576 58327
rect 42524 58284 42576 58293
rect 43260 58327 43312 58336
rect 43260 58293 43269 58327
rect 43269 58293 43303 58327
rect 43303 58293 43312 58327
rect 43260 58284 43312 58293
rect 43812 58327 43864 58336
rect 43812 58293 43821 58327
rect 43821 58293 43855 58327
rect 43855 58293 43864 58327
rect 43812 58284 43864 58293
rect 66996 58284 67048 58336
rect 9246 58182 9298 58234
rect 9310 58182 9362 58234
rect 9374 58182 9426 58234
rect 9438 58182 9490 58234
rect 19246 58182 19298 58234
rect 19310 58182 19362 58234
rect 19374 58182 19426 58234
rect 19438 58182 19490 58234
rect 29246 58182 29298 58234
rect 29310 58182 29362 58234
rect 29374 58182 29426 58234
rect 29438 58182 29490 58234
rect 39246 58182 39298 58234
rect 39310 58182 39362 58234
rect 39374 58182 39426 58234
rect 39438 58182 39490 58234
rect 49246 58182 49298 58234
rect 49310 58182 49362 58234
rect 49374 58182 49426 58234
rect 49438 58182 49490 58234
rect 59246 58182 59298 58234
rect 59310 58182 59362 58234
rect 59374 58182 59426 58234
rect 59438 58182 59490 58234
rect 6920 58080 6972 58132
rect 8208 58080 8260 58132
rect 34520 58080 34572 58132
rect 46848 58080 46900 58132
rect 65524 58055 65576 58064
rect 4712 57944 4764 57996
rect 6920 57944 6972 57996
rect 6368 57919 6420 57928
rect 6368 57885 6377 57919
rect 6377 57885 6411 57919
rect 6411 57885 6420 57919
rect 6368 57876 6420 57885
rect 65524 58021 65533 58055
rect 65533 58021 65567 58055
rect 65567 58021 65576 58055
rect 65524 58012 65576 58021
rect 27988 57944 28040 57996
rect 48872 57944 48924 57996
rect 65064 57987 65116 57996
rect 65064 57953 65073 57987
rect 65073 57953 65107 57987
rect 65107 57953 65116 57987
rect 65064 57944 65116 57953
rect 50252 57876 50304 57928
rect 4712 57783 4764 57792
rect 4712 57749 4721 57783
rect 4721 57749 4755 57783
rect 4755 57749 4764 57783
rect 4712 57740 4764 57749
rect 8208 57783 8260 57792
rect 8208 57749 8217 57783
rect 8217 57749 8251 57783
rect 8251 57749 8260 57783
rect 8208 57740 8260 57749
rect 26976 57808 27028 57860
rect 27804 57740 27856 57792
rect 36176 57783 36228 57792
rect 36176 57749 36185 57783
rect 36185 57749 36219 57783
rect 36219 57749 36228 57783
rect 36176 57740 36228 57749
rect 43444 57783 43496 57792
rect 43444 57749 43453 57783
rect 43453 57749 43487 57783
rect 43487 57749 43496 57783
rect 43444 57740 43496 57749
rect 44088 57740 44140 57792
rect 45284 57783 45336 57792
rect 45284 57749 45293 57783
rect 45293 57749 45327 57783
rect 45327 57749 45336 57783
rect 45284 57740 45336 57749
rect 55128 57783 55180 57792
rect 55128 57749 55137 57783
rect 55137 57749 55171 57783
rect 55171 57749 55180 57783
rect 55128 57740 55180 57749
rect 58624 57740 58676 57792
rect 65064 57740 65116 57792
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 14246 57638 14298 57690
rect 14310 57638 14362 57690
rect 14374 57638 14426 57690
rect 14438 57638 14490 57690
rect 24246 57638 24298 57690
rect 24310 57638 24362 57690
rect 24374 57638 24426 57690
rect 24438 57638 24490 57690
rect 34246 57638 34298 57690
rect 34310 57638 34362 57690
rect 34374 57638 34426 57690
rect 34438 57638 34490 57690
rect 44246 57638 44298 57690
rect 44310 57638 44362 57690
rect 44374 57638 44426 57690
rect 44438 57638 44490 57690
rect 54246 57638 54298 57690
rect 54310 57638 54362 57690
rect 54374 57638 54426 57690
rect 54438 57638 54490 57690
rect 64246 57638 64298 57690
rect 64310 57638 64362 57690
rect 64374 57638 64426 57690
rect 64438 57638 64490 57690
rect 8208 57536 8260 57588
rect 44916 57536 44968 57588
rect 45284 57536 45336 57588
rect 63960 57536 64012 57588
rect 67272 57579 67324 57588
rect 67272 57545 67281 57579
rect 67281 57545 67315 57579
rect 67315 57545 67324 57579
rect 67272 57536 67324 57545
rect 11704 57468 11756 57520
rect 36176 57468 36228 57520
rect 51448 57468 51500 57520
rect 8852 57400 8904 57452
rect 1584 57375 1636 57384
rect 1584 57341 1593 57375
rect 1593 57341 1627 57375
rect 1627 57341 1636 57375
rect 1584 57332 1636 57341
rect 25504 57375 25556 57384
rect 25504 57341 25513 57375
rect 25513 57341 25547 57375
rect 25547 57341 25556 57375
rect 25504 57332 25556 57341
rect 67272 57332 67324 57384
rect 68100 57307 68152 57316
rect 68100 57273 68109 57307
rect 68109 57273 68143 57307
rect 68143 57273 68152 57307
rect 68100 57264 68152 57273
rect 6368 57196 6420 57248
rect 18328 57196 18380 57248
rect 50252 57196 50304 57248
rect 66168 57196 66220 57248
rect 9246 57094 9298 57146
rect 9310 57094 9362 57146
rect 9374 57094 9426 57146
rect 9438 57094 9490 57146
rect 19246 57094 19298 57146
rect 19310 57094 19362 57146
rect 19374 57094 19426 57146
rect 19438 57094 19490 57146
rect 29246 57094 29298 57146
rect 29310 57094 29362 57146
rect 29374 57094 29426 57146
rect 29438 57094 29490 57146
rect 39246 57094 39298 57146
rect 39310 57094 39362 57146
rect 39374 57094 39426 57146
rect 39438 57094 39490 57146
rect 49246 57094 49298 57146
rect 49310 57094 49362 57146
rect 49374 57094 49426 57146
rect 49438 57094 49490 57146
rect 59246 57094 59298 57146
rect 59310 57094 59362 57146
rect 59374 57094 59426 57146
rect 59438 57094 59490 57146
rect 12624 56652 12676 56704
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 14246 56550 14298 56602
rect 14310 56550 14362 56602
rect 14374 56550 14426 56602
rect 14438 56550 14490 56602
rect 24246 56550 24298 56602
rect 24310 56550 24362 56602
rect 24374 56550 24426 56602
rect 24438 56550 24490 56602
rect 34246 56550 34298 56602
rect 34310 56550 34362 56602
rect 34374 56550 34426 56602
rect 34438 56550 34490 56602
rect 44246 56550 44298 56602
rect 44310 56550 44362 56602
rect 44374 56550 44426 56602
rect 44438 56550 44490 56602
rect 54246 56550 54298 56602
rect 54310 56550 54362 56602
rect 54374 56550 54426 56602
rect 54438 56550 54490 56602
rect 64246 56550 64298 56602
rect 64310 56550 64362 56602
rect 64374 56550 64426 56602
rect 64438 56550 64490 56602
rect 1768 56355 1820 56364
rect 1768 56321 1777 56355
rect 1777 56321 1811 56355
rect 1811 56321 1820 56355
rect 1768 56312 1820 56321
rect 30288 56287 30340 56296
rect 30288 56253 30297 56287
rect 30297 56253 30331 56287
rect 30331 56253 30340 56287
rect 30288 56244 30340 56253
rect 44640 56244 44692 56296
rect 68100 56287 68152 56296
rect 68100 56253 68109 56287
rect 68109 56253 68143 56287
rect 68143 56253 68152 56287
rect 68100 56244 68152 56253
rect 2504 56151 2556 56160
rect 2504 56117 2513 56151
rect 2513 56117 2547 56151
rect 2547 56117 2556 56151
rect 2504 56108 2556 56117
rect 9246 56006 9298 56058
rect 9310 56006 9362 56058
rect 9374 56006 9426 56058
rect 9438 56006 9490 56058
rect 19246 56006 19298 56058
rect 19310 56006 19362 56058
rect 19374 56006 19426 56058
rect 19438 56006 19490 56058
rect 29246 56006 29298 56058
rect 29310 56006 29362 56058
rect 29374 56006 29426 56058
rect 29438 56006 29490 56058
rect 39246 56006 39298 56058
rect 39310 56006 39362 56058
rect 39374 56006 39426 56058
rect 39438 56006 39490 56058
rect 49246 56006 49298 56058
rect 49310 56006 49362 56058
rect 49374 56006 49426 56058
rect 49438 56006 49490 56058
rect 59246 56006 59298 56058
rect 59310 56006 59362 56058
rect 59374 56006 59426 56058
rect 59438 56006 59490 56058
rect 2688 55632 2740 55684
rect 9956 55811 10008 55820
rect 9956 55777 9965 55811
rect 9965 55777 9999 55811
rect 9999 55777 10008 55811
rect 9956 55768 10008 55777
rect 11060 55607 11112 55616
rect 11060 55573 11069 55607
rect 11069 55573 11103 55607
rect 11103 55573 11112 55607
rect 11060 55564 11112 55573
rect 13084 55607 13136 55616
rect 13084 55573 13093 55607
rect 13093 55573 13127 55607
rect 13127 55573 13136 55607
rect 13084 55564 13136 55573
rect 31300 55836 31352 55888
rect 51632 55836 51684 55888
rect 25504 55632 25556 55684
rect 47584 55632 47636 55684
rect 38016 55607 38068 55616
rect 38016 55573 38025 55607
rect 38025 55573 38059 55607
rect 38059 55573 38068 55607
rect 38016 55564 38068 55573
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 14246 55462 14298 55514
rect 14310 55462 14362 55514
rect 14374 55462 14426 55514
rect 14438 55462 14490 55514
rect 24246 55462 24298 55514
rect 24310 55462 24362 55514
rect 24374 55462 24426 55514
rect 24438 55462 24490 55514
rect 34246 55462 34298 55514
rect 34310 55462 34362 55514
rect 34374 55462 34426 55514
rect 34438 55462 34490 55514
rect 44246 55462 44298 55514
rect 44310 55462 44362 55514
rect 44374 55462 44426 55514
rect 44438 55462 44490 55514
rect 54246 55462 54298 55514
rect 54310 55462 54362 55514
rect 54374 55462 54426 55514
rect 54438 55462 54490 55514
rect 64246 55462 64298 55514
rect 64310 55462 64362 55514
rect 64374 55462 64426 55514
rect 64438 55462 64490 55514
rect 11060 55360 11112 55412
rect 42340 55360 42392 55412
rect 9956 55292 10008 55344
rect 31300 55292 31352 55344
rect 39948 55292 40000 55344
rect 67456 55292 67508 55344
rect 2688 55224 2740 55276
rect 38016 55156 38068 55208
rect 38752 55156 38804 55208
rect 37464 55088 37516 55140
rect 41696 55224 41748 55276
rect 67088 55224 67140 55276
rect 1860 55063 1912 55072
rect 1860 55029 1869 55063
rect 1869 55029 1903 55063
rect 1903 55029 1912 55063
rect 1860 55020 1912 55029
rect 38384 55063 38436 55072
rect 38384 55029 38393 55063
rect 38393 55029 38427 55063
rect 38427 55029 38436 55063
rect 38384 55020 38436 55029
rect 62764 55020 62816 55072
rect 9246 54918 9298 54970
rect 9310 54918 9362 54970
rect 9374 54918 9426 54970
rect 9438 54918 9490 54970
rect 19246 54918 19298 54970
rect 19310 54918 19362 54970
rect 19374 54918 19426 54970
rect 19438 54918 19490 54970
rect 29246 54918 29298 54970
rect 29310 54918 29362 54970
rect 29374 54918 29426 54970
rect 29438 54918 29490 54970
rect 39246 54918 39298 54970
rect 39310 54918 39362 54970
rect 39374 54918 39426 54970
rect 39438 54918 39490 54970
rect 49246 54918 49298 54970
rect 49310 54918 49362 54970
rect 49374 54918 49426 54970
rect 49438 54918 49490 54970
rect 59246 54918 59298 54970
rect 59310 54918 59362 54970
rect 59374 54918 59426 54970
rect 59438 54918 59490 54970
rect 33876 54476 33928 54528
rect 38752 54476 38804 54528
rect 44824 54519 44876 54528
rect 44824 54485 44833 54519
rect 44833 54485 44867 54519
rect 44867 54485 44876 54519
rect 44824 54476 44876 54485
rect 62120 54519 62172 54528
rect 62120 54485 62129 54519
rect 62129 54485 62163 54519
rect 62163 54485 62172 54519
rect 62120 54476 62172 54485
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 14246 54374 14298 54426
rect 14310 54374 14362 54426
rect 14374 54374 14426 54426
rect 14438 54374 14490 54426
rect 24246 54374 24298 54426
rect 24310 54374 24362 54426
rect 24374 54374 24426 54426
rect 24438 54374 24490 54426
rect 34246 54374 34298 54426
rect 34310 54374 34362 54426
rect 34374 54374 34426 54426
rect 34438 54374 34490 54426
rect 44246 54374 44298 54426
rect 44310 54374 44362 54426
rect 44374 54374 44426 54426
rect 44438 54374 44490 54426
rect 54246 54374 54298 54426
rect 54310 54374 54362 54426
rect 54374 54374 54426 54426
rect 54438 54374 54490 54426
rect 64246 54374 64298 54426
rect 64310 54374 64362 54426
rect 64374 54374 64426 54426
rect 64438 54374 64490 54426
rect 2412 54272 2464 54324
rect 44824 54272 44876 54324
rect 48780 54111 48832 54120
rect 48780 54077 48789 54111
rect 48789 54077 48823 54111
rect 48823 54077 48832 54111
rect 48780 54068 48832 54077
rect 66904 54068 66956 54120
rect 9246 53830 9298 53882
rect 9310 53830 9362 53882
rect 9374 53830 9426 53882
rect 9438 53830 9490 53882
rect 19246 53830 19298 53882
rect 19310 53830 19362 53882
rect 19374 53830 19426 53882
rect 19438 53830 19490 53882
rect 29246 53830 29298 53882
rect 29310 53830 29362 53882
rect 29374 53830 29426 53882
rect 29438 53830 29490 53882
rect 39246 53830 39298 53882
rect 39310 53830 39362 53882
rect 39374 53830 39426 53882
rect 39438 53830 39490 53882
rect 49246 53830 49298 53882
rect 49310 53830 49362 53882
rect 49374 53830 49426 53882
rect 49438 53830 49490 53882
rect 59246 53830 59298 53882
rect 59310 53830 59362 53882
rect 59374 53830 59426 53882
rect 59438 53830 59490 53882
rect 37464 53728 37516 53780
rect 12164 53388 12216 53440
rect 19984 53388 20036 53440
rect 29092 53524 29144 53576
rect 29552 53524 29604 53576
rect 32864 53567 32916 53576
rect 32864 53533 32873 53567
rect 32873 53533 32907 53567
rect 32907 53533 32916 53567
rect 32864 53524 32916 53533
rect 33140 53567 33192 53576
rect 33140 53533 33149 53567
rect 33149 53533 33183 53567
rect 33183 53533 33192 53567
rect 33140 53524 33192 53533
rect 43260 53592 43312 53644
rect 37188 53388 37240 53440
rect 43444 53388 43496 53440
rect 53932 53431 53984 53440
rect 53932 53397 53941 53431
rect 53941 53397 53975 53431
rect 53975 53397 53984 53431
rect 53932 53388 53984 53397
rect 55588 53388 55640 53440
rect 55864 53388 55916 53440
rect 68100 53499 68152 53508
rect 68100 53465 68109 53499
rect 68109 53465 68143 53499
rect 68143 53465 68152 53499
rect 68100 53456 68152 53465
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 14246 53286 14298 53338
rect 14310 53286 14362 53338
rect 14374 53286 14426 53338
rect 14438 53286 14490 53338
rect 24246 53286 24298 53338
rect 24310 53286 24362 53338
rect 24374 53286 24426 53338
rect 24438 53286 24490 53338
rect 34246 53286 34298 53338
rect 34310 53286 34362 53338
rect 34374 53286 34426 53338
rect 34438 53286 34490 53338
rect 44246 53286 44298 53338
rect 44310 53286 44362 53338
rect 44374 53286 44426 53338
rect 44438 53286 44490 53338
rect 54246 53286 54298 53338
rect 54310 53286 54362 53338
rect 54374 53286 54426 53338
rect 54438 53286 54490 53338
rect 64246 53286 64298 53338
rect 64310 53286 64362 53338
rect 64374 53286 64426 53338
rect 64438 53286 64490 53338
rect 2688 53184 2740 53236
rect 53932 53116 53984 53168
rect 66352 53048 66404 53100
rect 45100 52980 45152 53032
rect 52000 52980 52052 53032
rect 53012 52980 53064 53032
rect 54576 53023 54628 53032
rect 54576 52989 54585 53023
rect 54585 52989 54619 53023
rect 54619 52989 54628 53023
rect 54576 52980 54628 52989
rect 54668 52980 54720 53032
rect 55588 53023 55640 53032
rect 32864 52912 32916 52964
rect 36912 52912 36964 52964
rect 33140 52844 33192 52896
rect 53012 52887 53064 52896
rect 53012 52853 53021 52887
rect 53021 52853 53055 52887
rect 53055 52853 53064 52887
rect 53012 52844 53064 52853
rect 53840 52887 53892 52896
rect 53840 52853 53849 52887
rect 53849 52853 53883 52887
rect 53883 52853 53892 52887
rect 55588 52989 55597 53023
rect 55597 52989 55631 53023
rect 55631 52989 55640 53023
rect 55588 52980 55640 52989
rect 62856 53023 62908 53032
rect 62856 52989 62865 53023
rect 62865 52989 62899 53023
rect 62899 52989 62908 53023
rect 62856 52980 62908 52989
rect 65248 53023 65300 53032
rect 65248 52989 65257 53023
rect 65257 52989 65291 53023
rect 65291 52989 65300 53023
rect 65248 52980 65300 52989
rect 62764 52955 62816 52964
rect 62764 52921 62773 52955
rect 62773 52921 62807 52955
rect 62807 52921 62816 52955
rect 62764 52912 62816 52921
rect 53840 52844 53892 52853
rect 9246 52742 9298 52794
rect 9310 52742 9362 52794
rect 9374 52742 9426 52794
rect 9438 52742 9490 52794
rect 19246 52742 19298 52794
rect 19310 52742 19362 52794
rect 19374 52742 19426 52794
rect 19438 52742 19490 52794
rect 29246 52742 29298 52794
rect 29310 52742 29362 52794
rect 29374 52742 29426 52794
rect 29438 52742 29490 52794
rect 39246 52742 39298 52794
rect 39310 52742 39362 52794
rect 39374 52742 39426 52794
rect 39438 52742 39490 52794
rect 49246 52742 49298 52794
rect 49310 52742 49362 52794
rect 49374 52742 49426 52794
rect 49438 52742 49490 52794
rect 59246 52742 59298 52794
rect 59310 52742 59362 52794
rect 59374 52742 59426 52794
rect 59438 52742 59490 52794
rect 39948 52640 40000 52692
rect 48228 52640 48280 52692
rect 55588 52640 55640 52692
rect 62396 52640 62448 52692
rect 62856 52640 62908 52692
rect 1584 52547 1636 52556
rect 1584 52513 1593 52547
rect 1593 52513 1627 52547
rect 1627 52513 1636 52547
rect 1584 52504 1636 52513
rect 11244 52504 11296 52556
rect 53840 52504 53892 52556
rect 54668 52504 54720 52556
rect 19984 52436 20036 52488
rect 20628 52436 20680 52488
rect 54024 52479 54076 52488
rect 54024 52445 54033 52479
rect 54033 52445 54067 52479
rect 54067 52445 54076 52479
rect 54024 52436 54076 52445
rect 54576 52436 54628 52488
rect 55312 52479 55364 52488
rect 55312 52445 55321 52479
rect 55321 52445 55355 52479
rect 55355 52445 55364 52479
rect 55312 52436 55364 52445
rect 65984 52368 66036 52420
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 14246 52198 14298 52250
rect 14310 52198 14362 52250
rect 14374 52198 14426 52250
rect 14438 52198 14490 52250
rect 24246 52198 24298 52250
rect 24310 52198 24362 52250
rect 24374 52198 24426 52250
rect 24438 52198 24490 52250
rect 34246 52198 34298 52250
rect 34310 52198 34362 52250
rect 34374 52198 34426 52250
rect 34438 52198 34490 52250
rect 44246 52198 44298 52250
rect 44310 52198 44362 52250
rect 44374 52198 44426 52250
rect 44438 52198 44490 52250
rect 54246 52198 54298 52250
rect 54310 52198 54362 52250
rect 54374 52198 54426 52250
rect 54438 52198 54490 52250
rect 64246 52198 64298 52250
rect 64310 52198 64362 52250
rect 64374 52198 64426 52250
rect 64438 52198 64490 52250
rect 67180 52096 67232 52148
rect 15844 51935 15896 51944
rect 15844 51901 15853 51935
rect 15853 51901 15887 51935
rect 15887 51901 15896 51935
rect 15844 51892 15896 51901
rect 68100 52003 68152 52012
rect 68100 51969 68109 52003
rect 68109 51969 68143 52003
rect 68143 51969 68152 52003
rect 68100 51960 68152 51969
rect 31300 51756 31352 51808
rect 32036 51756 32088 51808
rect 53932 51756 53984 51808
rect 9246 51654 9298 51706
rect 9310 51654 9362 51706
rect 9374 51654 9426 51706
rect 9438 51654 9490 51706
rect 19246 51654 19298 51706
rect 19310 51654 19362 51706
rect 19374 51654 19426 51706
rect 19438 51654 19490 51706
rect 29246 51654 29298 51706
rect 29310 51654 29362 51706
rect 29374 51654 29426 51706
rect 29438 51654 29490 51706
rect 39246 51654 39298 51706
rect 39310 51654 39362 51706
rect 39374 51654 39426 51706
rect 39438 51654 39490 51706
rect 49246 51654 49298 51706
rect 49310 51654 49362 51706
rect 49374 51654 49426 51706
rect 49438 51654 49490 51706
rect 59246 51654 59298 51706
rect 59310 51654 59362 51706
rect 59374 51654 59426 51706
rect 59438 51654 59490 51706
rect 39948 51416 40000 51468
rect 31300 51348 31352 51400
rect 46204 51391 46256 51400
rect 46204 51357 46213 51391
rect 46213 51357 46247 51391
rect 46247 51357 46256 51391
rect 46204 51348 46256 51357
rect 2504 51212 2556 51264
rect 66444 51280 66496 51332
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 14246 51110 14298 51162
rect 14310 51110 14362 51162
rect 14374 51110 14426 51162
rect 14438 51110 14490 51162
rect 24246 51110 24298 51162
rect 24310 51110 24362 51162
rect 24374 51110 24426 51162
rect 24438 51110 24490 51162
rect 34246 51110 34298 51162
rect 34310 51110 34362 51162
rect 34374 51110 34426 51162
rect 34438 51110 34490 51162
rect 44246 51110 44298 51162
rect 44310 51110 44362 51162
rect 44374 51110 44426 51162
rect 44438 51110 44490 51162
rect 54246 51110 54298 51162
rect 54310 51110 54362 51162
rect 54374 51110 54426 51162
rect 54438 51110 54490 51162
rect 64246 51110 64298 51162
rect 64310 51110 64362 51162
rect 64374 51110 64426 51162
rect 64438 51110 64490 51162
rect 1860 51051 1912 51060
rect 1860 51017 1869 51051
rect 1869 51017 1903 51051
rect 1903 51017 1912 51051
rect 1860 51008 1912 51017
rect 2688 51008 2740 51060
rect 16580 50872 16632 50924
rect 17868 50736 17920 50788
rect 55956 50804 56008 50856
rect 68100 50847 68152 50856
rect 68100 50813 68109 50847
rect 68109 50813 68143 50847
rect 68143 50813 68152 50847
rect 68100 50804 68152 50813
rect 49608 50668 49660 50720
rect 50436 50668 50488 50720
rect 9246 50566 9298 50618
rect 9310 50566 9362 50618
rect 9374 50566 9426 50618
rect 9438 50566 9490 50618
rect 19246 50566 19298 50618
rect 19310 50566 19362 50618
rect 19374 50566 19426 50618
rect 19438 50566 19490 50618
rect 29246 50566 29298 50618
rect 29310 50566 29362 50618
rect 29374 50566 29426 50618
rect 29438 50566 29490 50618
rect 39246 50566 39298 50618
rect 39310 50566 39362 50618
rect 39374 50566 39426 50618
rect 39438 50566 39490 50618
rect 49246 50566 49298 50618
rect 49310 50566 49362 50618
rect 49374 50566 49426 50618
rect 49438 50566 49490 50618
rect 59246 50566 59298 50618
rect 59310 50566 59362 50618
rect 59374 50566 59426 50618
rect 59438 50566 59490 50618
rect 30932 50328 30984 50380
rect 54024 50328 54076 50380
rect 34152 50192 34204 50244
rect 3148 50167 3200 50176
rect 3148 50133 3157 50167
rect 3157 50133 3191 50167
rect 3191 50133 3200 50167
rect 3148 50124 3200 50133
rect 23296 50167 23348 50176
rect 23296 50133 23305 50167
rect 23305 50133 23339 50167
rect 23339 50133 23348 50167
rect 23296 50124 23348 50133
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 14246 50022 14298 50074
rect 14310 50022 14362 50074
rect 14374 50022 14426 50074
rect 14438 50022 14490 50074
rect 24246 50022 24298 50074
rect 24310 50022 24362 50074
rect 24374 50022 24426 50074
rect 24438 50022 24490 50074
rect 34246 50022 34298 50074
rect 34310 50022 34362 50074
rect 34374 50022 34426 50074
rect 34438 50022 34490 50074
rect 44246 50022 44298 50074
rect 44310 50022 44362 50074
rect 44374 50022 44426 50074
rect 44438 50022 44490 50074
rect 54246 50022 54298 50074
rect 54310 50022 54362 50074
rect 54374 50022 54426 50074
rect 54438 50022 54490 50074
rect 64246 50022 64298 50074
rect 64310 50022 64362 50074
rect 64374 50022 64426 50074
rect 64438 50022 64490 50074
rect 23296 49920 23348 49972
rect 65432 49920 65484 49972
rect 1768 49827 1820 49836
rect 1768 49793 1777 49827
rect 1777 49793 1811 49827
rect 1811 49793 1820 49827
rect 1768 49784 1820 49793
rect 11796 49784 11848 49836
rect 30932 49852 30984 49904
rect 34980 49852 35032 49904
rect 6920 49716 6972 49768
rect 33876 49784 33928 49836
rect 33968 49648 34020 49700
rect 34704 49759 34756 49768
rect 34704 49725 34718 49759
rect 34718 49725 34752 49759
rect 34752 49725 34756 49759
rect 34704 49716 34756 49725
rect 62764 49716 62816 49768
rect 28264 49580 28316 49632
rect 40132 49648 40184 49700
rect 9246 49478 9298 49530
rect 9310 49478 9362 49530
rect 9374 49478 9426 49530
rect 9438 49478 9490 49530
rect 19246 49478 19298 49530
rect 19310 49478 19362 49530
rect 19374 49478 19426 49530
rect 19438 49478 19490 49530
rect 29246 49478 29298 49530
rect 29310 49478 29362 49530
rect 29374 49478 29426 49530
rect 29438 49478 29490 49530
rect 39246 49478 39298 49530
rect 39310 49478 39362 49530
rect 39374 49478 39426 49530
rect 39438 49478 39490 49530
rect 49246 49478 49298 49530
rect 49310 49478 49362 49530
rect 49374 49478 49426 49530
rect 49438 49478 49490 49530
rect 59246 49478 59298 49530
rect 59310 49478 59362 49530
rect 59374 49478 59426 49530
rect 59438 49478 59490 49530
rect 33968 49079 34020 49088
rect 33968 49045 33977 49079
rect 33977 49045 34011 49079
rect 34011 49045 34020 49079
rect 33968 49036 34020 49045
rect 40132 49036 40184 49088
rect 65800 49036 65852 49088
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 14246 48934 14298 48986
rect 14310 48934 14362 48986
rect 14374 48934 14426 48986
rect 14438 48934 14490 48986
rect 24246 48934 24298 48986
rect 24310 48934 24362 48986
rect 24374 48934 24426 48986
rect 24438 48934 24490 48986
rect 34246 48934 34298 48986
rect 34310 48934 34362 48986
rect 34374 48934 34426 48986
rect 34438 48934 34490 48986
rect 44246 48934 44298 48986
rect 44310 48934 44362 48986
rect 44374 48934 44426 48986
rect 44438 48934 44490 48986
rect 54246 48934 54298 48986
rect 54310 48934 54362 48986
rect 54374 48934 54426 48986
rect 54438 48934 54490 48986
rect 64246 48934 64298 48986
rect 64310 48934 64362 48986
rect 64374 48934 64426 48986
rect 64438 48934 64490 48986
rect 9246 48390 9298 48442
rect 9310 48390 9362 48442
rect 9374 48390 9426 48442
rect 9438 48390 9490 48442
rect 19246 48390 19298 48442
rect 19310 48390 19362 48442
rect 19374 48390 19426 48442
rect 19438 48390 19490 48442
rect 29246 48390 29298 48442
rect 29310 48390 29362 48442
rect 29374 48390 29426 48442
rect 29438 48390 29490 48442
rect 39246 48390 39298 48442
rect 39310 48390 39362 48442
rect 39374 48390 39426 48442
rect 39438 48390 39490 48442
rect 49246 48390 49298 48442
rect 49310 48390 49362 48442
rect 49374 48390 49426 48442
rect 49438 48390 49490 48442
rect 59246 48390 59298 48442
rect 59310 48390 59362 48442
rect 59374 48390 59426 48442
rect 59438 48390 59490 48442
rect 26332 48152 26384 48204
rect 27528 48152 27580 48204
rect 66812 48152 66864 48204
rect 68100 48059 68152 48068
rect 68100 48025 68109 48059
rect 68109 48025 68143 48059
rect 68143 48025 68152 48059
rect 68100 48016 68152 48025
rect 45008 47991 45060 48000
rect 45008 47957 45017 47991
rect 45017 47957 45051 47991
rect 45051 47957 45060 47991
rect 45008 47948 45060 47957
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 14246 47846 14298 47898
rect 14310 47846 14362 47898
rect 14374 47846 14426 47898
rect 14438 47846 14490 47898
rect 24246 47846 24298 47898
rect 24310 47846 24362 47898
rect 24374 47846 24426 47898
rect 24438 47846 24490 47898
rect 34246 47846 34298 47898
rect 34310 47846 34362 47898
rect 34374 47846 34426 47898
rect 34438 47846 34490 47898
rect 44246 47846 44298 47898
rect 44310 47846 44362 47898
rect 44374 47846 44426 47898
rect 44438 47846 44490 47898
rect 54246 47846 54298 47898
rect 54310 47846 54362 47898
rect 54374 47846 54426 47898
rect 54438 47846 54490 47898
rect 64246 47846 64298 47898
rect 64310 47846 64362 47898
rect 64374 47846 64426 47898
rect 64438 47846 64490 47898
rect 33232 47608 33284 47660
rect 40408 47608 40460 47660
rect 40316 47540 40368 47592
rect 65340 47540 65392 47592
rect 9246 47302 9298 47354
rect 9310 47302 9362 47354
rect 9374 47302 9426 47354
rect 9438 47302 9490 47354
rect 19246 47302 19298 47354
rect 19310 47302 19362 47354
rect 19374 47302 19426 47354
rect 19438 47302 19490 47354
rect 29246 47302 29298 47354
rect 29310 47302 29362 47354
rect 29374 47302 29426 47354
rect 29438 47302 29490 47354
rect 39246 47302 39298 47354
rect 39310 47302 39362 47354
rect 39374 47302 39426 47354
rect 39438 47302 39490 47354
rect 49246 47302 49298 47354
rect 49310 47302 49362 47354
rect 49374 47302 49426 47354
rect 49438 47302 49490 47354
rect 59246 47302 59298 47354
rect 59310 47302 59362 47354
rect 59374 47302 59426 47354
rect 59438 47302 59490 47354
rect 27528 47200 27580 47252
rect 1860 47175 1912 47184
rect 1860 47141 1869 47175
rect 1869 47141 1903 47175
rect 1903 47141 1912 47175
rect 1860 47132 1912 47141
rect 31668 47132 31720 47184
rect 31852 47132 31904 47184
rect 40776 47132 40828 47184
rect 44824 46996 44876 47048
rect 32588 46971 32640 46980
rect 32588 46937 32597 46971
rect 32597 46937 32631 46971
rect 32631 46937 32640 46971
rect 32588 46928 32640 46937
rect 33968 46928 34020 46980
rect 46756 46928 46808 46980
rect 48688 46928 48740 46980
rect 67180 46928 67232 46980
rect 68100 46971 68152 46980
rect 68100 46937 68109 46971
rect 68109 46937 68143 46971
rect 68143 46937 68152 46971
rect 68100 46928 68152 46937
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 14246 46758 14298 46810
rect 14310 46758 14362 46810
rect 14374 46758 14426 46810
rect 14438 46758 14490 46810
rect 24246 46758 24298 46810
rect 24310 46758 24362 46810
rect 24374 46758 24426 46810
rect 24438 46758 24490 46810
rect 34246 46758 34298 46810
rect 34310 46758 34362 46810
rect 34374 46758 34426 46810
rect 34438 46758 34490 46810
rect 44246 46758 44298 46810
rect 44310 46758 44362 46810
rect 44374 46758 44426 46810
rect 44438 46758 44490 46810
rect 54246 46758 54298 46810
rect 54310 46758 54362 46810
rect 54374 46758 54426 46810
rect 54438 46758 54490 46810
rect 64246 46758 64298 46810
rect 64310 46758 64362 46810
rect 64374 46758 64426 46810
rect 64438 46758 64490 46810
rect 1860 46656 1912 46708
rect 60740 46452 60792 46504
rect 63684 46384 63736 46436
rect 9246 46214 9298 46266
rect 9310 46214 9362 46266
rect 9374 46214 9426 46266
rect 9438 46214 9490 46266
rect 19246 46214 19298 46266
rect 19310 46214 19362 46266
rect 19374 46214 19426 46266
rect 19438 46214 19490 46266
rect 29246 46214 29298 46266
rect 29310 46214 29362 46266
rect 29374 46214 29426 46266
rect 29438 46214 29490 46266
rect 39246 46214 39298 46266
rect 39310 46214 39362 46266
rect 39374 46214 39426 46266
rect 39438 46214 39490 46266
rect 49246 46214 49298 46266
rect 49310 46214 49362 46266
rect 49374 46214 49426 46266
rect 49438 46214 49490 46266
rect 59246 46214 59298 46266
rect 59310 46214 59362 46266
rect 59374 46214 59426 46266
rect 59438 46214 59490 46266
rect 2412 46112 2464 46164
rect 1768 45951 1820 45960
rect 1768 45917 1777 45951
rect 1777 45917 1811 45951
rect 1811 45917 1820 45951
rect 1768 45908 1820 45917
rect 39120 45772 39172 45824
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 14246 45670 14298 45722
rect 14310 45670 14362 45722
rect 14374 45670 14426 45722
rect 14438 45670 14490 45722
rect 24246 45670 24298 45722
rect 24310 45670 24362 45722
rect 24374 45670 24426 45722
rect 24438 45670 24490 45722
rect 34246 45670 34298 45722
rect 34310 45670 34362 45722
rect 34374 45670 34426 45722
rect 34438 45670 34490 45722
rect 44246 45670 44298 45722
rect 44310 45670 44362 45722
rect 44374 45670 44426 45722
rect 44438 45670 44490 45722
rect 54246 45670 54298 45722
rect 54310 45670 54362 45722
rect 54374 45670 54426 45722
rect 54438 45670 54490 45722
rect 64246 45670 64298 45722
rect 64310 45670 64362 45722
rect 64374 45670 64426 45722
rect 64438 45670 64490 45722
rect 39948 45543 40000 45552
rect 39948 45509 39957 45543
rect 39957 45509 39991 45543
rect 39991 45509 40000 45543
rect 39948 45500 40000 45509
rect 58624 45500 58676 45552
rect 12992 45407 13044 45416
rect 12992 45373 13001 45407
rect 13001 45373 13035 45407
rect 13035 45373 13044 45407
rect 12992 45364 13044 45373
rect 40132 45364 40184 45416
rect 40316 45407 40368 45416
rect 40316 45373 40325 45407
rect 40325 45373 40359 45407
rect 40359 45373 40368 45407
rect 40316 45364 40368 45373
rect 39120 45296 39172 45348
rect 39856 45228 39908 45280
rect 65616 45432 65668 45484
rect 68100 45407 68152 45416
rect 68100 45373 68109 45407
rect 68109 45373 68143 45407
rect 68143 45373 68152 45407
rect 68100 45364 68152 45373
rect 9246 45126 9298 45178
rect 9310 45126 9362 45178
rect 9374 45126 9426 45178
rect 9438 45126 9490 45178
rect 19246 45126 19298 45178
rect 19310 45126 19362 45178
rect 19374 45126 19426 45178
rect 19438 45126 19490 45178
rect 29246 45126 29298 45178
rect 29310 45126 29362 45178
rect 29374 45126 29426 45178
rect 29438 45126 29490 45178
rect 39246 45126 39298 45178
rect 39310 45126 39362 45178
rect 39374 45126 39426 45178
rect 39438 45126 39490 45178
rect 49246 45126 49298 45178
rect 49310 45126 49362 45178
rect 49374 45126 49426 45178
rect 49438 45126 49490 45178
rect 59246 45126 59298 45178
rect 59310 45126 59362 45178
rect 59374 45126 59426 45178
rect 59438 45126 59490 45178
rect 12992 45024 13044 45076
rect 66536 45024 66588 45076
rect 2136 44956 2188 45008
rect 13636 44956 13688 45008
rect 7288 44752 7340 44804
rect 1860 44727 1912 44736
rect 1860 44693 1869 44727
rect 1869 44693 1903 44727
rect 1903 44693 1912 44727
rect 1860 44684 1912 44693
rect 7012 44684 7064 44736
rect 17224 44888 17276 44940
rect 17684 44888 17736 44940
rect 17868 44888 17920 44940
rect 21364 44956 21416 45008
rect 30288 44956 30340 45008
rect 58716 44999 58768 45008
rect 58716 44965 58725 44999
rect 58725 44965 58759 44999
rect 58759 44965 58768 44999
rect 58716 44956 58768 44965
rect 34152 44888 34204 44940
rect 58624 44888 58676 44940
rect 58808 44931 58860 44940
rect 58808 44897 58817 44931
rect 58817 44897 58851 44931
rect 58851 44897 58860 44931
rect 58808 44888 58860 44897
rect 17868 44727 17920 44736
rect 17868 44693 17877 44727
rect 17877 44693 17911 44727
rect 17911 44693 17920 44727
rect 17868 44684 17920 44693
rect 40316 44684 40368 44736
rect 49608 44684 49660 44736
rect 60004 44752 60056 44804
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 14246 44582 14298 44634
rect 14310 44582 14362 44634
rect 14374 44582 14426 44634
rect 14438 44582 14490 44634
rect 24246 44582 24298 44634
rect 24310 44582 24362 44634
rect 24374 44582 24426 44634
rect 24438 44582 24490 44634
rect 34246 44582 34298 44634
rect 34310 44582 34362 44634
rect 34374 44582 34426 44634
rect 34438 44582 34490 44634
rect 44246 44582 44298 44634
rect 44310 44582 44362 44634
rect 44374 44582 44426 44634
rect 44438 44582 44490 44634
rect 54246 44582 54298 44634
rect 54310 44582 54362 44634
rect 54374 44582 54426 44634
rect 54438 44582 54490 44634
rect 64246 44582 64298 44634
rect 64310 44582 64362 44634
rect 64374 44582 64426 44634
rect 64438 44582 64490 44634
rect 58808 44480 58860 44532
rect 11704 44344 11756 44396
rect 21364 44344 21416 44396
rect 10692 44319 10744 44328
rect 10692 44285 10701 44319
rect 10701 44285 10735 44319
rect 10735 44285 10744 44319
rect 10692 44276 10744 44285
rect 48964 44208 49016 44260
rect 49608 44208 49660 44260
rect 33140 44140 33192 44192
rect 9246 44038 9298 44090
rect 9310 44038 9362 44090
rect 9374 44038 9426 44090
rect 9438 44038 9490 44090
rect 19246 44038 19298 44090
rect 19310 44038 19362 44090
rect 19374 44038 19426 44090
rect 19438 44038 19490 44090
rect 29246 44038 29298 44090
rect 29310 44038 29362 44090
rect 29374 44038 29426 44090
rect 29438 44038 29490 44090
rect 39246 44038 39298 44090
rect 39310 44038 39362 44090
rect 39374 44038 39426 44090
rect 39438 44038 39490 44090
rect 49246 44038 49298 44090
rect 49310 44038 49362 44090
rect 49374 44038 49426 44090
rect 49438 44038 49490 44090
rect 59246 44038 59298 44090
rect 59310 44038 59362 44090
rect 59374 44038 59426 44090
rect 59438 44038 59490 44090
rect 55312 43936 55364 43988
rect 56048 43936 56100 43988
rect 30564 43800 30616 43852
rect 62396 43843 62448 43852
rect 62396 43809 62405 43843
rect 62405 43809 62439 43843
rect 62439 43809 62448 43843
rect 62396 43800 62448 43809
rect 56048 43732 56100 43784
rect 17868 43596 17920 43648
rect 30748 43596 30800 43648
rect 35716 43639 35768 43648
rect 35716 43605 35725 43639
rect 35725 43605 35759 43639
rect 35759 43605 35768 43639
rect 35716 43596 35768 43605
rect 67548 43596 67600 43648
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 14246 43494 14298 43546
rect 14310 43494 14362 43546
rect 14374 43494 14426 43546
rect 14438 43494 14490 43546
rect 24246 43494 24298 43546
rect 24310 43494 24362 43546
rect 24374 43494 24426 43546
rect 24438 43494 24490 43546
rect 34246 43494 34298 43546
rect 34310 43494 34362 43546
rect 34374 43494 34426 43546
rect 34438 43494 34490 43546
rect 44246 43494 44298 43546
rect 44310 43494 44362 43546
rect 44374 43494 44426 43546
rect 44438 43494 44490 43546
rect 54246 43494 54298 43546
rect 54310 43494 54362 43546
rect 54374 43494 54426 43546
rect 54438 43494 54490 43546
rect 64246 43494 64298 43546
rect 64310 43494 64362 43546
rect 64374 43494 64426 43546
rect 64438 43494 64490 43546
rect 3700 43256 3752 43308
rect 17868 43256 17920 43308
rect 12992 43231 13044 43240
rect 12992 43197 13001 43231
rect 13001 43197 13035 43231
rect 13035 43197 13044 43231
rect 12992 43188 13044 43197
rect 60832 43188 60884 43240
rect 3700 43095 3752 43104
rect 3700 43061 3709 43095
rect 3709 43061 3743 43095
rect 3743 43061 3752 43095
rect 3700 43052 3752 43061
rect 13360 43052 13412 43104
rect 33140 43052 33192 43104
rect 9246 42950 9298 43002
rect 9310 42950 9362 43002
rect 9374 42950 9426 43002
rect 9438 42950 9490 43002
rect 19246 42950 19298 43002
rect 19310 42950 19362 43002
rect 19374 42950 19426 43002
rect 19438 42950 19490 43002
rect 29246 42950 29298 43002
rect 29310 42950 29362 43002
rect 29374 42950 29426 43002
rect 29438 42950 29490 43002
rect 39246 42950 39298 43002
rect 39310 42950 39362 43002
rect 39374 42950 39426 43002
rect 39438 42950 39490 43002
rect 49246 42950 49298 43002
rect 49310 42950 49362 43002
rect 49374 42950 49426 43002
rect 49438 42950 49490 43002
rect 59246 42950 59298 43002
rect 59310 42950 59362 43002
rect 59374 42950 59426 43002
rect 59438 42950 59490 43002
rect 13360 42848 13412 42900
rect 27252 42848 27304 42900
rect 37188 42576 37240 42628
rect 66720 42712 66772 42764
rect 68100 42755 68152 42764
rect 68100 42721 68109 42755
rect 68109 42721 68143 42755
rect 68143 42721 68152 42755
rect 68100 42712 68152 42721
rect 50252 42687 50304 42696
rect 50252 42653 50261 42687
rect 50261 42653 50295 42687
rect 50295 42653 50304 42687
rect 50252 42644 50304 42653
rect 7840 42508 7892 42560
rect 12808 42551 12860 42560
rect 12808 42517 12817 42551
rect 12817 42517 12851 42551
rect 12851 42517 12860 42551
rect 12808 42508 12860 42517
rect 60188 42576 60240 42628
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 14246 42406 14298 42458
rect 14310 42406 14362 42458
rect 14374 42406 14426 42458
rect 14438 42406 14490 42458
rect 24246 42406 24298 42458
rect 24310 42406 24362 42458
rect 24374 42406 24426 42458
rect 24438 42406 24490 42458
rect 34246 42406 34298 42458
rect 34310 42406 34362 42458
rect 34374 42406 34426 42458
rect 34438 42406 34490 42458
rect 44246 42406 44298 42458
rect 44310 42406 44362 42458
rect 44374 42406 44426 42458
rect 44438 42406 44490 42458
rect 54246 42406 54298 42458
rect 54310 42406 54362 42458
rect 54374 42406 54426 42458
rect 54438 42406 54490 42458
rect 64246 42406 64298 42458
rect 64310 42406 64362 42458
rect 64374 42406 64426 42458
rect 64438 42406 64490 42458
rect 12808 42304 12860 42356
rect 49976 42304 50028 42356
rect 18328 42236 18380 42288
rect 22928 42236 22980 42288
rect 1584 42143 1636 42152
rect 1584 42109 1593 42143
rect 1593 42109 1627 42143
rect 1627 42109 1636 42143
rect 1584 42100 1636 42109
rect 51356 42143 51408 42152
rect 51356 42109 51365 42143
rect 51365 42109 51399 42143
rect 51399 42109 51408 42143
rect 51356 42100 51408 42109
rect 65524 42100 65576 42152
rect 22928 42032 22980 42084
rect 39120 42032 39172 42084
rect 21364 41964 21416 42016
rect 53472 41964 53524 42016
rect 9246 41862 9298 41914
rect 9310 41862 9362 41914
rect 9374 41862 9426 41914
rect 9438 41862 9490 41914
rect 19246 41862 19298 41914
rect 19310 41862 19362 41914
rect 19374 41862 19426 41914
rect 19438 41862 19490 41914
rect 29246 41862 29298 41914
rect 29310 41862 29362 41914
rect 29374 41862 29426 41914
rect 29438 41862 29490 41914
rect 39246 41862 39298 41914
rect 39310 41862 39362 41914
rect 39374 41862 39426 41914
rect 39438 41862 39490 41914
rect 49246 41862 49298 41914
rect 49310 41862 49362 41914
rect 49374 41862 49426 41914
rect 49438 41862 49490 41914
rect 59246 41862 59298 41914
rect 59310 41862 59362 41914
rect 59374 41862 59426 41914
rect 59438 41862 59490 41914
rect 37832 41760 37884 41812
rect 66904 41760 66956 41812
rect 21364 41692 21416 41744
rect 30748 41735 30800 41744
rect 30748 41701 30757 41735
rect 30757 41701 30791 41735
rect 30791 41701 30800 41735
rect 30748 41692 30800 41701
rect 31392 41692 31444 41744
rect 17684 41624 17736 41676
rect 16948 41420 17000 41472
rect 17960 41667 18012 41676
rect 17960 41633 17969 41667
rect 17969 41633 18003 41667
rect 18003 41633 18012 41667
rect 17960 41624 18012 41633
rect 18144 41624 18196 41676
rect 18604 41624 18656 41676
rect 52092 41624 52144 41676
rect 41604 41556 41656 41608
rect 28264 41488 28316 41540
rect 28448 41488 28500 41540
rect 62304 41488 62356 41540
rect 68100 41531 68152 41540
rect 68100 41497 68109 41531
rect 68109 41497 68143 41531
rect 68143 41497 68152 41531
rect 68100 41488 68152 41497
rect 36728 41420 36780 41472
rect 37188 41420 37240 41472
rect 57704 41463 57756 41472
rect 57704 41429 57713 41463
rect 57713 41429 57747 41463
rect 57747 41429 57756 41463
rect 57704 41420 57756 41429
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 14246 41318 14298 41370
rect 14310 41318 14362 41370
rect 14374 41318 14426 41370
rect 14438 41318 14490 41370
rect 24246 41318 24298 41370
rect 24310 41318 24362 41370
rect 24374 41318 24426 41370
rect 24438 41318 24490 41370
rect 34246 41318 34298 41370
rect 34310 41318 34362 41370
rect 34374 41318 34426 41370
rect 34438 41318 34490 41370
rect 44246 41318 44298 41370
rect 44310 41318 44362 41370
rect 44374 41318 44426 41370
rect 44438 41318 44490 41370
rect 54246 41318 54298 41370
rect 54310 41318 54362 41370
rect 54374 41318 54426 41370
rect 54438 41318 54490 41370
rect 64246 41318 64298 41370
rect 64310 41318 64362 41370
rect 64374 41318 64426 41370
rect 64438 41318 64490 41370
rect 13820 41012 13872 41064
rect 47032 41055 47084 41064
rect 47032 41021 47041 41055
rect 47041 41021 47075 41055
rect 47075 41021 47084 41055
rect 47032 41012 47084 41021
rect 65340 41012 65392 41064
rect 17500 40919 17552 40928
rect 17500 40885 17509 40919
rect 17509 40885 17543 40919
rect 17543 40885 17552 40919
rect 17500 40876 17552 40885
rect 18604 40919 18656 40928
rect 18604 40885 18613 40919
rect 18613 40885 18647 40919
rect 18647 40885 18656 40919
rect 18604 40876 18656 40885
rect 39120 40876 39172 40928
rect 9246 40774 9298 40826
rect 9310 40774 9362 40826
rect 9374 40774 9426 40826
rect 9438 40774 9490 40826
rect 19246 40774 19298 40826
rect 19310 40774 19362 40826
rect 19374 40774 19426 40826
rect 19438 40774 19490 40826
rect 29246 40774 29298 40826
rect 29310 40774 29362 40826
rect 29374 40774 29426 40826
rect 29438 40774 29490 40826
rect 39246 40774 39298 40826
rect 39310 40774 39362 40826
rect 39374 40774 39426 40826
rect 39438 40774 39490 40826
rect 49246 40774 49298 40826
rect 49310 40774 49362 40826
rect 49374 40774 49426 40826
rect 49438 40774 49490 40826
rect 59246 40774 59298 40826
rect 59310 40774 59362 40826
rect 59374 40774 59426 40826
rect 59438 40774 59490 40826
rect 1860 40715 1912 40724
rect 1860 40681 1869 40715
rect 1869 40681 1903 40715
rect 1903 40681 1912 40715
rect 1860 40672 1912 40681
rect 17500 40672 17552 40724
rect 17960 40672 18012 40724
rect 50896 40672 50948 40724
rect 65708 40672 65760 40724
rect 2412 40536 2464 40588
rect 22928 40579 22980 40588
rect 22928 40545 22937 40579
rect 22937 40545 22971 40579
rect 22971 40545 22980 40579
rect 22928 40536 22980 40545
rect 39120 40468 39172 40520
rect 39856 40468 39908 40520
rect 2412 40332 2464 40384
rect 23020 40375 23072 40384
rect 23020 40341 23029 40375
rect 23029 40341 23063 40375
rect 23063 40341 23072 40375
rect 23020 40332 23072 40341
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 14246 40230 14298 40282
rect 14310 40230 14362 40282
rect 14374 40230 14426 40282
rect 14438 40230 14490 40282
rect 24246 40230 24298 40282
rect 24310 40230 24362 40282
rect 24374 40230 24426 40282
rect 24438 40230 24490 40282
rect 34246 40230 34298 40282
rect 34310 40230 34362 40282
rect 34374 40230 34426 40282
rect 34438 40230 34490 40282
rect 44246 40230 44298 40282
rect 44310 40230 44362 40282
rect 44374 40230 44426 40282
rect 44438 40230 44490 40282
rect 54246 40230 54298 40282
rect 54310 40230 54362 40282
rect 54374 40230 54426 40282
rect 54438 40230 54490 40282
rect 64246 40230 64298 40282
rect 64310 40230 64362 40282
rect 64374 40230 64426 40282
rect 64438 40230 64490 40282
rect 68100 39967 68152 39976
rect 68100 39933 68109 39967
rect 68109 39933 68143 39967
rect 68143 39933 68152 39967
rect 68100 39924 68152 39933
rect 9246 39686 9298 39738
rect 9310 39686 9362 39738
rect 9374 39686 9426 39738
rect 9438 39686 9490 39738
rect 19246 39686 19298 39738
rect 19310 39686 19362 39738
rect 19374 39686 19426 39738
rect 19438 39686 19490 39738
rect 29246 39686 29298 39738
rect 29310 39686 29362 39738
rect 29374 39686 29426 39738
rect 29438 39686 29490 39738
rect 39246 39686 39298 39738
rect 39310 39686 39362 39738
rect 39374 39686 39426 39738
rect 39438 39686 39490 39738
rect 49246 39686 49298 39738
rect 49310 39686 49362 39738
rect 49374 39686 49426 39738
rect 49438 39686 49490 39738
rect 59246 39686 59298 39738
rect 59310 39686 59362 39738
rect 59374 39686 59426 39738
rect 59438 39686 59490 39738
rect 2596 39627 2648 39636
rect 2596 39593 2605 39627
rect 2605 39593 2639 39627
rect 2639 39593 2648 39627
rect 2596 39584 2648 39593
rect 1768 39491 1820 39500
rect 1768 39457 1777 39491
rect 1777 39457 1811 39491
rect 1811 39457 1820 39491
rect 1768 39448 1820 39457
rect 9772 39380 9824 39432
rect 64788 39380 64840 39432
rect 2688 39312 2740 39364
rect 66996 39312 67048 39364
rect 29000 39244 29052 39296
rect 33416 39244 33468 39296
rect 33692 39244 33744 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 14246 39142 14298 39194
rect 14310 39142 14362 39194
rect 14374 39142 14426 39194
rect 14438 39142 14490 39194
rect 24246 39142 24298 39194
rect 24310 39142 24362 39194
rect 24374 39142 24426 39194
rect 24438 39142 24490 39194
rect 34246 39142 34298 39194
rect 34310 39142 34362 39194
rect 34374 39142 34426 39194
rect 34438 39142 34490 39194
rect 44246 39142 44298 39194
rect 44310 39142 44362 39194
rect 44374 39142 44426 39194
rect 44438 39142 44490 39194
rect 54246 39142 54298 39194
rect 54310 39142 54362 39194
rect 54374 39142 54426 39194
rect 54438 39142 54490 39194
rect 64246 39142 64298 39194
rect 64310 39142 64362 39194
rect 64374 39142 64426 39194
rect 64438 39142 64490 39194
rect 33140 38972 33192 39024
rect 33600 38972 33652 39024
rect 33692 38904 33744 38956
rect 17040 38700 17092 38752
rect 34704 38811 34756 38820
rect 34704 38777 34713 38811
rect 34713 38777 34747 38811
rect 34747 38777 34756 38811
rect 34704 38768 34756 38777
rect 63316 38836 63368 38888
rect 55680 38700 55732 38752
rect 9246 38598 9298 38650
rect 9310 38598 9362 38650
rect 9374 38598 9426 38650
rect 9438 38598 9490 38650
rect 19246 38598 19298 38650
rect 19310 38598 19362 38650
rect 19374 38598 19426 38650
rect 19438 38598 19490 38650
rect 29246 38598 29298 38650
rect 29310 38598 29362 38650
rect 29374 38598 29426 38650
rect 29438 38598 29490 38650
rect 39246 38598 39298 38650
rect 39310 38598 39362 38650
rect 39374 38598 39426 38650
rect 39438 38598 39490 38650
rect 49246 38598 49298 38650
rect 49310 38598 49362 38650
rect 49374 38598 49426 38650
rect 49438 38598 49490 38650
rect 59246 38598 59298 38650
rect 59310 38598 59362 38650
rect 59374 38598 59426 38650
rect 59438 38598 59490 38650
rect 40776 38496 40828 38548
rect 43720 38496 43772 38548
rect 33600 38199 33652 38208
rect 33600 38165 33609 38199
rect 33609 38165 33643 38199
rect 33643 38165 33652 38199
rect 33600 38156 33652 38165
rect 40960 38199 41012 38208
rect 40960 38165 40969 38199
rect 40969 38165 41003 38199
rect 41003 38165 41012 38199
rect 40960 38156 41012 38165
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 14246 38054 14298 38106
rect 14310 38054 14362 38106
rect 14374 38054 14426 38106
rect 14438 38054 14490 38106
rect 24246 38054 24298 38106
rect 24310 38054 24362 38106
rect 24374 38054 24426 38106
rect 24438 38054 24490 38106
rect 34246 38054 34298 38106
rect 34310 38054 34362 38106
rect 34374 38054 34426 38106
rect 34438 38054 34490 38106
rect 44246 38054 44298 38106
rect 44310 38054 44362 38106
rect 44374 38054 44426 38106
rect 44438 38054 44490 38106
rect 54246 38054 54298 38106
rect 54310 38054 54362 38106
rect 54374 38054 54426 38106
rect 54438 38054 54490 38106
rect 64246 38054 64298 38106
rect 64310 38054 64362 38106
rect 64374 38054 64426 38106
rect 64438 38054 64490 38106
rect 5724 37952 5776 38004
rect 40960 37952 41012 38004
rect 12808 37884 12860 37936
rect 29000 37884 29052 37936
rect 4896 37748 4948 37800
rect 40684 37791 40736 37800
rect 40684 37757 40693 37791
rect 40693 37757 40727 37791
rect 40727 37757 40736 37791
rect 40684 37748 40736 37757
rect 62212 37680 62264 37732
rect 66904 37680 66956 37732
rect 68100 37723 68152 37732
rect 68100 37689 68109 37723
rect 68109 37689 68143 37723
rect 68143 37689 68152 37723
rect 68100 37680 68152 37689
rect 9246 37510 9298 37562
rect 9310 37510 9362 37562
rect 9374 37510 9426 37562
rect 9438 37510 9490 37562
rect 19246 37510 19298 37562
rect 19310 37510 19362 37562
rect 19374 37510 19426 37562
rect 19438 37510 19490 37562
rect 29246 37510 29298 37562
rect 29310 37510 29362 37562
rect 29374 37510 29426 37562
rect 29438 37510 29490 37562
rect 39246 37510 39298 37562
rect 39310 37510 39362 37562
rect 39374 37510 39426 37562
rect 39438 37510 39490 37562
rect 49246 37510 49298 37562
rect 49310 37510 49362 37562
rect 49374 37510 49426 37562
rect 49438 37510 49490 37562
rect 59246 37510 59298 37562
rect 59310 37510 59362 37562
rect 59374 37510 59426 37562
rect 59438 37510 59490 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 14246 36966 14298 37018
rect 14310 36966 14362 37018
rect 14374 36966 14426 37018
rect 14438 36966 14490 37018
rect 24246 36966 24298 37018
rect 24310 36966 24362 37018
rect 24374 36966 24426 37018
rect 24438 36966 24490 37018
rect 34246 36966 34298 37018
rect 34310 36966 34362 37018
rect 34374 36966 34426 37018
rect 34438 36966 34490 37018
rect 44246 36966 44298 37018
rect 44310 36966 44362 37018
rect 44374 36966 44426 37018
rect 44438 36966 44490 37018
rect 54246 36966 54298 37018
rect 54310 36966 54362 37018
rect 54374 36966 54426 37018
rect 54438 36966 54490 37018
rect 64246 36966 64298 37018
rect 64310 36966 64362 37018
rect 64374 36966 64426 37018
rect 64438 36966 64490 37018
rect 1584 36703 1636 36712
rect 1584 36669 1593 36703
rect 1593 36669 1627 36703
rect 1627 36669 1636 36703
rect 1584 36660 1636 36669
rect 9246 36422 9298 36474
rect 9310 36422 9362 36474
rect 9374 36422 9426 36474
rect 9438 36422 9490 36474
rect 19246 36422 19298 36474
rect 19310 36422 19362 36474
rect 19374 36422 19426 36474
rect 19438 36422 19490 36474
rect 29246 36422 29298 36474
rect 29310 36422 29362 36474
rect 29374 36422 29426 36474
rect 29438 36422 29490 36474
rect 39246 36422 39298 36474
rect 39310 36422 39362 36474
rect 39374 36422 39426 36474
rect 39438 36422 39490 36474
rect 49246 36422 49298 36474
rect 49310 36422 49362 36474
rect 49374 36422 49426 36474
rect 49438 36422 49490 36474
rect 59246 36422 59298 36474
rect 59310 36422 59362 36474
rect 59374 36422 59426 36474
rect 59438 36422 59490 36474
rect 59544 36184 59596 36236
rect 66996 36184 67048 36236
rect 68100 36227 68152 36236
rect 68100 36193 68109 36227
rect 68109 36193 68143 36227
rect 68143 36193 68152 36227
rect 68100 36184 68152 36193
rect 41604 36116 41656 36168
rect 42064 36159 42116 36168
rect 42064 36125 42073 36159
rect 42073 36125 42107 36159
rect 42107 36125 42116 36159
rect 42064 36116 42116 36125
rect 2872 36023 2924 36032
rect 2872 35989 2881 36023
rect 2881 35989 2915 36023
rect 2915 35989 2924 36023
rect 2872 35980 2924 35989
rect 38200 35980 38252 36032
rect 42064 35980 42116 36032
rect 43168 36023 43220 36032
rect 43168 35989 43177 36023
rect 43177 35989 43211 36023
rect 43211 35989 43220 36023
rect 43168 35980 43220 35989
rect 51264 35980 51316 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 14246 35878 14298 35930
rect 14310 35878 14362 35930
rect 14374 35878 14426 35930
rect 14438 35878 14490 35930
rect 24246 35878 24298 35930
rect 24310 35878 24362 35930
rect 24374 35878 24426 35930
rect 24438 35878 24490 35930
rect 34246 35878 34298 35930
rect 34310 35878 34362 35930
rect 34374 35878 34426 35930
rect 34438 35878 34490 35930
rect 44246 35878 44298 35930
rect 44310 35878 44362 35930
rect 44374 35878 44426 35930
rect 44438 35878 44490 35930
rect 54246 35878 54298 35930
rect 54310 35878 54362 35930
rect 54374 35878 54426 35930
rect 54438 35878 54490 35930
rect 64246 35878 64298 35930
rect 64310 35878 64362 35930
rect 64374 35878 64426 35930
rect 64438 35878 64490 35930
rect 60004 35776 60056 35828
rect 61568 35776 61620 35828
rect 58716 35708 58768 35760
rect 60924 35708 60976 35760
rect 5356 35640 5408 35692
rect 67916 35640 67968 35692
rect 1768 35615 1820 35624
rect 1768 35581 1777 35615
rect 1777 35581 1811 35615
rect 1811 35581 1820 35615
rect 1768 35572 1820 35581
rect 7196 35615 7248 35624
rect 7196 35581 7205 35615
rect 7205 35581 7239 35615
rect 7239 35581 7248 35615
rect 7196 35572 7248 35581
rect 50160 35572 50212 35624
rect 60372 35572 60424 35624
rect 10324 35436 10376 35488
rect 41604 35436 41656 35488
rect 61568 35615 61620 35624
rect 61568 35581 61577 35615
rect 61577 35581 61611 35615
rect 61611 35581 61620 35615
rect 61568 35572 61620 35581
rect 60924 35436 60976 35488
rect 9246 35334 9298 35386
rect 9310 35334 9362 35386
rect 9374 35334 9426 35386
rect 9438 35334 9490 35386
rect 19246 35334 19298 35386
rect 19310 35334 19362 35386
rect 19374 35334 19426 35386
rect 19438 35334 19490 35386
rect 29246 35334 29298 35386
rect 29310 35334 29362 35386
rect 29374 35334 29426 35386
rect 29438 35334 29490 35386
rect 39246 35334 39298 35386
rect 39310 35334 39362 35386
rect 39374 35334 39426 35386
rect 39438 35334 39490 35386
rect 49246 35334 49298 35386
rect 49310 35334 49362 35386
rect 49374 35334 49426 35386
rect 49438 35334 49490 35386
rect 59246 35334 59298 35386
rect 59310 35334 59362 35386
rect 59374 35334 59426 35386
rect 59438 35334 59490 35386
rect 2504 35164 2556 35216
rect 44088 35164 44140 35216
rect 60372 35164 60424 35216
rect 65892 35164 65944 35216
rect 1308 35096 1360 35148
rect 32956 35096 33008 35148
rect 36452 35096 36504 35148
rect 67916 35139 67968 35148
rect 67916 35105 67925 35139
rect 67925 35105 67959 35139
rect 67959 35105 67968 35139
rect 67916 35096 67968 35105
rect 9036 35028 9088 35080
rect 39948 35028 40000 35080
rect 8392 34960 8444 35012
rect 12992 34960 13044 35012
rect 35072 34960 35124 35012
rect 67824 34960 67876 35012
rect 6092 34892 6144 34944
rect 11612 34892 11664 34944
rect 30564 34892 30616 34944
rect 34796 34892 34848 34944
rect 56048 34892 56100 34944
rect 57888 34892 57940 34944
rect 68928 34935 68980 34944
rect 68928 34901 68937 34935
rect 68937 34901 68971 34935
rect 68971 34901 68980 34935
rect 68928 34892 68980 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 14246 34790 14298 34842
rect 14310 34790 14362 34842
rect 14374 34790 14426 34842
rect 14438 34790 14490 34842
rect 24246 34790 24298 34842
rect 24310 34790 24362 34842
rect 24374 34790 24426 34842
rect 24438 34790 24490 34842
rect 34246 34790 34298 34842
rect 34310 34790 34362 34842
rect 34374 34790 34426 34842
rect 34438 34790 34490 34842
rect 44246 34790 44298 34842
rect 44310 34790 44362 34842
rect 44374 34790 44426 34842
rect 44438 34790 44490 34842
rect 54246 34790 54298 34842
rect 54310 34790 54362 34842
rect 54374 34790 54426 34842
rect 54438 34790 54490 34842
rect 64246 34790 64298 34842
rect 64310 34790 64362 34842
rect 64374 34790 64426 34842
rect 64438 34790 64490 34842
rect 7104 34688 7156 34740
rect 8392 34731 8444 34740
rect 8392 34697 8401 34731
rect 8401 34697 8435 34731
rect 8435 34697 8444 34731
rect 8392 34688 8444 34697
rect 9036 34731 9088 34740
rect 9036 34697 9045 34731
rect 9045 34697 9079 34731
rect 9079 34697 9088 34731
rect 9036 34688 9088 34697
rect 57888 34688 57940 34740
rect 66812 34688 66864 34740
rect 32036 34663 32088 34672
rect 32036 34629 32045 34663
rect 32045 34629 32079 34663
rect 32079 34629 32088 34663
rect 32036 34620 32088 34629
rect 33232 34620 33284 34672
rect 35072 34620 35124 34672
rect 36452 34620 36504 34672
rect 67272 34620 67324 34672
rect 9036 34552 9088 34604
rect 11612 34552 11664 34604
rect 32772 34552 32824 34604
rect 33140 34595 33192 34604
rect 33140 34561 33149 34595
rect 33149 34561 33183 34595
rect 33183 34561 33192 34595
rect 33140 34552 33192 34561
rect 33876 34552 33928 34604
rect 9588 34527 9640 34536
rect 9588 34493 9597 34527
rect 9597 34493 9631 34527
rect 9631 34493 9640 34527
rect 9588 34484 9640 34493
rect 32956 34484 33008 34536
rect 33324 34527 33376 34536
rect 33324 34493 33344 34527
rect 33344 34493 33376 34527
rect 33324 34484 33376 34493
rect 31760 34416 31812 34468
rect 32036 34416 32088 34468
rect 33140 34348 33192 34400
rect 35072 34484 35124 34536
rect 44088 34484 44140 34536
rect 34796 34348 34848 34400
rect 9246 34246 9298 34298
rect 9310 34246 9362 34298
rect 9374 34246 9426 34298
rect 9438 34246 9490 34298
rect 19246 34246 19298 34298
rect 19310 34246 19362 34298
rect 19374 34246 19426 34298
rect 19438 34246 19490 34298
rect 29246 34246 29298 34298
rect 29310 34246 29362 34298
rect 29374 34246 29426 34298
rect 29438 34246 29490 34298
rect 39246 34246 39298 34298
rect 39310 34246 39362 34298
rect 39374 34246 39426 34298
rect 39438 34246 39490 34298
rect 49246 34246 49298 34298
rect 49310 34246 49362 34298
rect 49374 34246 49426 34298
rect 49438 34246 49490 34298
rect 59246 34246 59298 34298
rect 59310 34246 59362 34298
rect 59374 34246 59426 34298
rect 59438 34246 59490 34298
rect 1860 34187 1912 34196
rect 1860 34153 1869 34187
rect 1869 34153 1903 34187
rect 1903 34153 1912 34187
rect 1860 34144 1912 34153
rect 32496 34144 32548 34196
rect 33324 34144 33376 34196
rect 33232 34076 33284 34128
rect 33784 34076 33836 34128
rect 2136 34008 2188 34060
rect 10140 34051 10192 34060
rect 10140 34017 10149 34051
rect 10149 34017 10183 34051
rect 10183 34017 10192 34051
rect 10140 34008 10192 34017
rect 2136 33804 2188 33856
rect 55312 33847 55364 33856
rect 55312 33813 55321 33847
rect 55321 33813 55355 33847
rect 55355 33813 55364 33847
rect 55312 33804 55364 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 14246 33702 14298 33754
rect 14310 33702 14362 33754
rect 14374 33702 14426 33754
rect 14438 33702 14490 33754
rect 24246 33702 24298 33754
rect 24310 33702 24362 33754
rect 24374 33702 24426 33754
rect 24438 33702 24490 33754
rect 34246 33702 34298 33754
rect 34310 33702 34362 33754
rect 34374 33702 34426 33754
rect 34438 33702 34490 33754
rect 44246 33702 44298 33754
rect 44310 33702 44362 33754
rect 44374 33702 44426 33754
rect 44438 33702 44490 33754
rect 54246 33702 54298 33754
rect 54310 33702 54362 33754
rect 54374 33702 54426 33754
rect 54438 33702 54490 33754
rect 64246 33702 64298 33754
rect 64310 33702 64362 33754
rect 64374 33702 64426 33754
rect 64438 33702 64490 33754
rect 67180 33464 67232 33516
rect 57336 33396 57388 33448
rect 62948 33439 63000 33448
rect 62948 33405 62957 33439
rect 62957 33405 62991 33439
rect 62991 33405 63000 33439
rect 62948 33396 63000 33405
rect 62856 33328 62908 33380
rect 9246 33158 9298 33210
rect 9310 33158 9362 33210
rect 9374 33158 9426 33210
rect 9438 33158 9490 33210
rect 19246 33158 19298 33210
rect 19310 33158 19362 33210
rect 19374 33158 19426 33210
rect 19438 33158 19490 33210
rect 29246 33158 29298 33210
rect 29310 33158 29362 33210
rect 29374 33158 29426 33210
rect 29438 33158 29490 33210
rect 39246 33158 39298 33210
rect 39310 33158 39362 33210
rect 39374 33158 39426 33210
rect 39438 33158 39490 33210
rect 49246 33158 49298 33210
rect 49310 33158 49362 33210
rect 49374 33158 49426 33210
rect 49438 33158 49490 33210
rect 59246 33158 59298 33210
rect 59310 33158 59362 33210
rect 59374 33158 59426 33210
rect 59438 33158 59490 33210
rect 64880 32759 64932 32768
rect 64880 32725 64889 32759
rect 64889 32725 64923 32759
rect 64923 32725 64932 32759
rect 64880 32716 64932 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 14246 32614 14298 32666
rect 14310 32614 14362 32666
rect 14374 32614 14426 32666
rect 14438 32614 14490 32666
rect 24246 32614 24298 32666
rect 24310 32614 24362 32666
rect 24374 32614 24426 32666
rect 24438 32614 24490 32666
rect 34246 32614 34298 32666
rect 34310 32614 34362 32666
rect 34374 32614 34426 32666
rect 34438 32614 34490 32666
rect 44246 32614 44298 32666
rect 44310 32614 44362 32666
rect 44374 32614 44426 32666
rect 44438 32614 44490 32666
rect 54246 32614 54298 32666
rect 54310 32614 54362 32666
rect 54374 32614 54426 32666
rect 54438 32614 54490 32666
rect 64246 32614 64298 32666
rect 64310 32614 64362 32666
rect 64374 32614 64426 32666
rect 64438 32614 64490 32666
rect 49884 32444 49936 32496
rect 62396 32444 62448 32496
rect 16764 32376 16816 32428
rect 30472 32376 30524 32428
rect 41236 32376 41288 32428
rect 65156 32376 65208 32428
rect 17684 32308 17736 32360
rect 66352 32240 66404 32292
rect 68100 32283 68152 32292
rect 68100 32249 68109 32283
rect 68109 32249 68143 32283
rect 68143 32249 68152 32283
rect 68100 32240 68152 32249
rect 9246 32070 9298 32122
rect 9310 32070 9362 32122
rect 9374 32070 9426 32122
rect 9438 32070 9490 32122
rect 19246 32070 19298 32122
rect 19310 32070 19362 32122
rect 19374 32070 19426 32122
rect 19438 32070 19490 32122
rect 29246 32070 29298 32122
rect 29310 32070 29362 32122
rect 29374 32070 29426 32122
rect 29438 32070 29490 32122
rect 39246 32070 39298 32122
rect 39310 32070 39362 32122
rect 39374 32070 39426 32122
rect 39438 32070 39490 32122
rect 49246 32070 49298 32122
rect 49310 32070 49362 32122
rect 49374 32070 49426 32122
rect 49438 32070 49490 32122
rect 59246 32070 59298 32122
rect 59310 32070 59362 32122
rect 59374 32070 59426 32122
rect 59438 32070 59490 32122
rect 1584 31875 1636 31884
rect 1584 31841 1593 31875
rect 1593 31841 1627 31875
rect 1627 31841 1636 31875
rect 1584 31832 1636 31841
rect 26884 31875 26936 31884
rect 26884 31841 26893 31875
rect 26893 31841 26927 31875
rect 26927 31841 26936 31875
rect 26884 31832 26936 31841
rect 39580 31968 39632 32020
rect 42432 31968 42484 32020
rect 61844 31968 61896 32020
rect 33784 31900 33836 31952
rect 36636 31943 36688 31952
rect 36636 31909 36645 31943
rect 36645 31909 36679 31943
rect 36679 31909 36688 31943
rect 36636 31900 36688 31909
rect 37004 31832 37056 31884
rect 39948 31900 40000 31952
rect 43812 31832 43864 31884
rect 47492 31832 47544 31884
rect 55680 31900 55732 31952
rect 56232 31832 56284 31884
rect 58716 31900 58768 31952
rect 49884 31764 49936 31816
rect 37648 31739 37700 31748
rect 37648 31705 37657 31739
rect 37657 31705 37691 31739
rect 37691 31705 37700 31739
rect 37648 31696 37700 31705
rect 42432 31739 42484 31748
rect 42432 31705 42441 31739
rect 42441 31705 42475 31739
rect 42475 31705 42484 31739
rect 42432 31696 42484 31705
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 14246 31526 14298 31578
rect 14310 31526 14362 31578
rect 14374 31526 14426 31578
rect 14438 31526 14490 31578
rect 24246 31526 24298 31578
rect 24310 31526 24362 31578
rect 24374 31526 24426 31578
rect 24438 31526 24490 31578
rect 34246 31526 34298 31578
rect 34310 31526 34362 31578
rect 34374 31526 34426 31578
rect 34438 31526 34490 31578
rect 44246 31526 44298 31578
rect 44310 31526 44362 31578
rect 44374 31526 44426 31578
rect 44438 31526 44490 31578
rect 54246 31526 54298 31578
rect 54310 31526 54362 31578
rect 54374 31526 54426 31578
rect 54438 31526 54490 31578
rect 64246 31526 64298 31578
rect 64310 31526 64362 31578
rect 64374 31526 64426 31578
rect 64438 31526 64490 31578
rect 31760 31424 31812 31476
rect 37648 31424 37700 31476
rect 9246 30982 9298 31034
rect 9310 30982 9362 31034
rect 9374 30982 9426 31034
rect 9438 30982 9490 31034
rect 19246 30982 19298 31034
rect 19310 30982 19362 31034
rect 19374 30982 19426 31034
rect 19438 30982 19490 31034
rect 29246 30982 29298 31034
rect 29310 30982 29362 31034
rect 29374 30982 29426 31034
rect 29438 30982 29490 31034
rect 39246 30982 39298 31034
rect 39310 30982 39362 31034
rect 39374 30982 39426 31034
rect 39438 30982 39490 31034
rect 49246 30982 49298 31034
rect 49310 30982 49362 31034
rect 49374 30982 49426 31034
rect 49438 30982 49490 31034
rect 59246 30982 59298 31034
rect 59310 30982 59362 31034
rect 59374 30982 59426 31034
rect 59438 30982 59490 31034
rect 30564 30880 30616 30932
rect 37096 30812 37148 30864
rect 40316 30812 40368 30864
rect 67548 30812 67600 30864
rect 68100 30855 68152 30864
rect 68100 30821 68109 30855
rect 68109 30821 68143 30855
rect 68143 30821 68152 30855
rect 68100 30812 68152 30821
rect 37648 30787 37700 30796
rect 37648 30753 37697 30787
rect 37697 30753 37700 30787
rect 37648 30744 37700 30753
rect 36452 30676 36504 30728
rect 38660 30744 38712 30796
rect 39120 30787 39172 30796
rect 39120 30753 39129 30787
rect 39129 30753 39163 30787
rect 39163 30753 39172 30787
rect 39120 30744 39172 30753
rect 10876 30608 10928 30660
rect 25228 30583 25280 30592
rect 25228 30549 25237 30583
rect 25237 30549 25271 30583
rect 25271 30549 25280 30583
rect 25228 30540 25280 30549
rect 33692 30540 33744 30592
rect 37556 30583 37608 30592
rect 37556 30549 37565 30583
rect 37565 30549 37599 30583
rect 37599 30549 37608 30583
rect 37556 30540 37608 30549
rect 37648 30540 37700 30592
rect 48964 30540 49016 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 14246 30438 14298 30490
rect 14310 30438 14362 30490
rect 14374 30438 14426 30490
rect 14438 30438 14490 30490
rect 24246 30438 24298 30490
rect 24310 30438 24362 30490
rect 24374 30438 24426 30490
rect 24438 30438 24490 30490
rect 34246 30438 34298 30490
rect 34310 30438 34362 30490
rect 34374 30438 34426 30490
rect 34438 30438 34490 30490
rect 44246 30438 44298 30490
rect 44310 30438 44362 30490
rect 44374 30438 44426 30490
rect 44438 30438 44490 30490
rect 54246 30438 54298 30490
rect 54310 30438 54362 30490
rect 54374 30438 54426 30490
rect 54438 30438 54490 30490
rect 64246 30438 64298 30490
rect 64310 30438 64362 30490
rect 64374 30438 64426 30490
rect 64438 30438 64490 30490
rect 12992 30336 13044 30388
rect 15200 30336 15252 30388
rect 1768 30311 1820 30320
rect 1768 30277 1777 30311
rect 1777 30277 1811 30311
rect 1811 30277 1820 30311
rect 1768 30268 1820 30277
rect 2688 30311 2740 30320
rect 2688 30277 2697 30311
rect 2697 30277 2731 30311
rect 2731 30277 2740 30311
rect 2688 30268 2740 30277
rect 36452 30336 36504 30388
rect 42432 30336 42484 30388
rect 37096 30311 37148 30320
rect 37096 30277 37105 30311
rect 37105 30277 37139 30311
rect 37139 30277 37148 30311
rect 37096 30268 37148 30277
rect 48964 30200 49016 30252
rect 12072 30175 12124 30184
rect 12072 30141 12081 30175
rect 12081 30141 12115 30175
rect 12115 30141 12124 30175
rect 12072 30132 12124 30141
rect 27620 30132 27672 30184
rect 38936 30175 38988 30184
rect 38936 30141 38945 30175
rect 38945 30141 38979 30175
rect 38979 30141 38988 30175
rect 38936 30132 38988 30141
rect 2228 30064 2280 30116
rect 17868 30064 17920 30116
rect 32864 30064 32916 30116
rect 32404 29996 32456 30048
rect 9246 29894 9298 29946
rect 9310 29894 9362 29946
rect 9374 29894 9426 29946
rect 9438 29894 9490 29946
rect 19246 29894 19298 29946
rect 19310 29894 19362 29946
rect 19374 29894 19426 29946
rect 19438 29894 19490 29946
rect 29246 29894 29298 29946
rect 29310 29894 29362 29946
rect 29374 29894 29426 29946
rect 29438 29894 29490 29946
rect 39246 29894 39298 29946
rect 39310 29894 39362 29946
rect 39374 29894 39426 29946
rect 39438 29894 39490 29946
rect 49246 29894 49298 29946
rect 49310 29894 49362 29946
rect 49374 29894 49426 29946
rect 49438 29894 49490 29946
rect 59246 29894 59298 29946
rect 59310 29894 59362 29946
rect 59374 29894 59426 29946
rect 59438 29894 59490 29946
rect 28540 29792 28592 29844
rect 29552 29724 29604 29776
rect 50712 29724 50764 29776
rect 2964 29656 3016 29708
rect 26884 29699 26936 29708
rect 26884 29665 26893 29699
rect 26893 29665 26927 29699
rect 26927 29665 26936 29699
rect 26884 29656 26936 29665
rect 54760 29656 54812 29708
rect 68100 29699 68152 29708
rect 68100 29665 68109 29699
rect 68109 29665 68143 29699
rect 68143 29665 68152 29699
rect 68100 29656 68152 29665
rect 28540 29588 28592 29640
rect 50252 29588 50304 29640
rect 53012 29520 53064 29572
rect 2228 29495 2280 29504
rect 2228 29461 2237 29495
rect 2237 29461 2271 29495
rect 2271 29461 2280 29495
rect 2228 29452 2280 29461
rect 7380 29452 7432 29504
rect 20996 29495 21048 29504
rect 20996 29461 21005 29495
rect 21005 29461 21039 29495
rect 21039 29461 21048 29495
rect 20996 29452 21048 29461
rect 26332 29495 26384 29504
rect 26332 29461 26341 29495
rect 26341 29461 26375 29495
rect 26375 29461 26384 29495
rect 26332 29452 26384 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 14246 29350 14298 29402
rect 14310 29350 14362 29402
rect 14374 29350 14426 29402
rect 14438 29350 14490 29402
rect 24246 29350 24298 29402
rect 24310 29350 24362 29402
rect 24374 29350 24426 29402
rect 24438 29350 24490 29402
rect 34246 29350 34298 29402
rect 34310 29350 34362 29402
rect 34374 29350 34426 29402
rect 34438 29350 34490 29402
rect 44246 29350 44298 29402
rect 44310 29350 44362 29402
rect 44374 29350 44426 29402
rect 44438 29350 44490 29402
rect 54246 29350 54298 29402
rect 54310 29350 54362 29402
rect 54374 29350 54426 29402
rect 54438 29350 54490 29402
rect 64246 29350 64298 29402
rect 64310 29350 64362 29402
rect 64374 29350 64426 29402
rect 64438 29350 64490 29402
rect 2228 29248 2280 29300
rect 16672 29248 16724 29300
rect 17868 29248 17920 29300
rect 20996 29248 21048 29300
rect 64052 29248 64104 29300
rect 26884 29180 26936 29232
rect 34888 29180 34940 29232
rect 1768 29087 1820 29096
rect 1768 29053 1777 29087
rect 1777 29053 1811 29087
rect 1811 29053 1820 29087
rect 1768 29044 1820 29053
rect 2044 29044 2096 29096
rect 4804 29044 4856 29096
rect 4988 28976 5040 29028
rect 9246 28806 9298 28858
rect 9310 28806 9362 28858
rect 9374 28806 9426 28858
rect 9438 28806 9490 28858
rect 19246 28806 19298 28858
rect 19310 28806 19362 28858
rect 19374 28806 19426 28858
rect 19438 28806 19490 28858
rect 29246 28806 29298 28858
rect 29310 28806 29362 28858
rect 29374 28806 29426 28858
rect 29438 28806 29490 28858
rect 39246 28806 39298 28858
rect 39310 28806 39362 28858
rect 39374 28806 39426 28858
rect 39438 28806 39490 28858
rect 49246 28806 49298 28858
rect 49310 28806 49362 28858
rect 49374 28806 49426 28858
rect 49438 28806 49490 28858
rect 59246 28806 59298 28858
rect 59310 28806 59362 28858
rect 59374 28806 59426 28858
rect 59438 28806 59490 28858
rect 23020 28704 23072 28756
rect 31484 28704 31536 28756
rect 66352 28500 66404 28552
rect 31760 28364 31812 28416
rect 38200 28364 38252 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 14246 28262 14298 28314
rect 14310 28262 14362 28314
rect 14374 28262 14426 28314
rect 14438 28262 14490 28314
rect 24246 28262 24298 28314
rect 24310 28262 24362 28314
rect 24374 28262 24426 28314
rect 24438 28262 24490 28314
rect 34246 28262 34298 28314
rect 34310 28262 34362 28314
rect 34374 28262 34426 28314
rect 34438 28262 34490 28314
rect 44246 28262 44298 28314
rect 44310 28262 44362 28314
rect 44374 28262 44426 28314
rect 44438 28262 44490 28314
rect 54246 28262 54298 28314
rect 54310 28262 54362 28314
rect 54374 28262 54426 28314
rect 54438 28262 54490 28314
rect 64246 28262 64298 28314
rect 64310 28262 64362 28314
rect 64374 28262 64426 28314
rect 64438 28262 64490 28314
rect 13544 28160 13596 28212
rect 31760 28160 31812 28212
rect 31668 28092 31720 28144
rect 2320 28024 2372 28076
rect 30932 28024 30984 28076
rect 31392 28024 31444 28076
rect 33140 28160 33192 28212
rect 32036 28092 32088 28144
rect 46112 28092 46164 28144
rect 31484 27956 31536 28008
rect 8484 27888 8536 27940
rect 31576 27888 31628 27940
rect 32036 27956 32088 28008
rect 60464 27999 60516 28008
rect 60464 27965 60473 27999
rect 60473 27965 60507 27999
rect 60507 27965 60516 27999
rect 60464 27956 60516 27965
rect 32220 27820 32272 27872
rect 33232 27863 33284 27872
rect 33232 27829 33241 27863
rect 33241 27829 33275 27863
rect 33275 27829 33284 27863
rect 33232 27820 33284 27829
rect 9246 27718 9298 27770
rect 9310 27718 9362 27770
rect 9374 27718 9426 27770
rect 9438 27718 9490 27770
rect 19246 27718 19298 27770
rect 19310 27718 19362 27770
rect 19374 27718 19426 27770
rect 19438 27718 19490 27770
rect 29246 27718 29298 27770
rect 29310 27718 29362 27770
rect 29374 27718 29426 27770
rect 29438 27718 29490 27770
rect 39246 27718 39298 27770
rect 39310 27718 39362 27770
rect 39374 27718 39426 27770
rect 39438 27718 39490 27770
rect 49246 27718 49298 27770
rect 49310 27718 49362 27770
rect 49374 27718 49426 27770
rect 49438 27718 49490 27770
rect 59246 27718 59298 27770
rect 59310 27718 59362 27770
rect 59374 27718 59426 27770
rect 59438 27718 59490 27770
rect 30196 27616 30248 27668
rect 33140 27616 33192 27668
rect 43628 27616 43680 27668
rect 66168 27616 66220 27668
rect 47584 27548 47636 27600
rect 48228 27548 48280 27600
rect 18236 27480 18288 27532
rect 18788 27412 18840 27464
rect 16672 27387 16724 27396
rect 16672 27353 16681 27387
rect 16681 27353 16715 27387
rect 16715 27353 16724 27387
rect 16672 27344 16724 27353
rect 7196 27276 7248 27328
rect 18512 27319 18564 27328
rect 18512 27285 18521 27319
rect 18521 27285 18555 27319
rect 18555 27285 18564 27319
rect 18512 27276 18564 27285
rect 31116 27319 31168 27328
rect 31116 27285 31125 27319
rect 31125 27285 31159 27319
rect 31159 27285 31168 27319
rect 31116 27276 31168 27285
rect 31576 27276 31628 27328
rect 60924 27276 60976 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 14246 27174 14298 27226
rect 14310 27174 14362 27226
rect 14374 27174 14426 27226
rect 14438 27174 14490 27226
rect 24246 27174 24298 27226
rect 24310 27174 24362 27226
rect 24374 27174 24426 27226
rect 24438 27174 24490 27226
rect 34246 27174 34298 27226
rect 34310 27174 34362 27226
rect 34374 27174 34426 27226
rect 34438 27174 34490 27226
rect 44246 27174 44298 27226
rect 44310 27174 44362 27226
rect 44374 27174 44426 27226
rect 44438 27174 44490 27226
rect 54246 27174 54298 27226
rect 54310 27174 54362 27226
rect 54374 27174 54426 27226
rect 54438 27174 54490 27226
rect 64246 27174 64298 27226
rect 64310 27174 64362 27226
rect 64374 27174 64426 27226
rect 64438 27174 64490 27226
rect 11060 27072 11112 27124
rect 18788 27115 18840 27124
rect 18788 27081 18797 27115
rect 18797 27081 18831 27115
rect 18831 27081 18840 27115
rect 18788 27072 18840 27081
rect 25228 27072 25280 27124
rect 26148 27072 26200 27124
rect 67272 27115 67324 27124
rect 67272 27081 67281 27115
rect 67281 27081 67315 27115
rect 67315 27081 67324 27115
rect 67272 27072 67324 27081
rect 27344 27004 27396 27056
rect 54576 27004 54628 27056
rect 32588 26936 32640 26988
rect 32956 26936 33008 26988
rect 53840 26936 53892 26988
rect 68100 26979 68152 26988
rect 68100 26945 68109 26979
rect 68109 26945 68143 26979
rect 68143 26945 68152 26979
rect 68100 26936 68152 26945
rect 1584 26911 1636 26920
rect 1584 26877 1593 26911
rect 1593 26877 1627 26911
rect 1627 26877 1636 26911
rect 1584 26868 1636 26877
rect 67180 26868 67232 26920
rect 67272 26868 67324 26920
rect 14004 26800 14056 26852
rect 27896 26800 27948 26852
rect 47216 26800 47268 26852
rect 57428 26800 57480 26852
rect 18236 26775 18288 26784
rect 18236 26741 18245 26775
rect 18245 26741 18279 26775
rect 18279 26741 18288 26775
rect 18236 26732 18288 26741
rect 38384 26732 38436 26784
rect 9246 26630 9298 26682
rect 9310 26630 9362 26682
rect 9374 26630 9426 26682
rect 9438 26630 9490 26682
rect 19246 26630 19298 26682
rect 19310 26630 19362 26682
rect 19374 26630 19426 26682
rect 19438 26630 19490 26682
rect 29246 26630 29298 26682
rect 29310 26630 29362 26682
rect 29374 26630 29426 26682
rect 29438 26630 29490 26682
rect 39246 26630 39298 26682
rect 39310 26630 39362 26682
rect 39374 26630 39426 26682
rect 39438 26630 39490 26682
rect 49246 26630 49298 26682
rect 49310 26630 49362 26682
rect 49374 26630 49426 26682
rect 49438 26630 49490 26682
rect 59246 26630 59298 26682
rect 59310 26630 59362 26682
rect 59374 26630 59426 26682
rect 59438 26630 59490 26682
rect 28172 26528 28224 26580
rect 30196 26528 30248 26580
rect 33600 26528 33652 26580
rect 42616 26528 42668 26580
rect 47492 26528 47544 26580
rect 27896 26503 27948 26512
rect 27896 26469 27905 26503
rect 27905 26469 27939 26503
rect 27939 26469 27948 26503
rect 27896 26460 27948 26469
rect 28172 26435 28224 26444
rect 28172 26401 28181 26435
rect 28181 26401 28215 26435
rect 28215 26401 28224 26435
rect 28172 26392 28224 26401
rect 28448 26435 28500 26444
rect 28448 26401 28457 26435
rect 28457 26401 28491 26435
rect 28491 26401 28500 26435
rect 28448 26392 28500 26401
rect 32956 26460 33008 26512
rect 30196 26435 30248 26444
rect 30196 26401 30205 26435
rect 30205 26401 30239 26435
rect 30239 26401 30248 26435
rect 30196 26392 30248 26401
rect 31392 26392 31444 26444
rect 31668 26392 31720 26444
rect 37924 26392 37976 26444
rect 39948 26392 40000 26444
rect 42616 26435 42668 26444
rect 42616 26401 42625 26435
rect 42625 26401 42659 26435
rect 42659 26401 42668 26435
rect 42616 26392 42668 26401
rect 48412 26392 48464 26444
rect 49332 26392 49384 26444
rect 49608 26435 49660 26444
rect 49608 26401 49617 26435
rect 49617 26401 49651 26435
rect 49651 26401 49660 26435
rect 49608 26392 49660 26401
rect 49884 26528 49936 26580
rect 48504 26367 48556 26376
rect 27344 26299 27396 26308
rect 27344 26265 27353 26299
rect 27353 26265 27387 26299
rect 27387 26265 27396 26299
rect 27344 26256 27396 26265
rect 47216 26256 47268 26308
rect 48504 26333 48513 26367
rect 48513 26333 48547 26367
rect 48547 26333 48556 26367
rect 48504 26324 48556 26333
rect 49424 26256 49476 26308
rect 49884 26256 49936 26308
rect 57244 26256 57296 26308
rect 62672 26299 62724 26308
rect 62672 26265 62681 26299
rect 62681 26265 62715 26299
rect 62715 26265 62724 26299
rect 62672 26256 62724 26265
rect 9588 26188 9640 26240
rect 11060 26188 11112 26240
rect 47584 26188 47636 26240
rect 49608 26188 49660 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 14246 26086 14298 26138
rect 14310 26086 14362 26138
rect 14374 26086 14426 26138
rect 14438 26086 14490 26138
rect 24246 26086 24298 26138
rect 24310 26086 24362 26138
rect 24374 26086 24426 26138
rect 24438 26086 24490 26138
rect 34246 26086 34298 26138
rect 34310 26086 34362 26138
rect 34374 26086 34426 26138
rect 34438 26086 34490 26138
rect 44246 26086 44298 26138
rect 44310 26086 44362 26138
rect 44374 26086 44426 26138
rect 44438 26086 44490 26138
rect 54246 26086 54298 26138
rect 54310 26086 54362 26138
rect 54374 26086 54426 26138
rect 54438 26086 54490 26138
rect 64246 26086 64298 26138
rect 64310 26086 64362 26138
rect 64374 26086 64426 26138
rect 64438 26086 64490 26138
rect 28448 25984 28500 26036
rect 67456 25984 67508 26036
rect 2412 25916 2464 25968
rect 15292 25848 15344 25900
rect 36728 25848 36780 25900
rect 13176 25780 13228 25832
rect 58440 25780 58492 25832
rect 67456 25780 67508 25832
rect 17868 25712 17920 25764
rect 42524 25712 42576 25764
rect 56416 25712 56468 25764
rect 68100 25755 68152 25764
rect 68100 25721 68109 25755
rect 68109 25721 68143 25755
rect 68143 25721 68152 25755
rect 68100 25712 68152 25721
rect 47584 25644 47636 25696
rect 48412 25687 48464 25696
rect 48412 25653 48421 25687
rect 48421 25653 48455 25687
rect 48455 25653 48464 25687
rect 48412 25644 48464 25653
rect 9246 25542 9298 25594
rect 9310 25542 9362 25594
rect 9374 25542 9426 25594
rect 9438 25542 9490 25594
rect 19246 25542 19298 25594
rect 19310 25542 19362 25594
rect 19374 25542 19426 25594
rect 19438 25542 19490 25594
rect 29246 25542 29298 25594
rect 29310 25542 29362 25594
rect 29374 25542 29426 25594
rect 29438 25542 29490 25594
rect 39246 25542 39298 25594
rect 39310 25542 39362 25594
rect 39374 25542 39426 25594
rect 39438 25542 39490 25594
rect 49246 25542 49298 25594
rect 49310 25542 49362 25594
rect 49374 25542 49426 25594
rect 49438 25542 49490 25594
rect 59246 25542 59298 25594
rect 59310 25542 59362 25594
rect 59374 25542 59426 25594
rect 59438 25542 59490 25594
rect 1768 25211 1820 25220
rect 1768 25177 1777 25211
rect 1777 25177 1811 25211
rect 1811 25177 1820 25211
rect 1768 25168 1820 25177
rect 13176 25440 13228 25492
rect 66904 25440 66956 25492
rect 15292 25236 15344 25288
rect 2596 25143 2648 25152
rect 2596 25109 2605 25143
rect 2605 25109 2639 25143
rect 2639 25109 2648 25143
rect 2596 25100 2648 25109
rect 7932 25143 7984 25152
rect 7932 25109 7941 25143
rect 7941 25109 7975 25143
rect 7975 25109 7984 25143
rect 7932 25100 7984 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 14246 24998 14298 25050
rect 14310 24998 14362 25050
rect 14374 24998 14426 25050
rect 14438 24998 14490 25050
rect 24246 24998 24298 25050
rect 24310 24998 24362 25050
rect 24374 24998 24426 25050
rect 24438 24998 24490 25050
rect 34246 24998 34298 25050
rect 34310 24998 34362 25050
rect 34374 24998 34426 25050
rect 34438 24998 34490 25050
rect 44246 24998 44298 25050
rect 44310 24998 44362 25050
rect 44374 24998 44426 25050
rect 44438 24998 44490 25050
rect 54246 24998 54298 25050
rect 54310 24998 54362 25050
rect 54374 24998 54426 25050
rect 54438 24998 54490 25050
rect 64246 24998 64298 25050
rect 64310 24998 64362 25050
rect 64374 24998 64426 25050
rect 64438 24998 64490 25050
rect 2596 24896 2648 24948
rect 16580 24896 16632 24948
rect 17868 24896 17920 24948
rect 7932 24828 7984 24880
rect 46480 24828 46532 24880
rect 23480 24760 23532 24812
rect 58532 24760 58584 24812
rect 36912 24735 36964 24744
rect 36912 24701 36921 24735
rect 36921 24701 36955 24735
rect 36955 24701 36964 24735
rect 36912 24692 36964 24701
rect 63500 24692 63552 24744
rect 68100 24735 68152 24744
rect 68100 24701 68109 24735
rect 68109 24701 68143 24735
rect 68143 24701 68152 24735
rect 68100 24692 68152 24701
rect 9246 24454 9298 24506
rect 9310 24454 9362 24506
rect 9374 24454 9426 24506
rect 9438 24454 9490 24506
rect 19246 24454 19298 24506
rect 19310 24454 19362 24506
rect 19374 24454 19426 24506
rect 19438 24454 19490 24506
rect 29246 24454 29298 24506
rect 29310 24454 29362 24506
rect 29374 24454 29426 24506
rect 29438 24454 29490 24506
rect 39246 24454 39298 24506
rect 39310 24454 39362 24506
rect 39374 24454 39426 24506
rect 39438 24454 39490 24506
rect 49246 24454 49298 24506
rect 49310 24454 49362 24506
rect 49374 24454 49426 24506
rect 49438 24454 49490 24506
rect 59246 24454 59298 24506
rect 59310 24454 59362 24506
rect 59374 24454 59426 24506
rect 59438 24454 59490 24506
rect 23480 24395 23532 24404
rect 19984 24216 20036 24268
rect 20628 24216 20680 24268
rect 23480 24361 23489 24395
rect 23489 24361 23523 24395
rect 23523 24361 23532 24395
rect 23480 24352 23532 24361
rect 36544 24216 36596 24268
rect 1860 24148 1912 24200
rect 7472 24080 7524 24132
rect 54760 24080 54812 24132
rect 12348 24055 12400 24064
rect 12348 24021 12357 24055
rect 12357 24021 12391 24055
rect 12391 24021 12400 24055
rect 12348 24012 12400 24021
rect 29092 24055 29144 24064
rect 29092 24021 29101 24055
rect 29101 24021 29135 24055
rect 29135 24021 29144 24055
rect 29092 24012 29144 24021
rect 54116 24055 54168 24064
rect 54116 24021 54125 24055
rect 54125 24021 54159 24055
rect 54159 24021 54168 24055
rect 54116 24012 54168 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 14246 23910 14298 23962
rect 14310 23910 14362 23962
rect 14374 23910 14426 23962
rect 14438 23910 14490 23962
rect 24246 23910 24298 23962
rect 24310 23910 24362 23962
rect 24374 23910 24426 23962
rect 24438 23910 24490 23962
rect 34246 23910 34298 23962
rect 34310 23910 34362 23962
rect 34374 23910 34426 23962
rect 34438 23910 34490 23962
rect 44246 23910 44298 23962
rect 44310 23910 44362 23962
rect 44374 23910 44426 23962
rect 44438 23910 44490 23962
rect 54246 23910 54298 23962
rect 54310 23910 54362 23962
rect 54374 23910 54426 23962
rect 54438 23910 54490 23962
rect 64246 23910 64298 23962
rect 64310 23910 64362 23962
rect 64374 23910 64426 23962
rect 64438 23910 64490 23962
rect 1860 23851 1912 23860
rect 1860 23817 1869 23851
rect 1869 23817 1903 23851
rect 1903 23817 1912 23851
rect 1860 23808 1912 23817
rect 3148 23808 3200 23860
rect 5448 23808 5500 23860
rect 54116 23808 54168 23860
rect 29092 23740 29144 23792
rect 66720 23740 66772 23792
rect 12348 23672 12400 23724
rect 37740 23672 37792 23724
rect 2320 23536 2372 23588
rect 47584 23604 47636 23656
rect 54392 23647 54444 23656
rect 54392 23613 54401 23647
rect 54401 23613 54435 23647
rect 54435 23613 54444 23647
rect 54392 23604 54444 23613
rect 36636 23536 36688 23588
rect 53840 23579 53892 23588
rect 53840 23545 53849 23579
rect 53849 23545 53883 23579
rect 53883 23545 53892 23579
rect 53840 23536 53892 23545
rect 53932 23468 53984 23520
rect 54392 23468 54444 23520
rect 54760 23511 54812 23520
rect 54760 23477 54769 23511
rect 54769 23477 54803 23511
rect 54803 23477 54812 23511
rect 54760 23468 54812 23477
rect 56508 23468 56560 23520
rect 9246 23366 9298 23418
rect 9310 23366 9362 23418
rect 9374 23366 9426 23418
rect 9438 23366 9490 23418
rect 19246 23366 19298 23418
rect 19310 23366 19362 23418
rect 19374 23366 19426 23418
rect 19438 23366 19490 23418
rect 29246 23366 29298 23418
rect 29310 23366 29362 23418
rect 29374 23366 29426 23418
rect 29438 23366 29490 23418
rect 39246 23366 39298 23418
rect 39310 23366 39362 23418
rect 39374 23366 39426 23418
rect 39438 23366 39490 23418
rect 49246 23366 49298 23418
rect 49310 23366 49362 23418
rect 49374 23366 49426 23418
rect 49438 23366 49490 23418
rect 59246 23366 59298 23418
rect 59310 23366 59362 23418
rect 59374 23366 59426 23418
rect 59438 23366 59490 23418
rect 13176 23264 13228 23316
rect 58440 23307 58492 23316
rect 9220 23196 9272 23248
rect 37556 23196 37608 23248
rect 53932 23239 53984 23248
rect 53932 23205 53941 23239
rect 53941 23205 53975 23239
rect 53975 23205 53984 23239
rect 53932 23196 53984 23205
rect 22928 23128 22980 23180
rect 39672 23128 39724 23180
rect 50068 23128 50120 23180
rect 58440 23273 58449 23307
rect 58449 23273 58483 23307
rect 58483 23273 58492 23307
rect 58440 23264 58492 23273
rect 67364 23307 67416 23316
rect 67364 23273 67373 23307
rect 67373 23273 67407 23307
rect 67407 23273 67416 23307
rect 67364 23264 67416 23273
rect 62396 23196 62448 23248
rect 30104 23060 30156 23112
rect 33692 23060 33744 23112
rect 56508 23060 56560 23112
rect 56968 23103 57020 23112
rect 56968 23069 56977 23103
rect 56977 23069 57011 23103
rect 57011 23069 57020 23103
rect 56968 23060 57020 23069
rect 54116 22992 54168 23044
rect 68100 23035 68152 23044
rect 68100 23001 68109 23035
rect 68109 23001 68143 23035
rect 68143 23001 68152 23035
rect 68100 22992 68152 23001
rect 29920 22924 29972 22976
rect 33600 22924 33652 22976
rect 37924 22967 37976 22976
rect 37924 22933 37933 22967
rect 37933 22933 37967 22967
rect 37967 22933 37976 22967
rect 37924 22924 37976 22933
rect 38200 22924 38252 22976
rect 38660 22924 38712 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 14246 22822 14298 22874
rect 14310 22822 14362 22874
rect 14374 22822 14426 22874
rect 14438 22822 14490 22874
rect 24246 22822 24298 22874
rect 24310 22822 24362 22874
rect 24374 22822 24426 22874
rect 24438 22822 24490 22874
rect 34246 22822 34298 22874
rect 34310 22822 34362 22874
rect 34374 22822 34426 22874
rect 34438 22822 34490 22874
rect 44246 22822 44298 22874
rect 44310 22822 44362 22874
rect 44374 22822 44426 22874
rect 44438 22822 44490 22874
rect 54246 22822 54298 22874
rect 54310 22822 54362 22874
rect 54374 22822 54426 22874
rect 54438 22822 54490 22874
rect 64246 22822 64298 22874
rect 64310 22822 64362 22874
rect 64374 22822 64426 22874
rect 64438 22822 64490 22874
rect 3700 22720 3752 22772
rect 9220 22695 9272 22704
rect 9220 22661 9229 22695
rect 9229 22661 9263 22695
rect 9263 22661 9272 22695
rect 9220 22652 9272 22661
rect 13176 22695 13228 22704
rect 13176 22661 13185 22695
rect 13185 22661 13219 22695
rect 13219 22661 13228 22695
rect 13176 22652 13228 22661
rect 29920 22695 29972 22704
rect 29920 22661 29929 22695
rect 29929 22661 29963 22695
rect 29963 22661 29972 22695
rect 29920 22652 29972 22661
rect 26148 22584 26200 22636
rect 31576 22720 31628 22772
rect 34980 22720 35032 22772
rect 38568 22720 38620 22772
rect 39672 22763 39724 22772
rect 39672 22729 39681 22763
rect 39681 22729 39715 22763
rect 39715 22729 39724 22763
rect 39672 22720 39724 22729
rect 64604 22720 64656 22772
rect 8576 22423 8628 22432
rect 8576 22389 8585 22423
rect 8585 22389 8619 22423
rect 8619 22389 8628 22423
rect 8576 22380 8628 22389
rect 30104 22448 30156 22500
rect 38200 22516 38252 22568
rect 56508 22584 56560 22636
rect 11060 22380 11112 22432
rect 11888 22380 11940 22432
rect 29920 22380 29972 22432
rect 31576 22448 31628 22500
rect 37924 22448 37976 22500
rect 37648 22380 37700 22432
rect 37832 22380 37884 22432
rect 46388 22559 46440 22568
rect 46388 22525 46397 22559
rect 46397 22525 46431 22559
rect 46431 22525 46440 22559
rect 46388 22516 46440 22525
rect 38568 22380 38620 22432
rect 56968 22380 57020 22432
rect 9246 22278 9298 22330
rect 9310 22278 9362 22330
rect 9374 22278 9426 22330
rect 9438 22278 9490 22330
rect 19246 22278 19298 22330
rect 19310 22278 19362 22330
rect 19374 22278 19426 22330
rect 19438 22278 19490 22330
rect 29246 22278 29298 22330
rect 29310 22278 29362 22330
rect 29374 22278 29426 22330
rect 29438 22278 29490 22330
rect 39246 22278 39298 22330
rect 39310 22278 39362 22330
rect 39374 22278 39426 22330
rect 39438 22278 39490 22330
rect 49246 22278 49298 22330
rect 49310 22278 49362 22330
rect 49374 22278 49426 22330
rect 49438 22278 49490 22330
rect 59246 22278 59298 22330
rect 59310 22278 59362 22330
rect 59374 22278 59426 22330
rect 59438 22278 59490 22330
rect 8576 22176 8628 22228
rect 30104 22219 30156 22228
rect 30104 22185 30113 22219
rect 30113 22185 30147 22219
rect 30147 22185 30156 22219
rect 30104 22176 30156 22185
rect 37832 22176 37884 22228
rect 11796 22040 11848 22092
rect 18880 22040 18932 22092
rect 22100 21836 22152 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 14246 21734 14298 21786
rect 14310 21734 14362 21786
rect 14374 21734 14426 21786
rect 14438 21734 14490 21786
rect 24246 21734 24298 21786
rect 24310 21734 24362 21786
rect 24374 21734 24426 21786
rect 24438 21734 24490 21786
rect 34246 21734 34298 21786
rect 34310 21734 34362 21786
rect 34374 21734 34426 21786
rect 34438 21734 34490 21786
rect 44246 21734 44298 21786
rect 44310 21734 44362 21786
rect 44374 21734 44426 21786
rect 44438 21734 44490 21786
rect 54246 21734 54298 21786
rect 54310 21734 54362 21786
rect 54374 21734 54426 21786
rect 54438 21734 54490 21786
rect 64246 21734 64298 21786
rect 64310 21734 64362 21786
rect 64374 21734 64426 21786
rect 64438 21734 64490 21786
rect 67272 21675 67324 21684
rect 67272 21641 67281 21675
rect 67281 21641 67315 21675
rect 67315 21641 67324 21675
rect 67272 21632 67324 21641
rect 15016 21564 15068 21616
rect 36912 21564 36964 21616
rect 38752 21564 38804 21616
rect 56232 21564 56284 21616
rect 68100 21607 68152 21616
rect 68100 21573 68109 21607
rect 68109 21573 68143 21607
rect 68143 21573 68152 21607
rect 68100 21564 68152 21573
rect 23940 21496 23992 21548
rect 62672 21496 62724 21548
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 11980 21428 12032 21480
rect 25596 21428 25648 21480
rect 39764 21428 39816 21480
rect 67272 21428 67324 21480
rect 39856 21360 39908 21412
rect 55404 21360 55456 21412
rect 67088 21360 67140 21412
rect 47860 21292 47912 21344
rect 9246 21190 9298 21242
rect 9310 21190 9362 21242
rect 9374 21190 9426 21242
rect 9438 21190 9490 21242
rect 19246 21190 19298 21242
rect 19310 21190 19362 21242
rect 19374 21190 19426 21242
rect 19438 21190 19490 21242
rect 29246 21190 29298 21242
rect 29310 21190 29362 21242
rect 29374 21190 29426 21242
rect 29438 21190 29490 21242
rect 39246 21190 39298 21242
rect 39310 21190 39362 21242
rect 39374 21190 39426 21242
rect 39438 21190 39490 21242
rect 49246 21190 49298 21242
rect 49310 21190 49362 21242
rect 49374 21190 49426 21242
rect 49438 21190 49490 21242
rect 59246 21190 59298 21242
rect 59310 21190 59362 21242
rect 59374 21190 59426 21242
rect 59438 21190 59490 21242
rect 1400 21131 1452 21140
rect 1400 21097 1409 21131
rect 1409 21097 1443 21131
rect 1443 21097 1452 21131
rect 1400 21088 1452 21097
rect 57980 20952 58032 21004
rect 60924 20952 60976 21004
rect 52552 20816 52604 20868
rect 38844 20748 38896 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 14246 20646 14298 20698
rect 14310 20646 14362 20698
rect 14374 20646 14426 20698
rect 14438 20646 14490 20698
rect 24246 20646 24298 20698
rect 24310 20646 24362 20698
rect 24374 20646 24426 20698
rect 24438 20646 24490 20698
rect 34246 20646 34298 20698
rect 34310 20646 34362 20698
rect 34374 20646 34426 20698
rect 34438 20646 34490 20698
rect 44246 20646 44298 20698
rect 44310 20646 44362 20698
rect 44374 20646 44426 20698
rect 44438 20646 44490 20698
rect 54246 20646 54298 20698
rect 54310 20646 54362 20698
rect 54374 20646 54426 20698
rect 54438 20646 54490 20698
rect 64246 20646 64298 20698
rect 64310 20646 64362 20698
rect 64374 20646 64426 20698
rect 64438 20646 64490 20698
rect 27804 20587 27856 20596
rect 27804 20553 27813 20587
rect 27813 20553 27847 20587
rect 27847 20553 27856 20587
rect 27804 20544 27856 20553
rect 31116 20544 31168 20596
rect 29000 20340 29052 20392
rect 67088 20340 67140 20392
rect 68100 20383 68152 20392
rect 68100 20349 68109 20383
rect 68109 20349 68143 20383
rect 68143 20349 68152 20383
rect 68100 20340 68152 20349
rect 9246 20102 9298 20154
rect 9310 20102 9362 20154
rect 9374 20102 9426 20154
rect 9438 20102 9490 20154
rect 19246 20102 19298 20154
rect 19310 20102 19362 20154
rect 19374 20102 19426 20154
rect 19438 20102 19490 20154
rect 29246 20102 29298 20154
rect 29310 20102 29362 20154
rect 29374 20102 29426 20154
rect 29438 20102 29490 20154
rect 39246 20102 39298 20154
rect 39310 20102 39362 20154
rect 39374 20102 39426 20154
rect 39438 20102 39490 20154
rect 49246 20102 49298 20154
rect 49310 20102 49362 20154
rect 49374 20102 49426 20154
rect 49438 20102 49490 20154
rect 59246 20102 59298 20154
rect 59310 20102 59362 20154
rect 59374 20102 59426 20154
rect 59438 20102 59490 20154
rect 1860 20043 1912 20052
rect 1860 20009 1869 20043
rect 1869 20009 1903 20043
rect 1903 20009 1912 20043
rect 1860 20000 1912 20009
rect 27252 20043 27304 20052
rect 27252 20009 27261 20043
rect 27261 20009 27295 20043
rect 27295 20009 27304 20043
rect 27252 20000 27304 20009
rect 14832 19864 14884 19916
rect 30104 20000 30156 20052
rect 32404 19932 32456 19984
rect 50068 19932 50120 19984
rect 31852 19907 31904 19916
rect 27804 19796 27856 19848
rect 31852 19873 31861 19907
rect 31861 19873 31895 19907
rect 31895 19873 31904 19907
rect 31852 19864 31904 19873
rect 36636 19796 36688 19848
rect 5080 19660 5132 19712
rect 28264 19703 28316 19712
rect 28264 19669 28273 19703
rect 28273 19669 28307 19703
rect 28307 19669 28316 19703
rect 31116 19728 31168 19780
rect 28264 19660 28316 19669
rect 31668 19660 31720 19712
rect 33968 19703 34020 19712
rect 33968 19669 33977 19703
rect 33977 19669 34011 19703
rect 34011 19669 34020 19703
rect 33968 19660 34020 19669
rect 50344 19660 50396 19712
rect 53288 19703 53340 19712
rect 53288 19669 53297 19703
rect 53297 19669 53331 19703
rect 53331 19669 53340 19703
rect 53288 19660 53340 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 14246 19558 14298 19610
rect 14310 19558 14362 19610
rect 14374 19558 14426 19610
rect 14438 19558 14490 19610
rect 24246 19558 24298 19610
rect 24310 19558 24362 19610
rect 24374 19558 24426 19610
rect 24438 19558 24490 19610
rect 34246 19558 34298 19610
rect 34310 19558 34362 19610
rect 34374 19558 34426 19610
rect 34438 19558 34490 19610
rect 44246 19558 44298 19610
rect 44310 19558 44362 19610
rect 44374 19558 44426 19610
rect 44438 19558 44490 19610
rect 54246 19558 54298 19610
rect 54310 19558 54362 19610
rect 54374 19558 54426 19610
rect 54438 19558 54490 19610
rect 64246 19558 64298 19610
rect 64310 19558 64362 19610
rect 64374 19558 64426 19610
rect 64438 19558 64490 19610
rect 18236 19456 18288 19508
rect 28264 19456 28316 19508
rect 61660 19320 61712 19372
rect 41328 19116 41380 19168
rect 68100 19227 68152 19236
rect 68100 19193 68109 19227
rect 68109 19193 68143 19227
rect 68143 19193 68152 19227
rect 68100 19184 68152 19193
rect 9246 19014 9298 19066
rect 9310 19014 9362 19066
rect 9374 19014 9426 19066
rect 9438 19014 9490 19066
rect 39246 19014 39298 19066
rect 39310 19014 39362 19066
rect 39374 19014 39426 19066
rect 39438 19014 39490 19066
rect 49246 19014 49298 19066
rect 49310 19014 49362 19066
rect 49374 19014 49426 19066
rect 49438 19014 49490 19066
rect 59246 19014 59298 19066
rect 59310 19014 59362 19066
rect 59374 19014 59426 19066
rect 59438 19014 59490 19066
rect 2228 18912 2280 18964
rect 15108 18912 15160 18964
rect 26332 18912 26384 18964
rect 33232 18912 33284 18964
rect 50528 18912 50580 18964
rect 16396 18844 16448 18896
rect 33968 18844 34020 18896
rect 13912 18776 13964 18828
rect 38936 18776 38988 18828
rect 50804 18776 50856 18828
rect 18328 18708 18380 18760
rect 45008 18708 45060 18760
rect 1768 18683 1820 18692
rect 1768 18649 1777 18683
rect 1777 18649 1811 18683
rect 1811 18649 1820 18683
rect 1768 18640 1820 18649
rect 2872 18640 2924 18692
rect 66076 18640 66128 18692
rect 8392 18572 8444 18624
rect 15752 18572 15804 18624
rect 48412 18572 48464 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 14246 18470 14298 18522
rect 14310 18470 14362 18522
rect 14374 18470 14426 18522
rect 14438 18470 14490 18522
rect 44246 18470 44298 18522
rect 44310 18470 44362 18522
rect 44374 18470 44426 18522
rect 44438 18470 44490 18522
rect 54246 18470 54298 18522
rect 54310 18470 54362 18522
rect 54374 18470 54426 18522
rect 54438 18470 54490 18522
rect 64246 18470 64298 18522
rect 64310 18470 64362 18522
rect 64374 18470 64426 18522
rect 64438 18470 64490 18522
rect 18236 18411 18288 18420
rect 18236 18377 18245 18411
rect 18245 18377 18279 18411
rect 18279 18377 18288 18411
rect 18236 18368 18288 18377
rect 61476 18411 61528 18420
rect 61476 18377 61485 18411
rect 61485 18377 61519 18411
rect 61519 18377 61528 18411
rect 61476 18368 61528 18377
rect 17868 18096 17920 18148
rect 34612 18096 34664 18148
rect 9246 17926 9298 17978
rect 9310 17926 9362 17978
rect 9374 17926 9426 17978
rect 9438 17926 9490 17978
rect 39246 17926 39298 17978
rect 39310 17926 39362 17978
rect 39374 17926 39426 17978
rect 39438 17926 39490 17978
rect 49246 17926 49298 17978
rect 49310 17926 49362 17978
rect 49374 17926 49426 17978
rect 49438 17926 49490 17978
rect 59246 17926 59298 17978
rect 59310 17926 59362 17978
rect 59374 17926 59426 17978
rect 59438 17926 59490 17978
rect 17776 17867 17828 17876
rect 17776 17833 17785 17867
rect 17785 17833 17819 17867
rect 17819 17833 17828 17867
rect 17776 17824 17828 17833
rect 66628 17824 66680 17876
rect 18236 17756 18288 17808
rect 17868 17731 17920 17740
rect 17868 17697 17877 17731
rect 17877 17697 17911 17731
rect 17911 17697 17920 17731
rect 17868 17688 17920 17697
rect 68100 17731 68152 17740
rect 68100 17697 68109 17731
rect 68109 17697 68143 17731
rect 68143 17697 68152 17731
rect 68100 17688 68152 17697
rect 17224 17620 17276 17672
rect 29000 17620 29052 17672
rect 11152 17552 11204 17604
rect 48504 17552 48556 17604
rect 18144 17484 18196 17536
rect 37004 17484 37056 17536
rect 56048 17484 56100 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 14246 17382 14298 17434
rect 14310 17382 14362 17434
rect 14374 17382 14426 17434
rect 14438 17382 14490 17434
rect 44246 17382 44298 17434
rect 44310 17382 44362 17434
rect 44374 17382 44426 17434
rect 44438 17382 44490 17434
rect 54246 17382 54298 17434
rect 54310 17382 54362 17434
rect 54374 17382 54426 17434
rect 54438 17382 54490 17434
rect 64246 17382 64298 17434
rect 64310 17382 64362 17434
rect 64374 17382 64426 17434
rect 64438 17382 64490 17434
rect 15844 17280 15896 17332
rect 65800 17280 65852 17332
rect 10232 17212 10284 17264
rect 63500 17212 63552 17264
rect 53932 17076 53984 17128
rect 42524 17008 42576 17060
rect 54944 17008 54996 17060
rect 63868 16940 63920 16992
rect 9246 16838 9298 16890
rect 9310 16838 9362 16890
rect 9374 16838 9426 16890
rect 9438 16838 9490 16890
rect 39246 16838 39298 16890
rect 39310 16838 39362 16890
rect 39374 16838 39426 16890
rect 39438 16838 39490 16890
rect 49246 16838 49298 16890
rect 49310 16838 49362 16890
rect 49374 16838 49426 16890
rect 49438 16838 49490 16890
rect 59246 16838 59298 16890
rect 59310 16838 59362 16890
rect 59374 16838 59426 16890
rect 59438 16838 59490 16890
rect 50712 16668 50764 16720
rect 56140 16600 56192 16652
rect 68100 16643 68152 16652
rect 68100 16609 68109 16643
rect 68109 16609 68143 16643
rect 68143 16609 68152 16643
rect 68100 16600 68152 16609
rect 27620 16575 27672 16584
rect 27620 16541 27629 16575
rect 27629 16541 27663 16575
rect 27663 16541 27672 16575
rect 27620 16532 27672 16541
rect 56508 16507 56560 16516
rect 56508 16473 56517 16507
rect 56517 16473 56551 16507
rect 56551 16473 56560 16507
rect 56508 16464 56560 16473
rect 63500 16396 63552 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 14246 16294 14298 16346
rect 14310 16294 14362 16346
rect 14374 16294 14426 16346
rect 14438 16294 14490 16346
rect 44246 16294 44298 16346
rect 44310 16294 44362 16346
rect 44374 16294 44426 16346
rect 44438 16294 44490 16346
rect 54246 16294 54298 16346
rect 54310 16294 54362 16346
rect 54374 16294 54426 16346
rect 54438 16294 54490 16346
rect 64246 16294 64298 16346
rect 64310 16294 64362 16346
rect 64374 16294 64426 16346
rect 64438 16294 64490 16346
rect 18052 16235 18104 16244
rect 18052 16201 18061 16235
rect 18061 16201 18095 16235
rect 18095 16201 18104 16235
rect 18052 16192 18104 16201
rect 56140 16235 56192 16244
rect 56140 16201 56149 16235
rect 56149 16201 56183 16235
rect 56183 16201 56192 16235
rect 56140 16192 56192 16201
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 66996 15988 67048 16040
rect 17316 15852 17368 15904
rect 32588 15852 32640 15904
rect 47584 15852 47636 15904
rect 50620 15852 50672 15904
rect 56140 15852 56192 15904
rect 9246 15750 9298 15802
rect 9310 15750 9362 15802
rect 9374 15750 9426 15802
rect 9438 15750 9490 15802
rect 39246 15750 39298 15802
rect 39310 15750 39362 15802
rect 39374 15750 39426 15802
rect 39438 15750 39490 15802
rect 49246 15750 49298 15802
rect 49310 15750 49362 15802
rect 49374 15750 49426 15802
rect 49438 15750 49490 15802
rect 59246 15750 59298 15802
rect 59310 15750 59362 15802
rect 59374 15750 59426 15802
rect 59438 15750 59490 15802
rect 11244 15648 11296 15700
rect 67732 15691 67784 15700
rect 67732 15657 67741 15691
rect 67741 15657 67775 15691
rect 67775 15657 67784 15691
rect 67732 15648 67784 15657
rect 2136 15512 2188 15564
rect 10784 15512 10836 15564
rect 17408 15512 17460 15564
rect 11888 15308 11940 15360
rect 12256 15308 12308 15360
rect 18236 15351 18288 15360
rect 18236 15317 18245 15351
rect 18245 15317 18279 15351
rect 18279 15317 18288 15351
rect 18236 15308 18288 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 14246 15206 14298 15258
rect 14310 15206 14362 15258
rect 14374 15206 14426 15258
rect 14438 15206 14490 15258
rect 44246 15206 44298 15258
rect 44310 15206 44362 15258
rect 44374 15206 44426 15258
rect 44438 15206 44490 15258
rect 54246 15206 54298 15258
rect 54310 15206 54362 15258
rect 54374 15206 54426 15258
rect 54438 15206 54490 15258
rect 64246 15206 64298 15258
rect 64310 15206 64362 15258
rect 64374 15206 64426 15258
rect 64438 15206 64490 15258
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 68100 15011 68152 15020
rect 68100 14977 68109 15011
rect 68109 14977 68143 15011
rect 68143 14977 68152 15011
rect 68100 14968 68152 14977
rect 53748 14900 53800 14952
rect 67180 14943 67232 14952
rect 67180 14909 67189 14943
rect 67189 14909 67223 14943
rect 67223 14909 67232 14943
rect 67180 14900 67232 14909
rect 67732 14900 67784 14952
rect 4712 14832 4764 14884
rect 18512 14832 18564 14884
rect 1860 14807 1912 14816
rect 1860 14773 1869 14807
rect 1869 14773 1903 14807
rect 1903 14773 1912 14807
rect 1860 14764 1912 14773
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 18788 14764 18840 14816
rect 9246 14662 9298 14714
rect 9310 14662 9362 14714
rect 9374 14662 9426 14714
rect 9438 14662 9490 14714
rect 39246 14662 39298 14714
rect 39310 14662 39362 14714
rect 39374 14662 39426 14714
rect 39438 14662 39490 14714
rect 49246 14662 49298 14714
rect 49310 14662 49362 14714
rect 49374 14662 49426 14714
rect 49438 14662 49490 14714
rect 59246 14662 59298 14714
rect 59310 14662 59362 14714
rect 59374 14662 59426 14714
rect 59438 14662 59490 14714
rect 16028 14560 16080 14612
rect 17132 14560 17184 14612
rect 17316 14603 17368 14612
rect 17316 14569 17325 14603
rect 17325 14569 17359 14603
rect 17359 14569 17368 14603
rect 17316 14560 17368 14569
rect 5632 14492 5684 14544
rect 18052 14492 18104 14544
rect 38108 14492 38160 14544
rect 48596 14492 48648 14544
rect 6736 14424 6788 14476
rect 12072 14424 12124 14476
rect 17132 14424 17184 14476
rect 18696 14424 18748 14476
rect 48780 14424 48832 14476
rect 55956 14424 56008 14476
rect 67272 14424 67324 14476
rect 48688 14356 48740 14408
rect 17408 14288 17460 14340
rect 35716 14288 35768 14340
rect 16488 14220 16540 14272
rect 17684 14220 17736 14272
rect 17960 14220 18012 14272
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 38384 14220 38436 14272
rect 51816 14220 51868 14272
rect 55864 14220 55916 14272
rect 58440 14220 58492 14272
rect 65340 14220 65392 14272
rect 67640 14220 67692 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 14246 14118 14298 14170
rect 14310 14118 14362 14170
rect 14374 14118 14426 14170
rect 14438 14118 14490 14170
rect 44246 14118 44298 14170
rect 44310 14118 44362 14170
rect 44374 14118 44426 14170
rect 44438 14118 44490 14170
rect 54246 14118 54298 14170
rect 54310 14118 54362 14170
rect 54374 14118 54426 14170
rect 54438 14118 54490 14170
rect 64246 14118 64298 14170
rect 64310 14118 64362 14170
rect 64374 14118 64426 14170
rect 64438 14118 64490 14170
rect 13084 14016 13136 14068
rect 17592 14016 17644 14068
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 14648 13991 14700 14000
rect 14648 13957 14657 13991
rect 14657 13957 14691 13991
rect 14691 13957 14700 13991
rect 14648 13948 14700 13957
rect 55128 14016 55180 14068
rect 66444 14016 66496 14068
rect 38108 13991 38160 14000
rect 38108 13957 38117 13991
rect 38117 13957 38151 13991
rect 38151 13957 38160 13991
rect 38108 13948 38160 13957
rect 38568 13948 38620 14000
rect 39764 13948 39816 14000
rect 46204 13948 46256 14000
rect 14096 13812 14148 13864
rect 15660 13812 15712 13864
rect 15844 13855 15896 13864
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 16304 13855 16356 13864
rect 15844 13812 15896 13821
rect 16304 13821 16313 13855
rect 16313 13821 16347 13855
rect 16347 13821 16356 13855
rect 16304 13812 16356 13821
rect 47400 13880 47452 13932
rect 17132 13812 17184 13864
rect 17592 13855 17644 13864
rect 17592 13821 17601 13855
rect 17601 13821 17635 13855
rect 17635 13821 17644 13855
rect 17592 13812 17644 13821
rect 18604 13812 18656 13864
rect 37648 13812 37700 13864
rect 37924 13812 37976 13864
rect 39764 13855 39816 13864
rect 39764 13821 39773 13855
rect 39773 13821 39807 13855
rect 39807 13821 39816 13855
rect 39764 13812 39816 13821
rect 68100 13855 68152 13864
rect 68100 13821 68109 13855
rect 68109 13821 68143 13855
rect 68143 13821 68152 13855
rect 68100 13812 68152 13821
rect 14096 13676 14148 13728
rect 53840 13744 53892 13796
rect 9246 13574 9298 13626
rect 9310 13574 9362 13626
rect 9374 13574 9426 13626
rect 9438 13574 9490 13626
rect 39246 13574 39298 13626
rect 39310 13574 39362 13626
rect 39374 13574 39426 13626
rect 39438 13574 39490 13626
rect 49246 13574 49298 13626
rect 49310 13574 49362 13626
rect 49374 13574 49426 13626
rect 49438 13574 49490 13626
rect 59246 13574 59298 13626
rect 59310 13574 59362 13626
rect 59374 13574 59426 13626
rect 59438 13574 59490 13626
rect 1860 13515 1912 13524
rect 1860 13481 1869 13515
rect 1869 13481 1903 13515
rect 1903 13481 1912 13515
rect 1860 13472 1912 13481
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 62948 13472 63000 13524
rect 2320 13404 2372 13456
rect 2412 13404 2464 13456
rect 13360 13336 13412 13388
rect 40040 13404 40092 13456
rect 40684 13404 40736 13456
rect 41144 13404 41196 13456
rect 37464 13268 37516 13320
rect 40040 13268 40092 13320
rect 40132 13268 40184 13320
rect 55312 13336 55364 13388
rect 43168 13268 43220 13320
rect 51908 13268 51960 13320
rect 15568 13200 15620 13252
rect 16304 13200 16356 13252
rect 55680 13200 55732 13252
rect 13544 13175 13596 13184
rect 13544 13141 13553 13175
rect 13553 13141 13587 13175
rect 13587 13141 13596 13175
rect 13544 13132 13596 13141
rect 15936 13132 15988 13184
rect 16396 13132 16448 13184
rect 16764 13175 16816 13184
rect 16764 13141 16773 13175
rect 16773 13141 16807 13175
rect 16807 13141 16816 13175
rect 16764 13132 16816 13141
rect 18420 13132 18472 13184
rect 37740 13132 37792 13184
rect 39212 13175 39264 13184
rect 39212 13141 39221 13175
rect 39221 13141 39255 13175
rect 39255 13141 39264 13175
rect 39212 13132 39264 13141
rect 39672 13132 39724 13184
rect 40316 13132 40368 13184
rect 41144 13132 41196 13184
rect 41972 13132 42024 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 14246 13030 14298 13082
rect 14310 13030 14362 13082
rect 14374 13030 14426 13082
rect 14438 13030 14490 13082
rect 44246 13030 44298 13082
rect 44310 13030 44362 13082
rect 44374 13030 44426 13082
rect 44438 13030 44490 13082
rect 54246 13030 54298 13082
rect 54310 13030 54362 13082
rect 54374 13030 54426 13082
rect 54438 13030 54490 13082
rect 64246 13030 64298 13082
rect 64310 13030 64362 13082
rect 64374 13030 64426 13082
rect 64438 13030 64490 13082
rect 2320 12928 2372 12980
rect 15476 12928 15528 12980
rect 18144 12928 18196 12980
rect 38292 12928 38344 12980
rect 38752 12928 38804 12980
rect 39948 12928 40000 12980
rect 53840 12971 53892 12980
rect 53840 12937 53849 12971
rect 53849 12937 53883 12971
rect 53883 12937 53892 12971
rect 53840 12928 53892 12937
rect 15752 12903 15804 12912
rect 15752 12869 15761 12903
rect 15761 12869 15795 12903
rect 15795 12869 15804 12903
rect 15752 12860 15804 12869
rect 40960 12860 41012 12912
rect 16304 12792 16356 12844
rect 23296 12792 23348 12844
rect 37556 12792 37608 12844
rect 40316 12792 40368 12844
rect 10508 12656 10560 12708
rect 12164 12588 12216 12640
rect 12716 12588 12768 12640
rect 13360 12631 13412 12640
rect 13360 12597 13369 12631
rect 13369 12597 13403 12631
rect 13403 12597 13412 12631
rect 13360 12588 13412 12597
rect 19984 12724 20036 12776
rect 40592 12724 40644 12776
rect 42616 12860 42668 12912
rect 16120 12656 16172 12708
rect 37188 12656 37240 12708
rect 40684 12656 40736 12708
rect 53288 12792 53340 12844
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 17592 12588 17644 12640
rect 37832 12588 37884 12640
rect 39120 12588 39172 12640
rect 39580 12631 39632 12640
rect 39580 12597 39589 12631
rect 39589 12597 39623 12631
rect 39623 12597 39632 12631
rect 39580 12588 39632 12597
rect 40868 12631 40920 12640
rect 40868 12597 40877 12631
rect 40877 12597 40911 12631
rect 40911 12597 40920 12631
rect 42616 12656 42668 12708
rect 65248 12724 65300 12776
rect 40868 12588 40920 12597
rect 53932 12588 53984 12640
rect 9246 12486 9298 12538
rect 9310 12486 9362 12538
rect 9374 12486 9426 12538
rect 9438 12486 9490 12538
rect 39246 12486 39298 12538
rect 39310 12486 39362 12538
rect 39374 12486 39426 12538
rect 39438 12486 39490 12538
rect 49246 12486 49298 12538
rect 49310 12486 49362 12538
rect 49374 12486 49426 12538
rect 49438 12486 49490 12538
rect 59246 12486 59298 12538
rect 59310 12486 59362 12538
rect 59374 12486 59426 12538
rect 59438 12486 59490 12538
rect 9680 12384 9732 12436
rect 23940 12384 23992 12436
rect 12624 12359 12676 12368
rect 12624 12325 12633 12359
rect 12633 12325 12667 12359
rect 12667 12325 12676 12359
rect 12624 12316 12676 12325
rect 16580 12359 16632 12368
rect 16580 12325 16589 12359
rect 16589 12325 16623 12359
rect 16623 12325 16632 12359
rect 16580 12316 16632 12325
rect 11428 12044 11480 12096
rect 11796 12044 11848 12096
rect 16948 12248 17000 12300
rect 18236 12291 18288 12300
rect 18236 12257 18245 12291
rect 18245 12257 18279 12291
rect 18279 12257 18288 12291
rect 18236 12248 18288 12257
rect 68100 12291 68152 12300
rect 68100 12257 68109 12291
rect 68109 12257 68143 12291
rect 68143 12257 68152 12291
rect 68100 12248 68152 12257
rect 13820 12180 13872 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 18052 12180 18104 12232
rect 39764 12180 39816 12232
rect 39856 12112 39908 12164
rect 13452 12044 13504 12096
rect 14740 12044 14792 12096
rect 15016 12044 15068 12096
rect 15200 12087 15252 12096
rect 15200 12053 15209 12087
rect 15209 12053 15243 12087
rect 15243 12053 15252 12087
rect 15200 12044 15252 12053
rect 38108 12087 38160 12096
rect 38108 12053 38117 12087
rect 38117 12053 38151 12087
rect 38151 12053 38160 12087
rect 38108 12044 38160 12053
rect 38200 12044 38252 12096
rect 39120 12087 39172 12096
rect 39120 12053 39129 12087
rect 39129 12053 39163 12087
rect 39163 12053 39172 12087
rect 39120 12044 39172 12053
rect 39764 12087 39816 12096
rect 39764 12053 39773 12087
rect 39773 12053 39807 12087
rect 39807 12053 39816 12087
rect 39764 12044 39816 12053
rect 40316 12044 40368 12096
rect 40960 12087 41012 12096
rect 40960 12053 40969 12087
rect 40969 12053 41003 12087
rect 41003 12053 41012 12087
rect 40960 12044 41012 12053
rect 42708 12087 42760 12096
rect 42708 12053 42717 12087
rect 42717 12053 42751 12087
rect 42751 12053 42760 12087
rect 42708 12044 42760 12053
rect 43260 12087 43312 12096
rect 43260 12053 43269 12087
rect 43269 12053 43303 12087
rect 43303 12053 43312 12087
rect 43260 12044 43312 12053
rect 48688 12044 48740 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 14246 11942 14298 11994
rect 14310 11942 14362 11994
rect 14374 11942 14426 11994
rect 14438 11942 14490 11994
rect 44246 11942 44298 11994
rect 44310 11942 44362 11994
rect 44374 11942 44426 11994
rect 44438 11942 44490 11994
rect 54246 11942 54298 11994
rect 54310 11942 54362 11994
rect 54374 11942 54426 11994
rect 54438 11942 54490 11994
rect 64246 11942 64298 11994
rect 64310 11942 64362 11994
rect 64374 11942 64426 11994
rect 64438 11942 64490 11994
rect 38016 11883 38068 11892
rect 38016 11849 38025 11883
rect 38025 11849 38059 11883
rect 38059 11849 38068 11883
rect 38016 11840 38068 11849
rect 42156 11840 42208 11892
rect 45652 11840 45704 11892
rect 38108 11772 38160 11824
rect 53012 11772 53064 11824
rect 62120 11772 62172 11824
rect 65064 11772 65116 11824
rect 45560 11704 45612 11756
rect 53196 11704 53248 11756
rect 38292 11636 38344 11688
rect 38660 11636 38712 11688
rect 9956 11568 10008 11620
rect 42248 11568 42300 11620
rect 42432 11568 42484 11620
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 11980 11500 12032 11552
rect 12348 11500 12400 11552
rect 12624 11500 12676 11552
rect 12992 11500 13044 11552
rect 14832 11500 14884 11552
rect 14924 11543 14976 11552
rect 14924 11509 14933 11543
rect 14933 11509 14967 11543
rect 14967 11509 14976 11543
rect 14924 11500 14976 11509
rect 15660 11500 15712 11552
rect 16488 11500 16540 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 17684 11543 17736 11552
rect 17684 11509 17693 11543
rect 17693 11509 17727 11543
rect 17727 11509 17736 11543
rect 17684 11500 17736 11509
rect 18052 11500 18104 11552
rect 38476 11500 38528 11552
rect 40132 11500 40184 11552
rect 40500 11500 40552 11552
rect 41052 11543 41104 11552
rect 41052 11509 41061 11543
rect 41061 11509 41095 11543
rect 41095 11509 41104 11543
rect 41052 11500 41104 11509
rect 42892 11500 42944 11552
rect 67180 11636 67232 11688
rect 45560 11568 45612 11620
rect 45652 11568 45704 11620
rect 57704 11568 57756 11620
rect 44640 11543 44692 11552
rect 44640 11509 44649 11543
rect 44649 11509 44683 11543
rect 44683 11509 44692 11543
rect 44640 11500 44692 11509
rect 65984 11500 66036 11552
rect 66352 11500 66404 11552
rect 66628 11543 66680 11552
rect 66628 11509 66637 11543
rect 66637 11509 66671 11543
rect 66671 11509 66680 11543
rect 66628 11500 66680 11509
rect 67088 11500 67140 11552
rect 67364 11500 67416 11552
rect 67640 11543 67692 11552
rect 67640 11509 67649 11543
rect 67649 11509 67683 11543
rect 67683 11509 67692 11543
rect 67640 11500 67692 11509
rect 9246 11398 9298 11450
rect 9310 11398 9362 11450
rect 9374 11398 9426 11450
rect 9438 11398 9490 11450
rect 39246 11398 39298 11450
rect 39310 11398 39362 11450
rect 39374 11398 39426 11450
rect 39438 11398 39490 11450
rect 49246 11398 49298 11450
rect 49310 11398 49362 11450
rect 49374 11398 49426 11450
rect 49438 11398 49490 11450
rect 59246 11398 59298 11450
rect 59310 11398 59362 11450
rect 59374 11398 59426 11450
rect 59438 11398 59490 11450
rect 67272 11339 67324 11348
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 9680 11160 9732 11212
rect 13360 11228 13412 11280
rect 15108 11160 15160 11212
rect 37924 11203 37976 11212
rect 37924 11169 37933 11203
rect 37933 11169 37967 11203
rect 37967 11169 37976 11203
rect 37924 11160 37976 11169
rect 39764 11160 39816 11212
rect 10968 11092 11020 11144
rect 10600 11024 10652 11076
rect 10876 11067 10928 11076
rect 10876 11033 10885 11067
rect 10885 11033 10919 11067
rect 10919 11033 10928 11067
rect 10876 11024 10928 11033
rect 11704 11024 11756 11076
rect 12716 11024 12768 11076
rect 13268 11024 13320 11076
rect 13912 11024 13964 11076
rect 15384 11024 15436 11076
rect 15476 11024 15528 11076
rect 16672 11024 16724 11076
rect 17132 11067 17184 11076
rect 17132 11033 17141 11067
rect 17141 11033 17175 11067
rect 17175 11033 17184 11067
rect 17132 11024 17184 11033
rect 17776 11067 17828 11076
rect 17776 11033 17785 11067
rect 17785 11033 17819 11067
rect 17819 11033 17828 11067
rect 17776 11024 17828 11033
rect 38108 11024 38160 11076
rect 38752 11024 38804 11076
rect 39764 11067 39816 11076
rect 39764 11033 39773 11067
rect 39773 11033 39807 11067
rect 39807 11033 39816 11067
rect 39764 11024 39816 11033
rect 39672 10956 39724 11008
rect 67272 11305 67281 11339
rect 67281 11305 67315 11339
rect 67315 11305 67324 11339
rect 67272 11296 67324 11305
rect 67640 11160 67692 11212
rect 42432 11092 42484 11144
rect 40040 11024 40092 11076
rect 40868 11024 40920 11076
rect 41420 11024 41472 11076
rect 42064 11067 42116 11076
rect 42064 11033 42073 11067
rect 42073 11033 42107 11067
rect 42107 11033 42116 11067
rect 42064 11024 42116 11033
rect 42156 11024 42208 11076
rect 42616 11067 42668 11076
rect 42616 11033 42625 11067
rect 42625 11033 42659 11067
rect 42659 11033 42668 11067
rect 42616 11024 42668 11033
rect 42708 11024 42760 11076
rect 43812 11067 43864 11076
rect 43812 11033 43821 11067
rect 43821 11033 43855 11067
rect 43855 11033 43864 11067
rect 43812 11024 43864 11033
rect 44548 11024 44600 11076
rect 51264 11092 51316 11144
rect 65432 11092 65484 11144
rect 66536 11092 66588 11144
rect 45100 11024 45152 11076
rect 45468 11024 45520 11076
rect 65892 11024 65944 11076
rect 66076 11067 66128 11076
rect 66076 11033 66085 11067
rect 66085 11033 66119 11067
rect 66119 11033 66128 11067
rect 66076 11024 66128 11033
rect 66812 11067 66864 11076
rect 66812 11033 66821 11067
rect 66821 11033 66855 11067
rect 66855 11033 66864 11067
rect 66812 11024 66864 11033
rect 68100 11067 68152 11076
rect 68100 11033 68109 11067
rect 68109 11033 68143 11067
rect 68143 11033 68152 11067
rect 68100 11024 68152 11033
rect 42340 10956 42392 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 14246 10854 14298 10906
rect 14310 10854 14362 10906
rect 14374 10854 14426 10906
rect 14438 10854 14490 10906
rect 44246 10854 44298 10906
rect 44310 10854 44362 10906
rect 44374 10854 44426 10906
rect 44438 10854 44490 10906
rect 54246 10854 54298 10906
rect 54310 10854 54362 10906
rect 54374 10854 54426 10906
rect 54438 10854 54490 10906
rect 64246 10854 64298 10906
rect 64310 10854 64362 10906
rect 64374 10854 64426 10906
rect 64438 10854 64490 10906
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 18236 10795 18288 10804
rect 18236 10761 18245 10795
rect 18245 10761 18279 10795
rect 18279 10761 18288 10795
rect 18236 10752 18288 10761
rect 14464 10684 14516 10736
rect 4804 10616 4856 10668
rect 12256 10616 12308 10668
rect 43996 10616 44048 10668
rect 51356 10684 51408 10736
rect 17224 10548 17276 10600
rect 37372 10548 37424 10600
rect 37740 10548 37792 10600
rect 38016 10548 38068 10600
rect 38568 10548 38620 10600
rect 42524 10548 42576 10600
rect 67456 10548 67508 10600
rect 8484 10480 8536 10532
rect 10692 10480 10744 10532
rect 11336 10480 11388 10532
rect 13084 10480 13136 10532
rect 15200 10480 15252 10532
rect 44824 10480 44876 10532
rect 45008 10480 45060 10532
rect 8668 10412 8720 10464
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 11244 10412 11296 10464
rect 12900 10412 12952 10464
rect 13820 10412 13872 10464
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 15844 10412 15896 10464
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 37924 10412 37976 10464
rect 38568 10412 38620 10464
rect 39028 10412 39080 10464
rect 40132 10412 40184 10464
rect 40776 10455 40828 10464
rect 40776 10421 40785 10455
rect 40785 10421 40819 10455
rect 40819 10421 40828 10455
rect 40776 10412 40828 10421
rect 41512 10412 41564 10464
rect 41880 10455 41932 10464
rect 41880 10421 41889 10455
rect 41889 10421 41923 10455
rect 41923 10421 41932 10455
rect 41880 10412 41932 10421
rect 42984 10455 43036 10464
rect 42984 10421 42993 10455
rect 42993 10421 43027 10455
rect 43027 10421 43036 10455
rect 42984 10412 43036 10421
rect 43536 10455 43588 10464
rect 43536 10421 43545 10455
rect 43545 10421 43579 10455
rect 43579 10421 43588 10455
rect 43536 10412 43588 10421
rect 44180 10455 44232 10464
rect 44180 10421 44189 10455
rect 44189 10421 44223 10455
rect 44223 10421 44232 10455
rect 44180 10412 44232 10421
rect 45100 10412 45152 10464
rect 46480 10412 46532 10464
rect 47676 10412 47728 10464
rect 64144 10480 64196 10532
rect 66168 10523 66220 10532
rect 66168 10489 66177 10523
rect 66177 10489 66211 10523
rect 66211 10489 66220 10523
rect 66168 10480 66220 10489
rect 67548 10480 67600 10532
rect 64696 10412 64748 10464
rect 64880 10412 64932 10464
rect 65524 10412 65576 10464
rect 65708 10412 65760 10464
rect 67180 10412 67232 10464
rect 68008 10455 68060 10464
rect 68008 10421 68017 10455
rect 68017 10421 68051 10455
rect 68051 10421 68060 10455
rect 68008 10412 68060 10421
rect 9246 10310 9298 10362
rect 9310 10310 9362 10362
rect 9374 10310 9426 10362
rect 9438 10310 9490 10362
rect 39246 10310 39298 10362
rect 39310 10310 39362 10362
rect 39374 10310 39426 10362
rect 39438 10310 39490 10362
rect 49246 10310 49298 10362
rect 49310 10310 49362 10362
rect 49374 10310 49426 10362
rect 49438 10310 49490 10362
rect 59246 10310 59298 10362
rect 59310 10310 59362 10362
rect 59374 10310 59426 10362
rect 59438 10310 59490 10362
rect 2412 10208 2464 10260
rect 14096 10208 14148 10260
rect 15292 10208 15344 10260
rect 16212 10140 16264 10192
rect 39396 10140 39448 10192
rect 39672 10140 39724 10192
rect 12532 10072 12584 10124
rect 14464 10072 14516 10124
rect 15200 10115 15252 10124
rect 15200 10081 15209 10115
rect 15209 10081 15243 10115
rect 15243 10081 15252 10115
rect 15200 10072 15252 10081
rect 18328 10072 18380 10124
rect 32680 10072 32732 10124
rect 37832 10072 37884 10124
rect 11612 10004 11664 10056
rect 36084 10004 36136 10056
rect 37188 10004 37240 10056
rect 47032 10208 47084 10260
rect 45100 10140 45152 10192
rect 64972 10140 65024 10192
rect 67640 10140 67692 10192
rect 44088 10115 44140 10124
rect 44088 10081 44097 10115
rect 44097 10081 44131 10115
rect 44131 10081 44140 10115
rect 44088 10072 44140 10081
rect 63776 10072 63828 10124
rect 63960 10072 64012 10124
rect 12532 9936 12584 9988
rect 18328 9936 18380 9988
rect 38292 9936 38344 9988
rect 41696 10004 41748 10056
rect 42524 10004 42576 10056
rect 44916 10004 44968 10056
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2780 9868 2832 9877
rect 3700 9868 3752 9920
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 5172 9868 5224 9920
rect 5448 9868 5500 9920
rect 6368 9868 6420 9920
rect 6736 9868 6788 9920
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 9772 9911 9824 9920
rect 9772 9877 9781 9911
rect 9781 9877 9815 9911
rect 9815 9877 9824 9911
rect 9772 9868 9824 9877
rect 10232 9868 10284 9920
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 11612 9868 11664 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 15568 9868 15620 9920
rect 16580 9868 16632 9920
rect 18144 9868 18196 9920
rect 32588 9868 32640 9920
rect 41236 9936 41288 9988
rect 45284 9936 45336 9988
rect 65800 9936 65852 9988
rect 66904 9936 66956 9988
rect 68100 9979 68152 9988
rect 68100 9945 68109 9979
rect 68109 9945 68143 9979
rect 68143 9945 68152 9979
rect 68100 9936 68152 9945
rect 39488 9868 39540 9920
rect 40868 9868 40920 9920
rect 41144 9911 41196 9920
rect 41144 9877 41153 9911
rect 41153 9877 41187 9911
rect 41187 9877 41196 9911
rect 41144 9868 41196 9877
rect 41696 9911 41748 9920
rect 41696 9877 41705 9911
rect 41705 9877 41739 9911
rect 41739 9877 41748 9911
rect 41696 9868 41748 9877
rect 42156 9868 42208 9920
rect 42800 9911 42852 9920
rect 42800 9877 42809 9911
rect 42809 9877 42843 9911
rect 42843 9877 42852 9911
rect 42800 9868 42852 9877
rect 43352 9911 43404 9920
rect 43352 9877 43361 9911
rect 43361 9877 43395 9911
rect 43395 9877 43404 9911
rect 43352 9868 43404 9877
rect 44916 9868 44968 9920
rect 46296 9911 46348 9920
rect 46296 9877 46305 9911
rect 46305 9877 46339 9911
rect 46339 9877 46348 9911
rect 46296 9868 46348 9877
rect 46756 9911 46808 9920
rect 46756 9877 46765 9911
rect 46765 9877 46799 9911
rect 46799 9877 46808 9911
rect 46756 9868 46808 9877
rect 47768 9868 47820 9920
rect 63960 9911 64012 9920
rect 63960 9877 63969 9911
rect 63969 9877 64003 9911
rect 64003 9877 64012 9911
rect 63960 9868 64012 9877
rect 64972 9868 65024 9920
rect 65892 9868 65944 9920
rect 66996 9911 67048 9920
rect 66996 9877 67005 9911
rect 67005 9877 67039 9911
rect 67039 9877 67048 9911
rect 66996 9868 67048 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 14246 9766 14298 9818
rect 14310 9766 14362 9818
rect 14374 9766 14426 9818
rect 14438 9766 14490 9818
rect 44246 9766 44298 9818
rect 44310 9766 44362 9818
rect 44374 9766 44426 9818
rect 44438 9766 44490 9818
rect 54246 9766 54298 9818
rect 54310 9766 54362 9818
rect 54374 9766 54426 9818
rect 54438 9766 54490 9818
rect 64246 9766 64298 9818
rect 64310 9766 64362 9818
rect 64374 9766 64426 9818
rect 64438 9766 64490 9818
rect 6552 9664 6604 9716
rect 13084 9664 13136 9716
rect 14832 9664 14884 9716
rect 15200 9664 15252 9716
rect 39764 9664 39816 9716
rect 41328 9664 41380 9716
rect 1768 9639 1820 9648
rect 1768 9605 1777 9639
rect 1777 9605 1811 9639
rect 1811 9605 1820 9639
rect 1768 9596 1820 9605
rect 2596 9639 2648 9648
rect 2596 9605 2605 9639
rect 2605 9605 2639 9639
rect 2639 9605 2648 9639
rect 2596 9596 2648 9605
rect 5080 9596 5132 9648
rect 18880 9596 18932 9648
rect 37740 9596 37792 9648
rect 38016 9596 38068 9648
rect 2412 9460 2464 9512
rect 23940 9528 23992 9580
rect 4160 9460 4212 9512
rect 4804 9460 4856 9512
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 5816 9460 5868 9512
rect 6828 9460 6880 9512
rect 9680 9460 9732 9512
rect 11980 9460 12032 9512
rect 13820 9460 13872 9512
rect 14924 9460 14976 9512
rect 15200 9460 15252 9512
rect 15476 9460 15528 9512
rect 17500 9460 17552 9512
rect 13636 9392 13688 9444
rect 37280 9460 37332 9512
rect 4988 9324 5040 9376
rect 5264 9324 5316 9376
rect 5632 9324 5684 9376
rect 6644 9324 6696 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8392 9324 8444 9376
rect 8760 9324 8812 9376
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 13176 9324 13228 9376
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 15476 9324 15528 9376
rect 16212 9324 16264 9376
rect 23848 9392 23900 9444
rect 39120 9460 39172 9512
rect 43904 9528 43956 9580
rect 44088 9528 44140 9580
rect 39396 9503 39448 9512
rect 39396 9469 39405 9503
rect 39405 9469 39439 9503
rect 39439 9469 39448 9503
rect 39396 9460 39448 9469
rect 18236 9324 18288 9376
rect 38016 9324 38068 9376
rect 40316 9460 40368 9512
rect 41236 9460 41288 9512
rect 42064 9460 42116 9512
rect 43168 9460 43220 9512
rect 45376 9460 45428 9512
rect 44824 9392 44876 9444
rect 46020 9392 46072 9444
rect 46388 9392 46440 9444
rect 48596 9392 48648 9444
rect 48872 9392 48924 9444
rect 40316 9324 40368 9376
rect 40500 9324 40552 9376
rect 41604 9324 41656 9376
rect 42064 9367 42116 9376
rect 42064 9333 42073 9367
rect 42073 9333 42107 9367
rect 42107 9333 42116 9367
rect 42064 9324 42116 9333
rect 43076 9324 43128 9376
rect 44732 9367 44784 9376
rect 44732 9333 44741 9367
rect 44741 9333 44775 9367
rect 44775 9333 44784 9367
rect 44732 9324 44784 9333
rect 45192 9367 45244 9376
rect 45192 9333 45201 9367
rect 45201 9333 45235 9367
rect 45235 9333 45244 9367
rect 45192 9324 45244 9333
rect 45836 9367 45888 9376
rect 45836 9333 45845 9367
rect 45845 9333 45879 9367
rect 45879 9333 45888 9367
rect 45836 9324 45888 9333
rect 46572 9367 46624 9376
rect 46572 9333 46581 9367
rect 46581 9333 46615 9367
rect 46615 9333 46624 9367
rect 46572 9324 46624 9333
rect 48780 9324 48832 9376
rect 49148 9367 49200 9376
rect 49148 9333 49157 9367
rect 49157 9333 49191 9367
rect 49191 9333 49200 9367
rect 49148 9324 49200 9333
rect 49608 9324 49660 9376
rect 60464 9392 60516 9444
rect 68100 9392 68152 9444
rect 50252 9367 50304 9376
rect 50252 9333 50261 9367
rect 50261 9333 50295 9367
rect 50295 9333 50304 9367
rect 50252 9324 50304 9333
rect 62672 9324 62724 9376
rect 63316 9367 63368 9376
rect 63316 9333 63325 9367
rect 63325 9333 63359 9367
rect 63359 9333 63368 9367
rect 63316 9324 63368 9333
rect 63592 9324 63644 9376
rect 64236 9324 64288 9376
rect 65248 9324 65300 9376
rect 65984 9324 66036 9376
rect 66720 9367 66772 9376
rect 66720 9333 66729 9367
rect 66729 9333 66763 9367
rect 66763 9333 66772 9367
rect 66720 9324 66772 9333
rect 67272 9324 67324 9376
rect 9246 9222 9298 9274
rect 9310 9222 9362 9274
rect 9374 9222 9426 9274
rect 9438 9222 9490 9274
rect 39246 9222 39298 9274
rect 39310 9222 39362 9274
rect 39374 9222 39426 9274
rect 39438 9222 39490 9274
rect 49246 9222 49298 9274
rect 49310 9222 49362 9274
rect 49374 9222 49426 9274
rect 49438 9222 49490 9274
rect 59246 9222 59298 9274
rect 59310 9222 59362 9274
rect 59374 9222 59426 9274
rect 59438 9222 59490 9274
rect 7472 9163 7524 9172
rect 7472 9129 7481 9163
rect 7481 9129 7515 9163
rect 7515 9129 7524 9163
rect 7472 9120 7524 9129
rect 8760 9120 8812 9172
rect 17868 9120 17920 9172
rect 63684 9120 63736 9172
rect 67824 9120 67876 9172
rect 50896 9095 50948 9104
rect 13452 8984 13504 9036
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 15660 8984 15712 9036
rect 17592 9027 17644 9036
rect 17592 8993 17601 9027
rect 17601 8993 17635 9027
rect 17635 8993 17644 9027
rect 17592 8984 17644 8993
rect 24952 8984 25004 9036
rect 14096 8916 14148 8968
rect 2412 8848 2464 8900
rect 6276 8848 6328 8900
rect 7288 8848 7340 8900
rect 17224 8916 17276 8968
rect 32772 8984 32824 9036
rect 38200 8984 38252 9036
rect 39028 8984 39080 9036
rect 50896 9061 50905 9095
rect 50905 9061 50939 9095
rect 50939 9061 50948 9095
rect 50896 9052 50948 9061
rect 51356 9052 51408 9104
rect 40500 8984 40552 9036
rect 34888 8916 34940 8968
rect 41052 8916 41104 8968
rect 48412 8984 48464 9036
rect 50344 8984 50396 9036
rect 68100 9027 68152 9036
rect 68100 8993 68109 9027
rect 68109 8993 68143 9027
rect 68143 8993 68152 9027
rect 68100 8984 68152 8993
rect 68836 8984 68888 9036
rect 46848 8916 46900 8968
rect 19340 8848 19392 8900
rect 32312 8848 32364 8900
rect 37740 8848 37792 8900
rect 61384 8848 61436 8900
rect 62304 8848 62356 8900
rect 65524 8848 65576 8900
rect 67732 8848 67784 8900
rect 1400 8823 1452 8832
rect 1400 8789 1409 8823
rect 1409 8789 1443 8823
rect 1443 8789 1452 8823
rect 1400 8780 1452 8789
rect 1676 8780 1728 8832
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 2964 8780 3016 8832
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 5908 8780 5960 8832
rect 6092 8823 6144 8832
rect 6092 8789 6101 8823
rect 6101 8789 6135 8823
rect 6135 8789 6144 8823
rect 6092 8780 6144 8789
rect 7104 8780 7156 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 8852 8780 8904 8832
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 11060 8780 11112 8832
rect 13544 8780 13596 8832
rect 16856 8780 16908 8832
rect 23572 8780 23624 8832
rect 39856 8780 39908 8832
rect 41788 8823 41840 8832
rect 41788 8789 41797 8823
rect 41797 8789 41831 8823
rect 41831 8789 41840 8823
rect 41788 8780 41840 8789
rect 42340 8823 42392 8832
rect 42340 8789 42349 8823
rect 42349 8789 42383 8823
rect 42383 8789 42392 8823
rect 42340 8780 42392 8789
rect 42892 8823 42944 8832
rect 42892 8789 42901 8823
rect 42901 8789 42935 8823
rect 42935 8789 42944 8823
rect 42892 8780 42944 8789
rect 43444 8823 43496 8832
rect 43444 8789 43453 8823
rect 43453 8789 43487 8823
rect 43487 8789 43496 8823
rect 43444 8780 43496 8789
rect 43812 8780 43864 8832
rect 44548 8823 44600 8832
rect 44548 8789 44557 8823
rect 44557 8789 44591 8823
rect 44591 8789 44600 8823
rect 44548 8780 44600 8789
rect 45652 8823 45704 8832
rect 45652 8789 45661 8823
rect 45661 8789 45695 8823
rect 45695 8789 45704 8823
rect 45652 8780 45704 8789
rect 46112 8780 46164 8832
rect 46388 8780 46440 8832
rect 47032 8780 47084 8832
rect 47492 8780 47544 8832
rect 48412 8823 48464 8832
rect 48412 8789 48421 8823
rect 48421 8789 48455 8823
rect 48455 8789 48464 8823
rect 48412 8780 48464 8789
rect 49056 8780 49108 8832
rect 49700 8780 49752 8832
rect 49976 8780 50028 8832
rect 50436 8780 50488 8832
rect 51448 8780 51500 8832
rect 51632 8780 51684 8832
rect 52000 8823 52052 8832
rect 52000 8789 52009 8823
rect 52009 8789 52043 8823
rect 52043 8789 52052 8823
rect 52000 8780 52052 8789
rect 52460 8780 52512 8832
rect 53012 8780 53064 8832
rect 54116 8823 54168 8832
rect 54116 8789 54125 8823
rect 54125 8789 54159 8823
rect 54159 8789 54168 8823
rect 54116 8780 54168 8789
rect 62856 8780 62908 8832
rect 63132 8780 63184 8832
rect 63500 8823 63552 8832
rect 63500 8789 63509 8823
rect 63509 8789 63543 8823
rect 63543 8789 63552 8823
rect 63500 8780 63552 8789
rect 63776 8780 63828 8832
rect 63868 8780 63920 8832
rect 64052 8823 64104 8832
rect 64052 8789 64061 8823
rect 64061 8789 64095 8823
rect 64095 8789 64104 8823
rect 64052 8780 64104 8789
rect 65064 8823 65116 8832
rect 65064 8789 65073 8823
rect 65073 8789 65107 8823
rect 65107 8789 65116 8823
rect 65064 8780 65116 8789
rect 65432 8780 65484 8832
rect 68100 8780 68152 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 14246 8678 14298 8730
rect 14310 8678 14362 8730
rect 14374 8678 14426 8730
rect 14438 8678 14490 8730
rect 44246 8678 44298 8730
rect 44310 8678 44362 8730
rect 44374 8678 44426 8730
rect 44438 8678 44490 8730
rect 54246 8678 54298 8730
rect 54310 8678 54362 8730
rect 54374 8678 54426 8730
rect 54438 8678 54490 8730
rect 64246 8678 64298 8730
rect 64310 8678 64362 8730
rect 64374 8678 64426 8730
rect 64438 8678 64490 8730
rect 4620 8576 4672 8628
rect 6920 8619 6972 8628
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 9680 8576 9732 8628
rect 10784 8576 10836 8628
rect 17040 8576 17092 8628
rect 2688 8508 2740 8560
rect 16304 8508 16356 8560
rect 14464 8440 14516 8492
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 15292 8440 15344 8492
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 2596 8372 2648 8424
rect 12992 8372 13044 8424
rect 3056 8304 3108 8356
rect 3332 8304 3384 8356
rect 5724 8304 5776 8356
rect 6184 8304 6236 8356
rect 7564 8304 7616 8356
rect 8116 8347 8168 8356
rect 8116 8313 8125 8347
rect 8125 8313 8159 8347
rect 8159 8313 8168 8347
rect 8116 8304 8168 8313
rect 9036 8304 9088 8356
rect 9864 8304 9916 8356
rect 10784 8347 10836 8356
rect 10784 8313 10793 8347
rect 10793 8313 10827 8347
rect 10827 8313 10836 8347
rect 10784 8304 10836 8313
rect 15016 8372 15068 8424
rect 24492 8440 24544 8492
rect 31944 8440 31996 8492
rect 14832 8304 14884 8356
rect 18052 8372 18104 8424
rect 37096 8372 37148 8424
rect 38476 8372 38528 8424
rect 39396 8415 39448 8424
rect 17684 8304 17736 8356
rect 21088 8304 21140 8356
rect 32956 8304 33008 8356
rect 38660 8304 38712 8356
rect 39396 8381 39405 8415
rect 39405 8381 39439 8415
rect 39439 8381 39448 8415
rect 39396 8372 39448 8381
rect 40040 8415 40092 8424
rect 40040 8381 40049 8415
rect 40049 8381 40083 8415
rect 40083 8381 40092 8415
rect 40040 8372 40092 8381
rect 41052 8576 41104 8628
rect 48412 8576 48464 8628
rect 50620 8576 50672 8628
rect 50712 8576 50764 8628
rect 51448 8576 51500 8628
rect 51816 8576 51868 8628
rect 51908 8576 51960 8628
rect 54024 8576 54076 8628
rect 55036 8576 55088 8628
rect 61384 8619 61436 8628
rect 61384 8585 61393 8619
rect 61393 8585 61427 8619
rect 61427 8585 61436 8619
rect 61384 8576 61436 8585
rect 40500 8508 40552 8560
rect 43536 8508 43588 8560
rect 43720 8508 43772 8560
rect 43996 8508 44048 8560
rect 40316 8372 40368 8424
rect 41420 8415 41472 8424
rect 41420 8381 41429 8415
rect 41429 8381 41463 8415
rect 41463 8381 41472 8415
rect 41420 8372 41472 8381
rect 41328 8304 41380 8356
rect 42616 8372 42668 8424
rect 43536 8415 43588 8424
rect 43536 8381 43545 8415
rect 43545 8381 43579 8415
rect 43579 8381 43588 8415
rect 43536 8372 43588 8381
rect 45100 8372 45152 8424
rect 67088 8372 67140 8424
rect 67456 8415 67508 8424
rect 67456 8381 67465 8415
rect 67465 8381 67499 8415
rect 67499 8381 67508 8415
rect 67456 8372 67508 8381
rect 68100 8415 68152 8424
rect 68100 8381 68109 8415
rect 68109 8381 68143 8415
rect 68143 8381 68152 8415
rect 68100 8372 68152 8381
rect 45744 8347 45796 8356
rect 45744 8313 45753 8347
rect 45753 8313 45787 8347
rect 45787 8313 45796 8347
rect 45744 8304 45796 8313
rect 46664 8304 46716 8356
rect 47124 8304 47176 8356
rect 48136 8304 48188 8356
rect 48504 8304 48556 8356
rect 49056 8304 49108 8356
rect 52276 8304 52328 8356
rect 53380 8304 53432 8356
rect 54668 8347 54720 8356
rect 54668 8313 54677 8347
rect 54677 8313 54711 8347
rect 54711 8313 54720 8347
rect 54668 8304 54720 8313
rect 55220 8347 55272 8356
rect 55220 8313 55229 8347
rect 55229 8313 55263 8347
rect 55263 8313 55272 8347
rect 55220 8304 55272 8313
rect 55680 8347 55732 8356
rect 55680 8313 55689 8347
rect 55689 8313 55723 8347
rect 55723 8313 55732 8347
rect 55680 8304 55732 8313
rect 62212 8347 62264 8356
rect 62212 8313 62221 8347
rect 62221 8313 62255 8347
rect 62255 8313 62264 8347
rect 62212 8304 62264 8313
rect 62580 8304 62632 8356
rect 64604 8304 64656 8356
rect 65616 8347 65668 8356
rect 65616 8313 65625 8347
rect 65625 8313 65659 8347
rect 65659 8313 65668 8347
rect 65616 8304 65668 8313
rect 66444 8304 66496 8356
rect 68192 8304 68244 8356
rect 2872 8236 2924 8288
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 12256 8236 12308 8288
rect 15200 8236 15252 8288
rect 15384 8236 15436 8288
rect 41420 8236 41472 8288
rect 41696 8236 41748 8288
rect 43996 8279 44048 8288
rect 43996 8245 44005 8279
rect 44005 8245 44039 8279
rect 44039 8245 44048 8279
rect 43996 8236 44048 8245
rect 45376 8236 45428 8288
rect 46204 8279 46256 8288
rect 46204 8245 46213 8279
rect 46213 8245 46247 8279
rect 46247 8245 46256 8279
rect 46204 8236 46256 8245
rect 57336 8236 57388 8288
rect 57520 8236 57572 8288
rect 64696 8236 64748 8288
rect 9246 8134 9298 8186
rect 9310 8134 9362 8186
rect 9374 8134 9426 8186
rect 9438 8134 9490 8186
rect 39246 8134 39298 8186
rect 39310 8134 39362 8186
rect 39374 8134 39426 8186
rect 39438 8134 39490 8186
rect 49246 8134 49298 8186
rect 49310 8134 49362 8186
rect 49374 8134 49426 8186
rect 49438 8134 49490 8186
rect 59246 8134 59298 8186
rect 59310 8134 59362 8186
rect 59374 8134 59426 8186
rect 59438 8134 59490 8186
rect 6276 8075 6328 8084
rect 6276 8041 6285 8075
rect 6285 8041 6319 8075
rect 6319 8041 6328 8075
rect 6276 8032 6328 8041
rect 14556 8032 14608 8084
rect 15016 8032 15068 8084
rect 11244 7896 11296 7948
rect 11704 7896 11756 7948
rect 12624 7896 12676 7948
rect 13912 7896 13964 7948
rect 17040 8032 17092 8084
rect 17224 8032 17276 8084
rect 36912 8032 36964 8084
rect 16488 7964 16540 8016
rect 23296 7964 23348 8016
rect 34980 7964 35032 8016
rect 38660 7964 38712 8016
rect 17132 7939 17184 7948
rect 12716 7828 12768 7880
rect 17132 7905 17141 7939
rect 17141 7905 17175 7939
rect 17175 7905 17184 7939
rect 17132 7896 17184 7905
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 23756 7896 23808 7948
rect 32036 7896 32088 7948
rect 37924 7896 37976 7948
rect 39028 7964 39080 8016
rect 40316 8032 40368 8084
rect 42984 8032 43036 8084
rect 55404 8032 55456 8084
rect 56048 8032 56100 8084
rect 57244 8032 57296 8084
rect 57428 8032 57480 8084
rect 16948 7828 17000 7880
rect 20996 7828 21048 7880
rect 39672 7896 39724 7948
rect 41420 7896 41472 7948
rect 41880 7896 41932 7948
rect 42800 7896 42852 7948
rect 42984 7896 43036 7948
rect 46204 7964 46256 8016
rect 43904 7896 43956 7948
rect 44088 7896 44140 7948
rect 44916 7896 44968 7948
rect 46940 7896 46992 7948
rect 55956 7896 56008 7948
rect 67180 7896 67232 7948
rect 67640 7896 67692 7948
rect 68008 7939 68060 7948
rect 68008 7905 68017 7939
rect 68017 7905 68051 7939
rect 68051 7905 68060 7939
rect 68008 7896 68060 7905
rect 43628 7828 43680 7880
rect 45560 7828 45612 7880
rect 48412 7828 48464 7880
rect 66628 7828 66680 7880
rect 68284 7828 68336 7880
rect 15200 7760 15252 7812
rect 15292 7760 15344 7812
rect 23664 7760 23716 7812
rect 38660 7760 38712 7812
rect 41880 7760 41932 7812
rect 48596 7760 48648 7812
rect 65340 7760 65392 7812
rect 66168 7760 66220 7812
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 4804 7692 4856 7744
rect 4896 7692 4948 7744
rect 5540 7692 5592 7744
rect 7380 7692 7432 7744
rect 7932 7692 7984 7744
rect 8392 7692 8444 7744
rect 8944 7692 8996 7744
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 11520 7692 11572 7744
rect 16488 7692 16540 7744
rect 39672 7692 39724 7744
rect 44732 7692 44784 7744
rect 45560 7692 45612 7744
rect 46204 7735 46256 7744
rect 46204 7701 46213 7735
rect 46213 7701 46247 7735
rect 46247 7701 46256 7735
rect 46204 7692 46256 7701
rect 46848 7735 46900 7744
rect 46848 7701 46857 7735
rect 46857 7701 46891 7735
rect 46891 7701 46900 7735
rect 46848 7692 46900 7701
rect 47216 7692 47268 7744
rect 47860 7735 47912 7744
rect 47860 7701 47869 7735
rect 47869 7701 47903 7735
rect 47903 7701 47912 7735
rect 47860 7692 47912 7701
rect 48320 7692 48372 7744
rect 50344 7692 50396 7744
rect 50896 7735 50948 7744
rect 50896 7701 50905 7735
rect 50905 7701 50939 7735
rect 50939 7701 50948 7735
rect 50896 7692 50948 7701
rect 51448 7735 51500 7744
rect 51448 7701 51457 7735
rect 51457 7701 51491 7735
rect 51491 7701 51500 7735
rect 51448 7692 51500 7701
rect 52092 7735 52144 7744
rect 52092 7701 52101 7735
rect 52101 7701 52135 7735
rect 52135 7701 52144 7735
rect 52092 7692 52144 7701
rect 52368 7692 52420 7744
rect 52828 7692 52880 7744
rect 53472 7692 53524 7744
rect 53748 7692 53800 7744
rect 54852 7692 54904 7744
rect 55956 7692 56008 7744
rect 60832 7735 60884 7744
rect 60832 7701 60841 7735
rect 60841 7701 60875 7735
rect 60875 7701 60884 7735
rect 60832 7692 60884 7701
rect 61936 7735 61988 7744
rect 61936 7701 61945 7735
rect 61945 7701 61979 7735
rect 61979 7701 61988 7735
rect 61936 7692 61988 7701
rect 62488 7735 62540 7744
rect 62488 7701 62497 7735
rect 62497 7701 62531 7735
rect 62531 7701 62540 7735
rect 62488 7692 62540 7701
rect 63040 7735 63092 7744
rect 63040 7701 63049 7735
rect 63049 7701 63083 7735
rect 63083 7701 63092 7735
rect 63040 7692 63092 7701
rect 63868 7692 63920 7744
rect 65156 7692 65208 7744
rect 65892 7735 65944 7744
rect 65892 7701 65901 7735
rect 65901 7701 65935 7735
rect 65935 7701 65944 7735
rect 65892 7692 65944 7701
rect 66628 7735 66680 7744
rect 66628 7701 66637 7735
rect 66637 7701 66671 7735
rect 66671 7701 66680 7735
rect 66628 7692 66680 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 14246 7590 14298 7642
rect 14310 7590 14362 7642
rect 14374 7590 14426 7642
rect 14438 7590 14490 7642
rect 44246 7590 44298 7642
rect 44310 7590 44362 7642
rect 44374 7590 44426 7642
rect 44438 7590 44490 7642
rect 54246 7590 54298 7642
rect 54310 7590 54362 7642
rect 54374 7590 54426 7642
rect 54438 7590 54490 7642
rect 64246 7590 64298 7642
rect 64310 7590 64362 7642
rect 64374 7590 64426 7642
rect 64438 7590 64490 7642
rect 4068 7488 4120 7540
rect 6828 7488 6880 7540
rect 7012 7488 7064 7540
rect 35256 7488 35308 7540
rect 39672 7488 39724 7540
rect 56784 7531 56836 7540
rect 56784 7497 56793 7531
rect 56793 7497 56827 7531
rect 56827 7497 56836 7531
rect 56784 7488 56836 7497
rect 57152 7488 57204 7540
rect 57520 7488 57572 7540
rect 57980 7531 58032 7540
rect 57980 7497 57989 7531
rect 57989 7497 58023 7531
rect 58023 7497 58032 7531
rect 57980 7488 58032 7497
rect 60188 7531 60240 7540
rect 60188 7497 60197 7531
rect 60197 7497 60231 7531
rect 60231 7497 60240 7531
rect 60188 7488 60240 7497
rect 60740 7531 60792 7540
rect 60740 7497 60749 7531
rect 60749 7497 60783 7531
rect 60783 7497 60792 7531
rect 60740 7488 60792 7497
rect 61108 7488 61160 7540
rect 61660 7531 61712 7540
rect 61660 7497 61669 7531
rect 61669 7497 61703 7531
rect 61703 7497 61712 7531
rect 61660 7488 61712 7497
rect 61844 7488 61896 7540
rect 4620 7352 4672 7404
rect 1860 7284 1912 7336
rect 2504 7284 2556 7336
rect 6920 7284 6972 7336
rect 7472 7284 7524 7336
rect 10416 7284 10468 7336
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11336 7284 11388 7336
rect 12900 7284 12952 7336
rect 13268 7284 13320 7336
rect 17684 7420 17736 7472
rect 35624 7420 35676 7472
rect 40316 7420 40368 7472
rect 61200 7420 61252 7472
rect 15292 7284 15344 7336
rect 15384 7284 15436 7336
rect 16672 7352 16724 7404
rect 19524 7352 19576 7404
rect 36268 7352 36320 7404
rect 6276 7216 6328 7268
rect 11428 7216 11480 7268
rect 2228 7148 2280 7200
rect 4068 7148 4120 7200
rect 5448 7148 5500 7200
rect 5724 7148 5776 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 11888 7148 11940 7200
rect 18236 7327 18288 7336
rect 18236 7293 18245 7327
rect 18245 7293 18279 7327
rect 18279 7293 18288 7327
rect 18236 7284 18288 7293
rect 38108 7327 38160 7336
rect 38108 7293 38117 7327
rect 38117 7293 38151 7327
rect 38151 7293 38160 7327
rect 38108 7284 38160 7293
rect 38752 7327 38804 7336
rect 17776 7216 17828 7268
rect 21732 7216 21784 7268
rect 33048 7216 33100 7268
rect 38752 7293 38761 7327
rect 38761 7293 38795 7327
rect 38795 7293 38804 7327
rect 38752 7284 38804 7293
rect 40132 7352 40184 7404
rect 39120 7216 39172 7268
rect 40316 7284 40368 7336
rect 40776 7327 40828 7336
rect 40776 7293 40785 7327
rect 40785 7293 40819 7327
rect 40819 7293 40828 7327
rect 40776 7284 40828 7293
rect 44088 7352 44140 7404
rect 41512 7284 41564 7336
rect 41696 7284 41748 7336
rect 43076 7284 43128 7336
rect 43352 7327 43404 7336
rect 43352 7293 43361 7327
rect 43361 7293 43395 7327
rect 43395 7293 43404 7327
rect 43352 7284 43404 7293
rect 44732 7284 44784 7336
rect 46388 7352 46440 7404
rect 65248 7352 65300 7404
rect 40132 7216 40184 7268
rect 44364 7216 44416 7268
rect 47584 7284 47636 7336
rect 50160 7284 50212 7336
rect 69296 7352 69348 7404
rect 65984 7284 66036 7336
rect 66260 7284 66312 7336
rect 66720 7327 66772 7336
rect 66720 7293 66729 7327
rect 66729 7293 66763 7327
rect 66763 7293 66772 7327
rect 66720 7284 66772 7293
rect 46112 7216 46164 7268
rect 49976 7216 50028 7268
rect 51724 7216 51776 7268
rect 53840 7216 53892 7268
rect 66996 7216 67048 7268
rect 67824 7284 67876 7336
rect 68100 7259 68152 7268
rect 68100 7225 68109 7259
rect 68109 7225 68143 7259
rect 68143 7225 68152 7259
rect 68100 7216 68152 7225
rect 19432 7148 19484 7200
rect 32496 7148 32548 7200
rect 38752 7148 38804 7200
rect 40776 7148 40828 7200
rect 41236 7148 41288 7200
rect 45928 7191 45980 7200
rect 45928 7157 45937 7191
rect 45937 7157 45971 7191
rect 45971 7157 45980 7191
rect 45928 7148 45980 7157
rect 46388 7148 46440 7200
rect 47400 7148 47452 7200
rect 48228 7191 48280 7200
rect 48228 7157 48237 7191
rect 48237 7157 48271 7191
rect 48271 7157 48280 7191
rect 48228 7148 48280 7157
rect 48964 7148 49016 7200
rect 49148 7148 49200 7200
rect 49884 7191 49936 7200
rect 49884 7157 49893 7191
rect 49893 7157 49927 7191
rect 49927 7157 49936 7191
rect 49884 7148 49936 7157
rect 50804 7148 50856 7200
rect 52184 7191 52236 7200
rect 52184 7157 52193 7191
rect 52193 7157 52227 7191
rect 52227 7157 52236 7191
rect 52184 7148 52236 7157
rect 52920 7148 52972 7200
rect 53748 7148 53800 7200
rect 55036 7148 55088 7200
rect 55496 7148 55548 7200
rect 56232 7191 56284 7200
rect 56232 7157 56241 7191
rect 56241 7157 56275 7191
rect 56275 7157 56284 7191
rect 56232 7148 56284 7157
rect 59544 7148 59596 7200
rect 62396 7148 62448 7200
rect 62764 7191 62816 7200
rect 62764 7157 62773 7191
rect 62773 7157 62807 7191
rect 62807 7157 62816 7191
rect 62764 7148 62816 7157
rect 63316 7191 63368 7200
rect 63316 7157 63325 7191
rect 63325 7157 63359 7191
rect 63359 7157 63368 7191
rect 63316 7148 63368 7157
rect 63500 7148 63552 7200
rect 64788 7191 64840 7200
rect 64788 7157 64797 7191
rect 64797 7157 64831 7191
rect 64831 7157 64840 7191
rect 64788 7148 64840 7157
rect 66720 7148 66772 7200
rect 9246 7046 9298 7098
rect 9310 7046 9362 7098
rect 9374 7046 9426 7098
rect 9438 7046 9490 7098
rect 39246 7046 39298 7098
rect 39310 7046 39362 7098
rect 39374 7046 39426 7098
rect 39438 7046 39490 7098
rect 49246 7046 49298 7098
rect 49310 7046 49362 7098
rect 49374 7046 49426 7098
rect 49438 7046 49490 7098
rect 59246 7046 59298 7098
rect 59310 7046 59362 7098
rect 59374 7046 59426 7098
rect 59438 7046 59490 7098
rect 12164 6944 12216 6996
rect 13084 6944 13136 6996
rect 31760 6944 31812 6996
rect 40316 6944 40368 6996
rect 41420 6944 41472 6996
rect 44364 6944 44416 6996
rect 62488 6944 62540 6996
rect 67824 6944 67876 6996
rect 38476 6876 38528 6928
rect 40132 6876 40184 6928
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 10232 6851 10284 6860
rect 10232 6817 10241 6851
rect 10241 6817 10275 6851
rect 10275 6817 10284 6851
rect 10232 6808 10284 6817
rect 11612 6808 11664 6860
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 12440 6808 12492 6817
rect 11980 6740 12032 6792
rect 12532 6740 12584 6792
rect 13728 6808 13780 6860
rect 15384 6851 15436 6860
rect 2504 6672 2556 6724
rect 6000 6672 6052 6724
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 15844 6808 15896 6860
rect 16120 6808 16172 6860
rect 16580 6808 16632 6860
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 18144 6808 18196 6860
rect 19064 6808 19116 6860
rect 38568 6851 38620 6860
rect 22652 6740 22704 6792
rect 38568 6817 38577 6851
rect 38577 6817 38611 6851
rect 38611 6817 38620 6851
rect 38568 6808 38620 6817
rect 38752 6808 38804 6860
rect 39856 6740 39908 6792
rect 2596 6647 2648 6656
rect 2596 6613 2605 6647
rect 2605 6613 2639 6647
rect 2639 6613 2648 6647
rect 2596 6604 2648 6613
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 3792 6604 3844 6656
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 6092 6604 6144 6656
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 7656 6604 7708 6656
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 13728 6604 13780 6656
rect 17040 6604 17092 6656
rect 17592 6672 17644 6724
rect 20904 6672 20956 6724
rect 37004 6672 37056 6724
rect 41144 6808 41196 6860
rect 41420 6808 41472 6860
rect 42156 6851 42208 6860
rect 42156 6817 42165 6851
rect 42165 6817 42199 6851
rect 42199 6817 42208 6851
rect 42156 6808 42208 6817
rect 43168 6876 43220 6928
rect 42892 6808 42944 6860
rect 40132 6740 40184 6792
rect 44732 6808 44784 6860
rect 44548 6740 44600 6792
rect 45192 6808 45244 6860
rect 18972 6604 19024 6656
rect 37832 6604 37884 6656
rect 45192 6672 45244 6724
rect 45560 6876 45612 6928
rect 45836 6808 45888 6860
rect 47492 6851 47544 6860
rect 45560 6740 45612 6792
rect 46572 6740 46624 6792
rect 47492 6817 47501 6851
rect 47501 6817 47535 6851
rect 47535 6817 47544 6851
rect 47492 6808 47544 6817
rect 59636 6808 59688 6860
rect 65340 6876 65392 6928
rect 65432 6808 65484 6860
rect 47124 6740 47176 6792
rect 47308 6740 47360 6792
rect 64144 6740 64196 6792
rect 65340 6740 65392 6792
rect 67272 6808 67324 6860
rect 67732 6808 67784 6860
rect 68468 6740 68520 6792
rect 46112 6672 46164 6724
rect 48044 6672 48096 6724
rect 57612 6672 57664 6724
rect 64052 6672 64104 6724
rect 65800 6672 65852 6724
rect 40316 6604 40368 6656
rect 46388 6604 46440 6656
rect 46572 6604 46624 6656
rect 47124 6604 47176 6656
rect 49792 6604 49844 6656
rect 50068 6604 50120 6656
rect 50712 6604 50764 6656
rect 51264 6604 51316 6656
rect 51816 6604 51868 6656
rect 52552 6647 52604 6656
rect 52552 6613 52561 6647
rect 52561 6613 52595 6647
rect 52595 6613 52604 6647
rect 52552 6604 52604 6613
rect 53196 6647 53248 6656
rect 53196 6613 53205 6647
rect 53205 6613 53239 6647
rect 53239 6613 53248 6647
rect 53196 6604 53248 6613
rect 53932 6647 53984 6656
rect 53932 6613 53941 6647
rect 53941 6613 53975 6647
rect 53975 6613 53984 6647
rect 53932 6604 53984 6613
rect 54576 6647 54628 6656
rect 54576 6613 54585 6647
rect 54585 6613 54619 6647
rect 54619 6613 54628 6647
rect 54576 6604 54628 6613
rect 54944 6604 54996 6656
rect 55404 6604 55456 6656
rect 56324 6604 56376 6656
rect 57244 6647 57296 6656
rect 57244 6613 57253 6647
rect 57253 6613 57287 6647
rect 57287 6613 57296 6647
rect 57244 6604 57296 6613
rect 57888 6647 57940 6656
rect 57888 6613 57897 6647
rect 57897 6613 57931 6647
rect 57931 6613 57940 6647
rect 57888 6604 57940 6613
rect 60188 6604 60240 6656
rect 60372 6647 60424 6656
rect 60372 6613 60381 6647
rect 60381 6613 60415 6647
rect 60415 6613 60424 6647
rect 60372 6604 60424 6613
rect 61384 6647 61436 6656
rect 61384 6613 61393 6647
rect 61393 6613 61427 6647
rect 61427 6613 61436 6647
rect 61384 6604 61436 6613
rect 62028 6647 62080 6656
rect 62028 6613 62037 6647
rect 62037 6613 62071 6647
rect 62071 6613 62080 6647
rect 62028 6604 62080 6613
rect 62856 6647 62908 6656
rect 62856 6613 62865 6647
rect 62865 6613 62899 6647
rect 62899 6613 62908 6647
rect 62856 6604 62908 6613
rect 63408 6647 63460 6656
rect 63408 6613 63417 6647
rect 63417 6613 63451 6647
rect 63451 6613 63460 6647
rect 63408 6604 63460 6613
rect 64144 6647 64196 6656
rect 64144 6613 64153 6647
rect 64153 6613 64187 6647
rect 64187 6613 64196 6647
rect 64144 6604 64196 6613
rect 67548 6604 67600 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 14246 6502 14298 6554
rect 14310 6502 14362 6554
rect 14374 6502 14426 6554
rect 14438 6502 14490 6554
rect 44246 6502 44298 6554
rect 44310 6502 44362 6554
rect 44374 6502 44426 6554
rect 44438 6502 44490 6554
rect 54246 6502 54298 6554
rect 54310 6502 54362 6554
rect 54374 6502 54426 6554
rect 54438 6502 54490 6554
rect 64246 6502 64298 6554
rect 64310 6502 64362 6554
rect 64374 6502 64426 6554
rect 64438 6502 64490 6554
rect 15384 6400 15436 6452
rect 16304 6400 16356 6452
rect 20444 6400 20496 6452
rect 39764 6400 39816 6452
rect 39856 6400 39908 6452
rect 5080 6264 5132 6316
rect 7012 6264 7064 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 1676 6196 1728 6248
rect 2964 6196 3016 6248
rect 9128 6196 9180 6248
rect 9588 6196 9640 6248
rect 9772 6196 9824 6248
rect 11060 6196 11112 6248
rect 13176 6239 13228 6248
rect 5080 6128 5132 6180
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 14464 6239 14516 6248
rect 13636 6128 13688 6180
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 16120 6264 16172 6316
rect 15568 6196 15620 6248
rect 16212 6196 16264 6248
rect 16304 6196 16356 6248
rect 22560 6332 22612 6384
rect 36544 6332 36596 6384
rect 45652 6400 45704 6452
rect 16856 6264 16908 6316
rect 19156 6264 19208 6316
rect 35532 6264 35584 6316
rect 37924 6307 37976 6316
rect 19340 6196 19392 6248
rect 19892 6196 19944 6248
rect 37924 6273 37933 6307
rect 37933 6273 37967 6307
rect 37967 6273 37976 6307
rect 37924 6264 37976 6273
rect 39856 6264 39908 6316
rect 42800 6332 42852 6384
rect 44180 6264 44232 6316
rect 47216 6332 47268 6384
rect 14096 6128 14148 6180
rect 23388 6128 23440 6180
rect 35348 6128 35400 6180
rect 40868 6196 40920 6248
rect 41604 6196 41656 6248
rect 42064 6239 42116 6248
rect 42064 6205 42073 6239
rect 42073 6205 42107 6239
rect 42107 6205 42116 6239
rect 42064 6196 42116 6205
rect 43076 6196 43128 6248
rect 43444 6196 43496 6248
rect 3608 6103 3660 6112
rect 3608 6069 3617 6103
rect 3617 6069 3651 6103
rect 3651 6069 3660 6103
rect 3608 6060 3660 6069
rect 4620 6060 4672 6112
rect 4988 6060 5040 6112
rect 5724 6060 5776 6112
rect 6736 6103 6788 6112
rect 6736 6069 6745 6103
rect 6745 6069 6779 6103
rect 6779 6069 6788 6103
rect 6736 6060 6788 6069
rect 10876 6060 10928 6112
rect 16580 6060 16632 6112
rect 35440 6060 35492 6112
rect 42984 6128 43036 6180
rect 43812 6128 43864 6180
rect 44732 6196 44784 6248
rect 45652 6196 45704 6248
rect 47032 6196 47084 6248
rect 49976 6196 50028 6248
rect 50896 6239 50948 6248
rect 50896 6205 50905 6239
rect 50905 6205 50939 6239
rect 50939 6205 50948 6239
rect 50896 6196 50948 6205
rect 55864 6196 55916 6248
rect 64696 6196 64748 6248
rect 65064 6196 65116 6248
rect 66444 6196 66496 6248
rect 66904 6196 66956 6248
rect 67088 6239 67140 6248
rect 67088 6205 67097 6239
rect 67097 6205 67131 6239
rect 67131 6205 67140 6239
rect 67088 6196 67140 6205
rect 67548 6196 67600 6248
rect 41144 6060 41196 6112
rect 47860 6128 47912 6180
rect 47952 6128 48004 6180
rect 56416 6128 56468 6180
rect 59912 6128 59964 6180
rect 46940 6060 46992 6112
rect 52644 6060 52696 6112
rect 53288 6060 53340 6112
rect 54760 6060 54812 6112
rect 55128 6060 55180 6112
rect 55588 6103 55640 6112
rect 55588 6069 55597 6103
rect 55597 6069 55631 6103
rect 55631 6069 55640 6103
rect 55588 6060 55640 6069
rect 56140 6103 56192 6112
rect 56140 6069 56149 6103
rect 56149 6069 56183 6103
rect 56183 6069 56192 6103
rect 56140 6060 56192 6069
rect 56876 6060 56928 6112
rect 57520 6103 57572 6112
rect 57520 6069 57529 6103
rect 57529 6069 57563 6103
rect 57563 6069 57572 6103
rect 57520 6060 57572 6069
rect 58900 6103 58952 6112
rect 58900 6069 58909 6103
rect 58909 6069 58943 6103
rect 58943 6069 58952 6103
rect 58900 6060 58952 6069
rect 59820 6060 59872 6112
rect 60096 6103 60148 6112
rect 60096 6069 60105 6103
rect 60105 6069 60139 6103
rect 60139 6069 60148 6103
rect 60096 6060 60148 6069
rect 61660 6103 61712 6112
rect 61660 6069 61669 6103
rect 61669 6069 61703 6103
rect 61703 6069 61712 6103
rect 61660 6060 61712 6069
rect 62304 6103 62356 6112
rect 62304 6069 62313 6103
rect 62313 6069 62347 6103
rect 62347 6069 62356 6103
rect 62304 6060 62356 6069
rect 63224 6060 63276 6112
rect 63684 6060 63736 6112
rect 64512 6060 64564 6112
rect 9246 5958 9298 6010
rect 9310 5958 9362 6010
rect 9374 5958 9426 6010
rect 9438 5958 9490 6010
rect 39246 5958 39298 6010
rect 39310 5958 39362 6010
rect 39374 5958 39426 6010
rect 39438 5958 39490 6010
rect 49246 5958 49298 6010
rect 49310 5958 49362 6010
rect 49374 5958 49426 6010
rect 49438 5958 49490 6010
rect 59246 5958 59298 6010
rect 59310 5958 59362 6010
rect 59374 5958 59426 6010
rect 59438 5958 59490 6010
rect 10048 5856 10100 5908
rect 1768 5831 1820 5840
rect 1768 5797 1777 5831
rect 1777 5797 1811 5831
rect 1811 5797 1820 5831
rect 1768 5788 1820 5797
rect 2780 5788 2832 5840
rect 2044 5720 2096 5772
rect 2688 5763 2740 5772
rect 2688 5729 2697 5763
rect 2697 5729 2731 5763
rect 2731 5729 2740 5763
rect 2688 5720 2740 5729
rect 3332 5763 3384 5772
rect 3332 5729 3341 5763
rect 3341 5729 3375 5763
rect 3375 5729 3384 5763
rect 3332 5720 3384 5729
rect 4896 5720 4948 5772
rect 5540 5720 5592 5772
rect 8300 5720 8352 5772
rect 3056 5652 3108 5704
rect 10324 5720 10376 5772
rect 10692 5720 10744 5772
rect 12072 5720 12124 5772
rect 13360 5856 13412 5908
rect 20352 5856 20404 5908
rect 35992 5856 36044 5908
rect 42064 5856 42116 5908
rect 42708 5856 42760 5908
rect 13728 5720 13780 5772
rect 15292 5788 15344 5840
rect 38384 5788 38436 5840
rect 43812 5788 43864 5840
rect 44088 5788 44140 5840
rect 44456 5856 44508 5908
rect 46112 5856 46164 5908
rect 15384 5763 15436 5772
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 2320 5516 2372 5568
rect 6276 5559 6328 5568
rect 6276 5525 6285 5559
rect 6285 5525 6319 5559
rect 6319 5525 6328 5559
rect 6276 5516 6328 5525
rect 7748 5516 7800 5568
rect 9404 5516 9456 5568
rect 9956 5584 10008 5636
rect 15476 5652 15528 5704
rect 16488 5720 16540 5772
rect 16580 5652 16632 5704
rect 17040 5720 17092 5772
rect 20076 5720 20128 5772
rect 33968 5720 34020 5772
rect 40316 5720 40368 5772
rect 41328 5720 41380 5772
rect 41788 5720 41840 5772
rect 42340 5763 42392 5772
rect 42340 5729 42349 5763
rect 42349 5729 42383 5763
rect 42383 5729 42392 5763
rect 42340 5720 42392 5729
rect 42800 5763 42852 5772
rect 42800 5729 42809 5763
rect 42809 5729 42843 5763
rect 42843 5729 42852 5763
rect 42800 5720 42852 5729
rect 19340 5652 19392 5704
rect 37924 5652 37976 5704
rect 43996 5720 44048 5772
rect 46940 5788 46992 5840
rect 14464 5584 14516 5636
rect 19616 5584 19668 5636
rect 31944 5627 31996 5636
rect 31944 5593 31953 5627
rect 31953 5593 31987 5627
rect 31987 5593 31996 5627
rect 31944 5584 31996 5593
rect 36820 5584 36872 5636
rect 39212 5627 39264 5636
rect 39212 5593 39221 5627
rect 39221 5593 39255 5627
rect 39255 5593 39264 5627
rect 39212 5584 39264 5593
rect 40316 5584 40368 5636
rect 40776 5584 40828 5636
rect 18144 5516 18196 5568
rect 24492 5559 24544 5568
rect 24492 5525 24501 5559
rect 24501 5525 24535 5559
rect 24535 5525 24544 5559
rect 24492 5516 24544 5525
rect 24952 5516 25004 5568
rect 31760 5559 31812 5568
rect 31760 5525 31769 5559
rect 31769 5525 31803 5559
rect 31803 5525 31812 5559
rect 32036 5559 32088 5568
rect 31760 5516 31812 5525
rect 32036 5525 32045 5559
rect 32045 5525 32079 5559
rect 32079 5525 32088 5559
rect 32036 5516 32088 5525
rect 32312 5559 32364 5568
rect 32312 5525 32321 5559
rect 32321 5525 32355 5559
rect 32355 5525 32364 5559
rect 32312 5516 32364 5525
rect 32496 5559 32548 5568
rect 32496 5525 32505 5559
rect 32505 5525 32539 5559
rect 32539 5525 32548 5559
rect 32496 5516 32548 5525
rect 37740 5516 37792 5568
rect 38568 5516 38620 5568
rect 39856 5516 39908 5568
rect 42156 5584 42208 5636
rect 42800 5584 42852 5636
rect 45376 5720 45428 5772
rect 46664 5720 46716 5772
rect 47676 5856 47728 5908
rect 47860 5856 47912 5908
rect 66536 5788 66588 5840
rect 67824 5788 67876 5840
rect 48136 5720 48188 5772
rect 48504 5720 48556 5772
rect 49056 5720 49108 5772
rect 50160 5720 50212 5772
rect 51172 5720 51224 5772
rect 51724 5720 51776 5772
rect 52368 5720 52420 5772
rect 52828 5720 52880 5772
rect 52920 5652 52972 5704
rect 53104 5652 53156 5704
rect 55036 5720 55088 5772
rect 55496 5720 55548 5772
rect 56416 5720 56468 5772
rect 62580 5720 62632 5772
rect 63500 5763 63552 5772
rect 63500 5729 63509 5763
rect 63509 5729 63543 5763
rect 63543 5729 63552 5763
rect 63500 5720 63552 5729
rect 64052 5720 64104 5772
rect 64604 5720 64656 5772
rect 54944 5652 54996 5704
rect 66168 5720 66220 5772
rect 68100 5763 68152 5772
rect 68100 5729 68109 5763
rect 68109 5729 68143 5763
rect 68143 5729 68152 5763
rect 68100 5720 68152 5729
rect 65616 5652 65668 5704
rect 69020 5652 69072 5704
rect 44456 5584 44508 5636
rect 45376 5584 45428 5636
rect 51724 5584 51776 5636
rect 52000 5584 52052 5636
rect 52368 5584 52420 5636
rect 60556 5584 60608 5636
rect 64512 5584 64564 5636
rect 69848 5584 69900 5636
rect 41696 5516 41748 5568
rect 44548 5516 44600 5568
rect 56784 5516 56836 5568
rect 57704 5559 57756 5568
rect 57704 5525 57713 5559
rect 57713 5525 57747 5559
rect 57747 5525 57756 5559
rect 57704 5516 57756 5525
rect 58808 5559 58860 5568
rect 58808 5525 58817 5559
rect 58817 5525 58851 5559
rect 58851 5525 58860 5559
rect 58808 5516 58860 5525
rect 60004 5516 60056 5568
rect 60280 5559 60332 5568
rect 60280 5525 60289 5559
rect 60289 5525 60323 5559
rect 60323 5525 60332 5559
rect 60280 5516 60332 5525
rect 60464 5516 60516 5568
rect 61752 5516 61804 5568
rect 64696 5516 64748 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 14246 5414 14298 5466
rect 14310 5414 14362 5466
rect 14374 5414 14426 5466
rect 14438 5414 14490 5466
rect 12164 5312 12216 5364
rect 37280 5448 37332 5500
rect 44246 5414 44298 5466
rect 44310 5414 44362 5466
rect 44374 5414 44426 5466
rect 44438 5414 44490 5466
rect 54246 5414 54298 5466
rect 54310 5414 54362 5466
rect 54374 5414 54426 5466
rect 54438 5414 54490 5466
rect 64246 5414 64298 5466
rect 64310 5414 64362 5466
rect 64374 5414 64426 5466
rect 64438 5414 64490 5466
rect 36176 5312 36228 5364
rect 40224 5312 40276 5364
rect 46204 5312 46256 5364
rect 4804 5244 4856 5296
rect 1492 5108 1544 5160
rect 1584 5108 1636 5160
rect 1952 5108 2004 5160
rect 2780 5108 2832 5160
rect 4068 5176 4120 5228
rect 3332 5108 3384 5160
rect 3884 5108 3936 5160
rect 4160 5151 4212 5160
rect 4160 5117 4169 5151
rect 4169 5117 4203 5151
rect 4203 5117 4212 5151
rect 4160 5108 4212 5117
rect 4804 5151 4856 5160
rect 4804 5117 4813 5151
rect 4813 5117 4847 5151
rect 4847 5117 4856 5151
rect 5448 5244 5500 5296
rect 9036 5244 9088 5296
rect 9404 5244 9456 5296
rect 5448 5151 5500 5160
rect 4804 5108 4856 5117
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 6092 5108 6144 5160
rect 6644 5108 6696 5160
rect 7288 5108 7340 5160
rect 7564 5151 7616 5160
rect 7564 5117 7573 5151
rect 7573 5117 7607 5151
rect 7607 5117 7616 5151
rect 7564 5108 7616 5117
rect 7472 5040 7524 5092
rect 8116 5108 8168 5160
rect 8852 5108 8904 5160
rect 9680 5108 9732 5160
rect 9864 5108 9916 5160
rect 20720 5244 20772 5296
rect 23572 5244 23624 5296
rect 42340 5244 42392 5296
rect 42616 5244 42668 5296
rect 44180 5244 44232 5296
rect 13360 5151 13412 5160
rect 7748 5040 7800 5092
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 13544 5108 13596 5160
rect 14556 5176 14608 5228
rect 14924 5176 14976 5228
rect 9864 4972 9916 5024
rect 10968 4972 11020 5024
rect 15568 5108 15620 5160
rect 21824 5176 21876 5228
rect 33048 5176 33100 5228
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 37740 5108 37792 5160
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 14464 5040 14516 5049
rect 14648 5083 14700 5092
rect 14648 5049 14657 5083
rect 14657 5049 14691 5083
rect 14691 5049 14700 5083
rect 14648 5040 14700 5049
rect 17684 5083 17736 5092
rect 17684 5049 17693 5083
rect 17693 5049 17727 5083
rect 17727 5049 17736 5083
rect 17684 5040 17736 5049
rect 38384 5040 38436 5092
rect 38844 5108 38896 5160
rect 39764 5108 39816 5160
rect 41972 5108 42024 5160
rect 44548 5176 44600 5228
rect 43352 5108 43404 5160
rect 17500 4972 17552 5024
rect 37188 4972 37240 5024
rect 40224 5040 40276 5092
rect 42524 5040 42576 5092
rect 42616 5040 42668 5092
rect 44456 5108 44508 5160
rect 45100 5244 45152 5296
rect 45652 5108 45704 5160
rect 45836 5108 45888 5160
rect 47952 5176 48004 5228
rect 46756 5151 46808 5160
rect 46756 5117 46765 5151
rect 46765 5117 46799 5151
rect 46799 5117 46808 5151
rect 46756 5108 46808 5117
rect 47308 5108 47360 5160
rect 46388 5040 46440 5092
rect 48320 5312 48372 5364
rect 50528 5244 50580 5296
rect 63592 5244 63644 5296
rect 64236 5244 64288 5296
rect 48320 5176 48372 5228
rect 51080 5176 51132 5228
rect 60832 5176 60884 5228
rect 48596 5108 48648 5160
rect 50344 5108 50396 5160
rect 50528 5108 50580 5160
rect 50620 5108 50672 5160
rect 51356 5083 51408 5092
rect 51356 5049 51365 5083
rect 51365 5049 51399 5083
rect 51399 5049 51408 5083
rect 51356 5040 51408 5049
rect 48136 4972 48188 5024
rect 51908 5108 51960 5160
rect 52092 5108 52144 5160
rect 53748 5108 53800 5160
rect 53840 5040 53892 5092
rect 54944 5108 54996 5160
rect 55404 5108 55456 5160
rect 55956 5151 56008 5160
rect 55956 5117 55965 5151
rect 55965 5117 55999 5151
rect 55999 5117 56008 5151
rect 55956 5108 56008 5117
rect 56324 5108 56376 5160
rect 55772 5040 55824 5092
rect 56232 5040 56284 5092
rect 56600 5108 56652 5160
rect 57244 5151 57296 5160
rect 57244 5117 57253 5151
rect 57253 5117 57287 5151
rect 57287 5117 57296 5151
rect 57244 5108 57296 5117
rect 57612 5108 57664 5160
rect 59912 5108 59964 5160
rect 60372 5108 60424 5160
rect 60740 5108 60792 5160
rect 61384 5151 61436 5160
rect 61384 5117 61393 5151
rect 61393 5117 61427 5151
rect 61427 5117 61436 5151
rect 61384 5108 61436 5117
rect 61292 5040 61344 5092
rect 62028 5108 62080 5160
rect 62120 5108 62172 5160
rect 62764 5108 62816 5160
rect 63040 5108 63092 5160
rect 63592 5108 63644 5160
rect 63868 5108 63920 5160
rect 65156 5151 65208 5160
rect 65156 5117 65165 5151
rect 65165 5117 65199 5151
rect 65199 5117 65208 5151
rect 65156 5108 65208 5117
rect 65616 5108 65668 5160
rect 65892 5108 65944 5160
rect 66628 5108 66680 5160
rect 51540 5015 51592 5024
rect 51540 4981 51549 5015
rect 51549 4981 51583 5015
rect 51583 4981 51592 5015
rect 51540 4972 51592 4981
rect 52000 4972 52052 5024
rect 58716 5015 58768 5024
rect 58716 4981 58725 5015
rect 58725 4981 58759 5015
rect 58759 4981 58768 5015
rect 58716 4972 58768 4981
rect 59544 4972 59596 5024
rect 66352 5040 66404 5092
rect 68744 5040 68796 5092
rect 66996 4972 67048 5024
rect 69664 4972 69716 5024
rect 9246 4870 9298 4922
rect 9310 4870 9362 4922
rect 9374 4870 9426 4922
rect 9438 4870 9490 4922
rect 23848 4904 23900 4956
rect 33048 4904 33100 4956
rect 24492 4879 24544 4888
rect 24492 4845 24501 4879
rect 24501 4845 24535 4879
rect 24535 4845 24544 4879
rect 24492 4836 24544 4845
rect 31760 4879 31812 4888
rect 31760 4845 31769 4879
rect 31769 4845 31803 4879
rect 31803 4845 31812 4879
rect 32036 4879 32088 4888
rect 31760 4836 31812 4845
rect 32036 4845 32045 4879
rect 32045 4845 32079 4879
rect 32079 4845 32088 4879
rect 32036 4836 32088 4845
rect 32312 4879 32364 4888
rect 32312 4845 32321 4879
rect 32321 4845 32355 4879
rect 32355 4845 32364 4879
rect 32312 4836 32364 4845
rect 32496 4879 32548 4888
rect 32496 4845 32505 4879
rect 32505 4845 32539 4879
rect 32539 4845 32548 4879
rect 32496 4836 32548 4845
rect 39246 4870 39298 4922
rect 39310 4870 39362 4922
rect 39374 4870 39426 4922
rect 39438 4870 39490 4922
rect 49246 4870 49298 4922
rect 49310 4870 49362 4922
rect 49374 4870 49426 4922
rect 49438 4870 49490 4922
rect 59246 4870 59298 4922
rect 59310 4870 59362 4922
rect 59374 4870 59426 4922
rect 59438 4870 59490 4922
rect 7012 4768 7064 4820
rect 7748 4768 7800 4820
rect 10784 4768 10836 4820
rect 3976 4700 4028 4752
rect 13636 4700 13688 4752
rect 2504 4632 2556 4684
rect 3240 4632 3292 4684
rect 4620 4675 4672 4684
rect 4620 4641 4629 4675
rect 4629 4641 4663 4675
rect 4663 4641 4672 4675
rect 4620 4632 4672 4641
rect 4988 4632 5040 4684
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 6000 4632 6052 4684
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 7380 4632 7432 4684
rect 7564 4632 7616 4684
rect 7932 4632 7984 4684
rect 8760 4632 8812 4684
rect 9220 4632 9272 4684
rect 9588 4632 9640 4684
rect 10784 4632 10836 4684
rect 11428 4632 11480 4684
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 12256 4632 12308 4684
rect 1952 4564 2004 4616
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 13544 4632 13596 4684
rect 14096 4632 14148 4684
rect 16028 4700 16080 4752
rect 16488 4768 16540 4820
rect 51908 4768 51960 4820
rect 52276 4768 52328 4820
rect 62672 4768 62724 4820
rect 15200 4632 15252 4684
rect 16304 4632 16356 4684
rect 13360 4564 13412 4616
rect 16672 4564 16724 4616
rect 14648 4496 14700 4548
rect 15200 4496 15252 4548
rect 16856 4539 16908 4548
rect 16856 4505 16865 4539
rect 16865 4505 16899 4539
rect 16899 4505 16908 4539
rect 16856 4496 16908 4505
rect 17224 4700 17276 4752
rect 59360 4700 59412 4752
rect 60648 4700 60700 4752
rect 18788 4632 18840 4684
rect 23756 4632 23808 4684
rect 24400 4632 24452 4684
rect 31944 4675 31996 4684
rect 31944 4641 31953 4675
rect 31953 4641 31987 4675
rect 31987 4641 31996 4675
rect 31944 4632 31996 4641
rect 37556 4632 37608 4684
rect 39672 4632 39724 4684
rect 39856 4675 39908 4684
rect 39856 4641 39865 4675
rect 39865 4641 39899 4675
rect 39899 4641 39908 4675
rect 39856 4632 39908 4641
rect 41052 4632 41104 4684
rect 42616 4632 42668 4684
rect 42892 4675 42944 4684
rect 42892 4641 42901 4675
rect 42901 4641 42935 4675
rect 42935 4641 42944 4675
rect 42892 4632 42944 4641
rect 18512 4564 18564 4616
rect 34612 4564 34664 4616
rect 45928 4632 45980 4684
rect 46112 4632 46164 4684
rect 46388 4632 46440 4684
rect 47400 4675 47452 4684
rect 47400 4641 47409 4675
rect 47409 4641 47443 4675
rect 47443 4641 47452 4675
rect 47400 4632 47452 4641
rect 48044 4675 48096 4684
rect 48044 4641 48053 4675
rect 48053 4641 48087 4675
rect 48087 4641 48096 4675
rect 48044 4632 48096 4641
rect 48136 4632 48188 4684
rect 49240 4632 49292 4684
rect 50344 4632 50396 4684
rect 50804 4632 50856 4684
rect 51448 4675 51500 4684
rect 51448 4641 51457 4675
rect 51457 4641 51491 4675
rect 51491 4641 51500 4675
rect 51448 4632 51500 4641
rect 52184 4632 52236 4684
rect 52828 4632 52880 4684
rect 53196 4632 53248 4684
rect 53932 4632 53984 4684
rect 54576 4632 54628 4684
rect 55404 4632 55456 4684
rect 56140 4632 56192 4684
rect 56692 4632 56744 4684
rect 56876 4675 56928 4684
rect 56876 4641 56885 4675
rect 56885 4641 56919 4675
rect 56919 4641 56928 4675
rect 56876 4632 56928 4641
rect 57060 4632 57112 4684
rect 57520 4675 57572 4684
rect 57520 4641 57529 4675
rect 57529 4641 57563 4675
rect 57563 4641 57572 4675
rect 57520 4632 57572 4641
rect 57888 4632 57940 4684
rect 58624 4632 58676 4684
rect 58900 4632 58952 4684
rect 59728 4675 59780 4684
rect 59728 4641 59737 4675
rect 59737 4641 59771 4675
rect 59771 4641 59780 4675
rect 59728 4632 59780 4641
rect 60096 4632 60148 4684
rect 62396 4675 62448 4684
rect 62396 4641 62405 4675
rect 62405 4641 62439 4675
rect 62439 4641 62448 4675
rect 62396 4632 62448 4641
rect 62488 4632 62540 4684
rect 63316 4632 63368 4684
rect 63868 4632 63920 4684
rect 64144 4632 64196 4684
rect 64696 4675 64748 4684
rect 64696 4641 64705 4675
rect 64705 4641 64739 4675
rect 64739 4641 64748 4675
rect 64696 4632 64748 4641
rect 64788 4632 64840 4684
rect 65248 4632 65300 4684
rect 60188 4564 60240 4616
rect 60648 4564 60700 4616
rect 17040 4496 17092 4548
rect 17224 4496 17276 4548
rect 17592 4496 17644 4548
rect 21456 4496 21508 4548
rect 35072 4496 35124 4548
rect 38844 4496 38896 4548
rect 40224 4496 40276 4548
rect 41052 4496 41104 4548
rect 41328 4496 41380 4548
rect 43444 4496 43496 4548
rect 46112 4496 46164 4548
rect 46204 4496 46256 4548
rect 64236 4496 64288 4548
rect 67824 4539 67876 4548
rect 67824 4505 67833 4539
rect 67833 4505 67867 4539
rect 67867 4505 67876 4539
rect 67824 4496 67876 4505
rect 43076 4428 43128 4480
rect 45652 4428 45704 4480
rect 46388 4428 46440 4480
rect 46756 4428 46808 4480
rect 47676 4428 47728 4480
rect 53932 4428 53984 4480
rect 54852 4428 54904 4480
rect 56232 4471 56284 4480
rect 56232 4437 56241 4471
rect 56241 4437 56275 4471
rect 56275 4437 56284 4471
rect 56232 4428 56284 4437
rect 56876 4428 56928 4480
rect 57888 4428 57940 4480
rect 59360 4428 59412 4480
rect 64052 4428 64104 4480
rect 69112 4428 69164 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 14246 4326 14298 4378
rect 14310 4326 14362 4378
rect 14374 4326 14426 4378
rect 14438 4326 14490 4378
rect 33048 4360 33100 4412
rect 35164 4360 35216 4412
rect 44246 4326 44298 4378
rect 44310 4326 44362 4378
rect 44374 4326 44426 4378
rect 44438 4326 44490 4378
rect 54246 4326 54298 4378
rect 54310 4326 54362 4378
rect 54374 4326 54426 4378
rect 54438 4326 54490 4378
rect 64246 4326 64298 4378
rect 64310 4326 64362 4378
rect 64374 4326 64426 4378
rect 64438 4326 64490 4378
rect 11428 4224 11480 4276
rect 16580 4224 16632 4276
rect 16672 4224 16724 4276
rect 18328 4224 18380 4276
rect 23296 4224 23348 4276
rect 6828 4156 6880 4208
rect 10968 4156 11020 4208
rect 12164 4156 12216 4208
rect 13636 4156 13688 4208
rect 19984 4156 20036 4208
rect 388 4088 440 4140
rect 1492 4088 1544 4140
rect 2136 4088 2188 4140
rect 3240 4088 3292 4140
rect 3976 4088 4028 4140
rect 4620 4088 4672 4140
rect 848 4020 900 4072
rect 2228 4020 2280 4072
rect 2412 4020 2464 4072
rect 2504 4020 2556 4072
rect 3148 4020 3200 4072
rect 572 3952 624 4004
rect 1676 3952 1728 4004
rect 3056 3952 3108 4004
rect 3516 4020 3568 4072
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 5080 4088 5132 4140
rect 8760 4088 8812 4140
rect 9496 4088 9548 4140
rect 11428 4088 11480 4140
rect 11888 4088 11940 4140
rect 11980 4088 12032 4140
rect 12440 4088 12492 4140
rect 12716 4088 12768 4140
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 6276 4020 6328 4072
rect 6460 4020 6512 4072
rect 6920 4020 6972 4072
rect 7380 4020 7432 4072
rect 7932 4020 7984 4072
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8944 4020 8996 4072
rect 4620 3952 4672 4004
rect 8208 3952 8260 4004
rect 940 3884 992 3936
rect 1952 3884 2004 3936
rect 2228 3884 2280 3936
rect 2412 3884 2464 3936
rect 3424 3884 3476 3936
rect 10692 4020 10744 4072
rect 10876 4020 10928 4072
rect 11520 4020 11572 4072
rect 12164 4020 12216 4072
rect 18144 4088 18196 4140
rect 23296 4088 23348 4140
rect 24952 4088 25004 4140
rect 40132 4224 40184 4276
rect 41788 4224 41840 4276
rect 42524 4224 42576 4276
rect 42616 4224 42668 4276
rect 33140 4156 33192 4208
rect 32588 4088 32640 4140
rect 38568 4156 38620 4208
rect 39120 4156 39172 4208
rect 10784 3952 10836 4004
rect 11060 3952 11112 4004
rect 11888 3952 11940 4004
rect 12256 3995 12308 4004
rect 12256 3961 12265 3995
rect 12265 3961 12299 3995
rect 12299 3961 12308 3995
rect 12256 3952 12308 3961
rect 12716 3952 12768 4004
rect 14372 4020 14424 4072
rect 15752 4020 15804 4072
rect 17408 4020 17460 4072
rect 17592 4020 17644 4072
rect 18696 4020 18748 4072
rect 24676 4020 24728 4072
rect 33968 4020 34020 4072
rect 13176 3952 13228 4004
rect 14004 3952 14056 4004
rect 14464 3995 14516 4004
rect 14464 3961 14473 3995
rect 14473 3961 14507 3995
rect 14507 3961 14516 3995
rect 14464 3952 14516 3961
rect 16028 3995 16080 4004
rect 16028 3961 16037 3995
rect 16037 3961 16071 3995
rect 16071 3961 16080 3995
rect 16028 3952 16080 3961
rect 21548 3952 21600 4004
rect 22652 3952 22704 4004
rect 23848 3952 23900 4004
rect 38108 4088 38160 4140
rect 38292 4088 38344 4140
rect 42064 4088 42116 4140
rect 42524 4088 42576 4140
rect 43904 4088 43956 4140
rect 45192 4088 45244 4140
rect 38660 4020 38712 4072
rect 39212 4063 39264 4072
rect 39212 4029 39221 4063
rect 39221 4029 39255 4063
rect 39255 4029 39264 4063
rect 39212 4020 39264 4029
rect 39396 4020 39448 4072
rect 40132 4020 40184 4072
rect 40316 4020 40368 4072
rect 40592 4020 40644 4072
rect 42432 4020 42484 4072
rect 43352 4020 43404 4072
rect 38476 3995 38528 4004
rect 38476 3961 38485 3995
rect 38485 3961 38519 3995
rect 38519 3961 38528 3995
rect 38476 3952 38528 3961
rect 38568 3952 38620 4004
rect 13636 3884 13688 3936
rect 18972 3884 19024 3936
rect 19616 3884 19668 3936
rect 21272 3884 21324 3936
rect 21732 3884 21784 3936
rect 24768 3884 24820 3936
rect 9246 3782 9298 3834
rect 9310 3782 9362 3834
rect 9374 3782 9426 3834
rect 9438 3782 9490 3834
rect 19340 3816 19392 3868
rect 21364 3816 21416 3868
rect 22560 3816 22612 3868
rect 24308 3816 24360 3868
rect 38752 3884 38804 3936
rect 39672 3952 39724 4004
rect 40040 3952 40092 4004
rect 42248 3952 42300 4004
rect 41512 3884 41564 3936
rect 43628 3952 43680 4004
rect 43720 3884 43772 3936
rect 45284 4020 45336 4072
rect 45652 4224 45704 4276
rect 45836 4224 45888 4276
rect 46940 4224 46992 4276
rect 50344 4224 50396 4276
rect 47584 4156 47636 4208
rect 48412 4156 48464 4208
rect 49240 4156 49292 4208
rect 56232 4224 56284 4276
rect 46572 4020 46624 4072
rect 48044 4088 48096 4140
rect 49056 4088 49108 4140
rect 47124 4020 47176 4072
rect 47584 4020 47636 4072
rect 49792 4088 49844 4140
rect 50620 4088 50672 4140
rect 51172 4088 51224 4140
rect 49240 4063 49292 4072
rect 49240 4029 49249 4063
rect 49249 4029 49283 4063
rect 49283 4029 49292 4063
rect 49884 4063 49936 4072
rect 49240 4020 49292 4029
rect 49884 4029 49893 4063
rect 49893 4029 49927 4063
rect 49927 4029 49936 4063
rect 49884 4020 49936 4029
rect 50712 4063 50764 4072
rect 50712 4029 50721 4063
rect 50721 4029 50755 4063
rect 50755 4029 50764 4063
rect 50712 4020 50764 4029
rect 50804 4020 50856 4072
rect 52644 4088 52696 4140
rect 55864 4156 55916 4208
rect 45836 3952 45888 4004
rect 47492 3952 47544 4004
rect 48596 3952 48648 4004
rect 51540 3952 51592 4004
rect 52092 4020 52144 4072
rect 52552 4020 52604 4072
rect 54852 4088 54904 4140
rect 55496 4088 55548 4140
rect 56324 4088 56376 4140
rect 63684 4156 63736 4208
rect 54760 4020 54812 4072
rect 55128 4063 55180 4072
rect 53748 3952 53800 4004
rect 45744 3884 45796 3936
rect 45928 3884 45980 3936
rect 47308 3884 47360 3936
rect 49056 3884 49108 3936
rect 50160 3884 50212 3936
rect 51080 3884 51132 3936
rect 52184 3884 52236 3936
rect 53932 3884 53984 3936
rect 55128 4029 55137 4063
rect 55137 4029 55171 4063
rect 55171 4029 55180 4063
rect 55128 4020 55180 4029
rect 55588 4020 55640 4072
rect 55864 4020 55916 4072
rect 56784 4020 56836 4072
rect 54944 3952 54996 4004
rect 56232 3952 56284 4004
rect 57704 4020 57756 4072
rect 58256 4020 58308 4072
rect 58808 4020 58860 4072
rect 59176 4020 59228 4072
rect 59820 4020 59872 4072
rect 60464 4020 60516 4072
rect 61384 4020 61436 4072
rect 61660 4020 61712 4072
rect 62580 4020 62632 4072
rect 62856 4020 62908 4072
rect 63040 4020 63092 4072
rect 63408 4063 63460 4072
rect 63408 4029 63417 4063
rect 63417 4029 63451 4063
rect 63451 4029 63460 4063
rect 63408 4020 63460 4029
rect 66168 4088 66220 4140
rect 68192 4088 68244 4140
rect 55588 3884 55640 3936
rect 55956 3884 56008 3936
rect 58992 3884 59044 3936
rect 63592 3884 63644 3936
rect 66076 4020 66128 4072
rect 66996 4020 67048 4072
rect 68560 4020 68612 4072
rect 66628 3995 66680 4004
rect 66628 3961 66637 3995
rect 66637 3961 66671 3995
rect 66671 3961 66680 3995
rect 66628 3952 66680 3961
rect 67456 3995 67508 4004
rect 67456 3961 67465 3995
rect 67465 3961 67499 3995
rect 67499 3961 67508 3995
rect 67456 3952 67508 3961
rect 68284 3952 68336 4004
rect 65984 3884 66036 3936
rect 69572 3884 69624 3936
rect 19432 3748 19484 3800
rect 23388 3748 23440 3800
rect 23480 3748 23532 3800
rect 23756 3748 23808 3800
rect 23940 3748 23992 3800
rect 32404 3748 32456 3800
rect 35440 3748 35492 3800
rect 39246 3782 39298 3834
rect 39310 3782 39362 3834
rect 39374 3782 39426 3834
rect 39438 3782 39490 3834
rect 49246 3782 49298 3834
rect 49310 3782 49362 3834
rect 49374 3782 49426 3834
rect 49438 3782 49490 3834
rect 59246 3782 59298 3834
rect 59310 3782 59362 3834
rect 59374 3782 59426 3834
rect 59438 3782 59490 3834
rect 1676 3680 1728 3732
rect 2320 3680 2372 3732
rect 3884 3612 3936 3664
rect 4712 3680 4764 3732
rect 5172 3680 5224 3732
rect 5724 3680 5776 3732
rect 6184 3680 6236 3732
rect 7564 3680 7616 3732
rect 7748 3680 7800 3732
rect 8392 3680 8444 3732
rect 10508 3680 10560 3732
rect 15384 3680 15436 3732
rect 5632 3655 5684 3664
rect 5632 3621 5641 3655
rect 5641 3621 5675 3655
rect 5675 3621 5684 3655
rect 5632 3612 5684 3621
rect 6368 3655 6420 3664
rect 6368 3621 6377 3655
rect 6377 3621 6411 3655
rect 6411 3621 6420 3655
rect 6368 3612 6420 3621
rect 11060 3612 11112 3664
rect 13084 3612 13136 3664
rect 13360 3655 13412 3664
rect 13360 3621 13369 3655
rect 13369 3621 13403 3655
rect 13403 3621 13412 3655
rect 13360 3612 13412 3621
rect 13544 3612 13596 3664
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 20 3476 72 3528
rect 1124 3476 1176 3528
rect 1400 3476 1452 3528
rect 2596 3544 2648 3596
rect 664 3408 716 3460
rect 1768 3408 1820 3460
rect 1952 3408 2004 3460
rect 3608 3544 3660 3596
rect 6736 3544 6788 3596
rect 5632 3476 5684 3528
rect 6092 3476 6144 3528
rect 7656 3544 7708 3596
rect 8024 3544 8076 3596
rect 10140 3544 10192 3596
rect 11152 3544 11204 3596
rect 15108 3587 15160 3596
rect 15108 3553 15117 3587
rect 15117 3553 15151 3587
rect 15151 3553 15160 3587
rect 15108 3544 15160 3553
rect 18144 3680 18196 3732
rect 18236 3680 18288 3732
rect 16396 3612 16448 3664
rect 17224 3612 17276 3664
rect 17960 3612 18012 3664
rect 16672 3544 16724 3596
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 17868 3544 17920 3596
rect 19708 3612 19760 3664
rect 20628 3544 20680 3596
rect 20996 3680 21048 3732
rect 33048 3680 33100 3732
rect 33968 3680 34020 3732
rect 35532 3680 35584 3732
rect 37280 3680 37332 3732
rect 38292 3680 38344 3732
rect 38568 3680 38620 3732
rect 21640 3612 21692 3664
rect 31668 3612 31720 3664
rect 36360 3612 36412 3664
rect 22652 3544 22704 3596
rect 24216 3544 24268 3596
rect 35072 3544 35124 3596
rect 35164 3544 35216 3596
rect 37188 3544 37240 3596
rect 37556 3612 37608 3664
rect 37648 3612 37700 3664
rect 39028 3587 39080 3596
rect 39028 3553 39037 3587
rect 39037 3553 39071 3587
rect 39071 3553 39080 3587
rect 39028 3544 39080 3553
rect 39212 3587 39264 3596
rect 39212 3553 39221 3587
rect 39221 3553 39255 3587
rect 39255 3553 39264 3587
rect 39212 3544 39264 3553
rect 40684 3612 40736 3664
rect 42156 3655 42208 3664
rect 42156 3621 42165 3655
rect 42165 3621 42199 3655
rect 42199 3621 42208 3655
rect 42156 3612 42208 3621
rect 42892 3680 42944 3732
rect 45192 3680 45244 3732
rect 46388 3680 46440 3732
rect 47216 3680 47268 3732
rect 48504 3680 48556 3732
rect 50160 3680 50212 3732
rect 51448 3680 51500 3732
rect 61660 3680 61712 3732
rect 62396 3680 62448 3732
rect 63960 3680 64012 3732
rect 3792 3408 3844 3460
rect 4804 3408 4856 3460
rect 6920 3408 6972 3460
rect 8944 3408 8996 3460
rect 5080 3340 5132 3392
rect 8024 3340 8076 3392
rect 8852 3340 8904 3392
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 10232 3340 10284 3392
rect 10600 3340 10652 3392
rect 11060 3340 11112 3392
rect 12256 3476 12308 3528
rect 15384 3476 15436 3528
rect 15936 3476 15988 3528
rect 20904 3476 20956 3528
rect 23480 3476 23532 3528
rect 32772 3476 32824 3528
rect 40868 3544 40920 3596
rect 42064 3544 42116 3596
rect 42340 3544 42392 3596
rect 43260 3544 43312 3596
rect 43720 3544 43772 3596
rect 45468 3612 45520 3664
rect 45652 3655 45704 3664
rect 45652 3621 45661 3655
rect 45661 3621 45695 3655
rect 45695 3621 45704 3655
rect 45652 3612 45704 3621
rect 45100 3544 45152 3596
rect 12440 3340 12492 3392
rect 13360 3340 13412 3392
rect 17960 3340 18012 3392
rect 19064 3408 19116 3460
rect 22652 3408 22704 3460
rect 23664 3408 23716 3460
rect 39120 3408 39172 3460
rect 39212 3408 39264 3460
rect 39488 3408 39540 3460
rect 42248 3476 42300 3528
rect 42800 3476 42852 3528
rect 44824 3476 44876 3528
rect 45744 3476 45796 3528
rect 19156 3340 19208 3392
rect 20904 3340 20956 3392
rect 21456 3340 21508 3392
rect 23940 3340 23992 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 14246 3238 14298 3290
rect 14310 3238 14362 3290
rect 14374 3238 14426 3290
rect 14438 3238 14490 3290
rect 38752 3340 38804 3392
rect 39856 3340 39908 3392
rect 43904 3408 43956 3460
rect 47124 3612 47176 3664
rect 47676 3655 47728 3664
rect 47676 3621 47685 3655
rect 47685 3621 47719 3655
rect 47719 3621 47728 3655
rect 47676 3612 47728 3621
rect 48136 3612 48188 3664
rect 46572 3544 46624 3596
rect 48228 3587 48280 3596
rect 46388 3476 46440 3528
rect 48228 3553 48237 3587
rect 48237 3553 48271 3587
rect 48271 3553 48280 3587
rect 48228 3544 48280 3553
rect 47308 3476 47360 3528
rect 48964 3544 49016 3596
rect 50068 3544 50120 3596
rect 52000 3612 52052 3664
rect 53380 3612 53432 3664
rect 54116 3612 54168 3664
rect 55680 3612 55732 3664
rect 57152 3612 57204 3664
rect 57428 3655 57480 3664
rect 57428 3621 57437 3655
rect 57437 3621 57471 3655
rect 57471 3621 57480 3655
rect 57428 3612 57480 3621
rect 49148 3476 49200 3528
rect 51264 3544 51316 3596
rect 51816 3544 51868 3596
rect 53012 3544 53064 3596
rect 57980 3544 58032 3596
rect 58716 3544 58768 3596
rect 58808 3544 58860 3596
rect 59544 3612 59596 3664
rect 61752 3612 61804 3664
rect 65984 3680 66036 3732
rect 66536 3680 66588 3732
rect 64880 3612 64932 3664
rect 65524 3612 65576 3664
rect 66812 3612 66864 3664
rect 67364 3612 67416 3664
rect 46572 3451 46624 3460
rect 46572 3417 46581 3451
rect 46581 3417 46615 3451
rect 46615 3417 46624 3451
rect 46572 3408 46624 3417
rect 47492 3451 47544 3460
rect 47492 3417 47501 3451
rect 47501 3417 47535 3451
rect 47535 3417 47544 3451
rect 47492 3408 47544 3417
rect 47676 3408 47728 3460
rect 41328 3340 41380 3392
rect 42708 3340 42760 3392
rect 42800 3340 42852 3392
rect 45744 3340 45796 3392
rect 50068 3340 50120 3392
rect 50344 3408 50396 3460
rect 51356 3476 51408 3528
rect 52276 3476 52328 3528
rect 53288 3476 53340 3528
rect 54760 3476 54812 3528
rect 57796 3476 57848 3528
rect 60004 3544 60056 3596
rect 60096 3544 60148 3596
rect 60556 3544 60608 3596
rect 60924 3544 60976 3596
rect 62304 3544 62356 3596
rect 62672 3544 62724 3596
rect 63224 3544 63276 3596
rect 61752 3476 61804 3528
rect 66812 3476 66864 3528
rect 67272 3476 67324 3528
rect 68284 3476 68336 3528
rect 51448 3408 51500 3460
rect 51724 3408 51776 3460
rect 52552 3451 52604 3460
rect 52552 3417 52561 3451
rect 52561 3417 52595 3451
rect 52595 3417 52604 3451
rect 52552 3408 52604 3417
rect 53380 3451 53432 3460
rect 53380 3417 53389 3451
rect 53389 3417 53423 3451
rect 53423 3417 53432 3451
rect 53380 3408 53432 3417
rect 54116 3408 54168 3460
rect 55128 3451 55180 3460
rect 55128 3417 55137 3451
rect 55137 3417 55171 3451
rect 55171 3417 55180 3451
rect 55128 3408 55180 3417
rect 56416 3408 56468 3460
rect 57244 3451 57296 3460
rect 57244 3417 57253 3451
rect 57253 3417 57287 3451
rect 57287 3417 57296 3451
rect 57244 3408 57296 3417
rect 64052 3451 64104 3460
rect 64052 3417 64061 3451
rect 64061 3417 64095 3451
rect 64095 3417 64104 3451
rect 64052 3408 64104 3417
rect 64880 3451 64932 3460
rect 64880 3417 64889 3451
rect 64889 3417 64923 3451
rect 64923 3417 64932 3451
rect 64880 3408 64932 3417
rect 65800 3408 65852 3460
rect 66352 3408 66404 3460
rect 66996 3408 67048 3460
rect 50528 3340 50580 3392
rect 50804 3340 50856 3392
rect 51080 3340 51132 3392
rect 51172 3340 51224 3392
rect 51816 3340 51868 3392
rect 52368 3340 52420 3392
rect 53196 3340 53248 3392
rect 53748 3340 53800 3392
rect 58532 3340 58584 3392
rect 66168 3340 66220 3392
rect 35532 3272 35584 3324
rect 19064 3204 19116 3256
rect 21640 3204 21692 3256
rect 33876 3204 33928 3256
rect 35348 3204 35400 3256
rect 35440 3204 35492 3256
rect 37096 3204 37148 3256
rect 44246 3238 44298 3290
rect 44310 3238 44362 3290
rect 44374 3238 44426 3290
rect 44438 3238 44490 3290
rect 54246 3238 54298 3290
rect 54310 3238 54362 3290
rect 54374 3238 54426 3290
rect 54438 3238 54490 3290
rect 64246 3238 64298 3290
rect 64310 3238 64362 3290
rect 64374 3238 64426 3290
rect 64438 3238 64490 3290
rect 2872 3136 2924 3188
rect 3332 3136 3384 3188
rect 10692 3136 10744 3188
rect 2780 3068 2832 3120
rect 8116 3068 8168 3120
rect 2228 3000 2280 3052
rect 4160 3000 4212 3052
rect 4712 3000 4764 3052
rect 1676 2932 1728 2984
rect 3700 2932 3752 2984
rect 5816 3000 5868 3052
rect 8484 3000 8536 3052
rect 5540 2932 5592 2984
rect 7196 2932 7248 2984
rect 8116 2932 8168 2984
rect 8668 2975 8720 2984
rect 8668 2941 8677 2975
rect 8677 2941 8711 2975
rect 8711 2941 8720 2975
rect 8668 2932 8720 2941
rect 2320 2864 2372 2916
rect 4068 2864 4120 2916
rect 5264 2864 5316 2916
rect 6552 2864 6604 2916
rect 8484 2907 8536 2916
rect 8484 2873 8493 2907
rect 8493 2873 8527 2907
rect 8527 2873 8536 2907
rect 8484 2864 8536 2873
rect 112 2796 164 2848
rect 1584 2796 1636 2848
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 2872 2796 2924 2848
rect 3700 2796 3752 2848
rect 5816 2796 5868 2848
rect 7012 2796 7064 2848
rect 8852 2932 8904 2984
rect 10140 3000 10192 3052
rect 11520 3068 11572 3120
rect 13544 3136 13596 3188
rect 23664 3136 23716 3188
rect 24492 3136 24544 3188
rect 21088 3068 21140 3120
rect 24400 3068 24452 3120
rect 34704 3136 34756 3188
rect 18512 3000 18564 3052
rect 18604 3000 18656 3052
rect 24952 3000 25004 3052
rect 35072 3068 35124 3120
rect 40040 3136 40092 3188
rect 40316 3136 40368 3188
rect 41420 3136 41472 3188
rect 41880 3136 41932 3188
rect 45652 3136 45704 3188
rect 47400 3136 47452 3188
rect 39764 3111 39816 3120
rect 39764 3077 39773 3111
rect 39773 3077 39807 3111
rect 39807 3077 39816 3111
rect 39764 3068 39816 3077
rect 39120 3000 39172 3052
rect 40132 3000 40184 3052
rect 10508 2932 10560 2984
rect 10600 2932 10652 2984
rect 12808 2932 12860 2984
rect 14004 2975 14056 2984
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 15016 2932 15068 2984
rect 15936 2932 15988 2984
rect 16212 2975 16264 2984
rect 16212 2941 16221 2975
rect 16221 2941 16255 2975
rect 16255 2941 16264 2975
rect 16212 2932 16264 2941
rect 16304 2932 16356 2984
rect 17500 2975 17552 2984
rect 8944 2864 8996 2916
rect 9772 2864 9824 2916
rect 10876 2907 10928 2916
rect 10876 2873 10885 2907
rect 10885 2873 10919 2907
rect 10919 2873 10928 2907
rect 10876 2864 10928 2873
rect 11796 2864 11848 2916
rect 16396 2864 16448 2916
rect 17500 2941 17509 2975
rect 17509 2941 17543 2975
rect 17543 2941 17552 2975
rect 17500 2932 17552 2941
rect 17960 2932 18012 2984
rect 22560 2932 22612 2984
rect 31852 2932 31904 2984
rect 17868 2864 17920 2916
rect 12808 2796 12860 2848
rect 15476 2839 15528 2848
rect 15476 2805 15485 2839
rect 15485 2805 15519 2839
rect 15519 2805 15528 2839
rect 15476 2796 15528 2805
rect 16120 2796 16172 2848
rect 17500 2796 17552 2848
rect 20260 2864 20312 2916
rect 20352 2864 20404 2916
rect 23572 2864 23624 2916
rect 31668 2864 31720 2916
rect 32956 2932 33008 2984
rect 37464 2932 37516 2984
rect 39212 2975 39264 2984
rect 39212 2941 39221 2975
rect 39221 2941 39255 2975
rect 39255 2941 39264 2975
rect 39212 2932 39264 2941
rect 39948 2975 40000 2984
rect 39948 2941 39957 2975
rect 39957 2941 39991 2975
rect 39991 2941 40000 2975
rect 39948 2932 40000 2941
rect 18696 2796 18748 2848
rect 9246 2694 9298 2746
rect 9310 2694 9362 2746
rect 9374 2694 9426 2746
rect 9438 2694 9490 2746
rect 16304 2592 16356 2644
rect 19800 2796 19852 2848
rect 21180 2796 21232 2848
rect 23388 2839 23440 2848
rect 23388 2805 23397 2839
rect 23397 2805 23431 2839
rect 23431 2805 23440 2839
rect 23388 2796 23440 2805
rect 24124 2796 24176 2848
rect 22744 2660 22796 2712
rect 23112 2660 23164 2712
rect 23388 2703 23440 2712
rect 23388 2669 23397 2703
rect 23397 2669 23431 2703
rect 23431 2669 23440 2703
rect 23388 2660 23440 2669
rect 31852 2660 31904 2712
rect 32036 2728 32088 2780
rect 24032 2592 24084 2644
rect 1124 2524 1176 2576
rect 5356 2524 5408 2576
rect 5908 2567 5960 2576
rect 5908 2533 5917 2567
rect 5917 2533 5951 2567
rect 5951 2533 5960 2567
rect 5908 2524 5960 2533
rect 7104 2567 7156 2576
rect 7104 2533 7113 2567
rect 7113 2533 7147 2567
rect 7147 2533 7156 2567
rect 7104 2524 7156 2533
rect 7840 2567 7892 2576
rect 7840 2533 7849 2567
rect 7849 2533 7883 2567
rect 7883 2533 7892 2567
rect 7840 2524 7892 2533
rect 8576 2567 8628 2576
rect 8576 2533 8585 2567
rect 8585 2533 8619 2567
rect 8619 2533 8628 2567
rect 8576 2524 8628 2533
rect 9772 2567 9824 2576
rect 9772 2533 9781 2567
rect 9781 2533 9815 2567
rect 9815 2533 9824 2567
rect 9772 2524 9824 2533
rect 10692 2524 10744 2576
rect 12348 2567 12400 2576
rect 12348 2533 12357 2567
rect 12357 2533 12391 2567
rect 12391 2533 12400 2567
rect 12348 2524 12400 2533
rect 13084 2567 13136 2576
rect 13084 2533 13093 2567
rect 13093 2533 13127 2567
rect 13127 2533 13136 2567
rect 13084 2524 13136 2533
rect 13820 2567 13872 2576
rect 13820 2533 13829 2567
rect 13829 2533 13863 2567
rect 13863 2533 13872 2567
rect 13820 2524 13872 2533
rect 15384 2524 15436 2576
rect 16764 2524 16816 2576
rect 18420 2524 18472 2576
rect 18788 2524 18840 2576
rect 32036 2524 32088 2576
rect 32128 2524 32180 2576
rect 32588 2864 32640 2916
rect 42892 3068 42944 3120
rect 44916 3068 44968 3120
rect 45284 3068 45336 3120
rect 40500 3043 40552 3052
rect 40500 3009 40509 3043
rect 40509 3009 40543 3043
rect 40543 3009 40552 3043
rect 40500 3000 40552 3009
rect 40776 3000 40828 3052
rect 44088 3000 44140 3052
rect 46112 3000 46164 3052
rect 40684 2975 40736 2984
rect 40684 2941 40693 2975
rect 40693 2941 40727 2975
rect 40727 2941 40736 2975
rect 40684 2932 40736 2941
rect 41420 2975 41472 2984
rect 41420 2941 41429 2975
rect 41429 2941 41463 2975
rect 41463 2941 41472 2975
rect 41420 2932 41472 2941
rect 41972 2975 42024 2984
rect 41972 2941 41981 2975
rect 41981 2941 42015 2975
rect 42015 2941 42024 2975
rect 41972 2932 42024 2941
rect 40500 2864 40552 2916
rect 43168 2932 43220 2984
rect 43720 2932 43772 2984
rect 44640 2932 44692 2984
rect 46480 2975 46532 2984
rect 46480 2941 46489 2975
rect 46489 2941 46523 2975
rect 46523 2941 46532 2975
rect 47768 3000 47820 3052
rect 46480 2932 46532 2941
rect 48228 3000 48280 3052
rect 48504 3000 48556 3052
rect 62856 3136 62908 3188
rect 48780 3068 48832 3120
rect 48688 2932 48740 2984
rect 42432 2864 42484 2916
rect 32772 2796 32824 2848
rect 32956 2839 33008 2848
rect 32956 2805 32965 2839
rect 32965 2805 32999 2839
rect 32999 2805 33008 2839
rect 32956 2796 33008 2805
rect 40132 2796 40184 2848
rect 41788 2796 41840 2848
rect 42984 2796 43036 2848
rect 43260 2796 43312 2848
rect 45008 2907 45060 2916
rect 45008 2873 45017 2907
rect 45017 2873 45051 2907
rect 45051 2873 45060 2907
rect 45008 2864 45060 2873
rect 45468 2864 45520 2916
rect 47860 2864 47912 2916
rect 44916 2796 44968 2848
rect 47032 2796 47084 2848
rect 49792 3068 49844 3120
rect 50528 3068 50580 3120
rect 54208 3068 54260 3120
rect 62764 3068 62816 3120
rect 65800 3068 65852 3120
rect 66076 3136 66128 3188
rect 69388 3136 69440 3188
rect 68100 3111 68152 3120
rect 68100 3077 68109 3111
rect 68109 3077 68143 3111
rect 68143 3077 68152 3111
rect 68100 3068 68152 3077
rect 50896 3000 50948 3052
rect 51724 3000 51776 3052
rect 53840 3000 53892 3052
rect 55496 3000 55548 3052
rect 50252 2975 50304 2984
rect 50252 2941 50261 2975
rect 50261 2941 50295 2975
rect 50295 2941 50304 2975
rect 50252 2932 50304 2941
rect 51356 2932 51408 2984
rect 49240 2864 49292 2916
rect 49608 2864 49660 2916
rect 51908 2932 51960 2984
rect 52460 2975 52512 2984
rect 52460 2941 52469 2975
rect 52469 2941 52503 2975
rect 52503 2941 52512 2975
rect 52460 2932 52512 2941
rect 54024 2975 54076 2984
rect 54024 2941 54033 2975
rect 54033 2941 54067 2975
rect 54067 2941 54076 2975
rect 54024 2932 54076 2941
rect 54668 2932 54720 2984
rect 56784 2932 56836 2984
rect 58348 2932 58400 2984
rect 63224 3000 63276 3052
rect 67916 3000 67968 3052
rect 51816 2864 51868 2916
rect 52920 2864 52972 2916
rect 53012 2864 53064 2916
rect 55220 2864 55272 2916
rect 56048 2864 56100 2916
rect 56324 2864 56376 2916
rect 57336 2864 57388 2916
rect 58992 2864 59044 2916
rect 60280 2932 60332 2984
rect 61200 2975 61252 2984
rect 61200 2941 61209 2975
rect 61209 2941 61243 2975
rect 61243 2941 61252 2975
rect 61200 2932 61252 2941
rect 62212 2932 62264 2984
rect 63960 2932 64012 2984
rect 64972 2932 65024 2984
rect 65708 2932 65760 2984
rect 59820 2864 59872 2916
rect 61016 2907 61068 2916
rect 61016 2873 61025 2907
rect 61025 2873 61059 2907
rect 61059 2873 61068 2907
rect 61016 2864 61068 2873
rect 62304 2907 62356 2916
rect 62304 2873 62313 2907
rect 62313 2873 62347 2907
rect 62347 2873 62356 2907
rect 62304 2864 62356 2873
rect 63132 2864 63184 2916
rect 63592 2864 63644 2916
rect 64696 2864 64748 2916
rect 65340 2864 65392 2916
rect 67088 2864 67140 2916
rect 48964 2796 49016 2848
rect 49976 2796 50028 2848
rect 51264 2796 51316 2848
rect 54484 2796 54536 2848
rect 54760 2796 54812 2848
rect 55956 2796 56008 2848
rect 62212 2796 62264 2848
rect 62672 2796 62724 2848
rect 65708 2796 65760 2848
rect 1584 2456 1636 2508
rect 6368 2456 6420 2508
rect 7656 2456 7708 2508
rect 10232 2456 10284 2508
rect 13912 2456 13964 2508
rect 14096 2456 14148 2508
rect 18604 2456 18656 2508
rect 31668 2456 31720 2508
rect 33324 2703 33376 2712
rect 33324 2669 33333 2703
rect 33333 2669 33367 2703
rect 33367 2669 33376 2703
rect 33324 2660 33376 2669
rect 36728 2660 36780 2712
rect 39246 2694 39298 2746
rect 39310 2694 39362 2746
rect 39374 2694 39426 2746
rect 39438 2694 39490 2746
rect 49246 2694 49298 2746
rect 49310 2694 49362 2746
rect 49374 2694 49426 2746
rect 49438 2694 49490 2746
rect 59246 2694 59298 2746
rect 59310 2694 59362 2746
rect 59374 2694 59426 2746
rect 59438 2694 59490 2746
rect 32772 2592 32824 2644
rect 48504 2592 48556 2644
rect 49792 2592 49844 2644
rect 54208 2635 54260 2644
rect 54208 2601 54217 2635
rect 54217 2601 54251 2635
rect 54251 2601 54260 2635
rect 54208 2592 54260 2601
rect 57520 2592 57572 2644
rect 58532 2592 58584 2644
rect 60648 2592 60700 2644
rect 66352 2592 66404 2644
rect 33416 2567 33468 2576
rect 33416 2533 33425 2567
rect 33425 2533 33459 2567
rect 33459 2533 33468 2567
rect 33416 2524 33468 2533
rect 33692 2524 33744 2576
rect 38936 2524 38988 2576
rect 39856 2524 39908 2576
rect 40316 2524 40368 2576
rect 40960 2567 41012 2576
rect 40960 2533 40969 2567
rect 40969 2533 41003 2567
rect 41003 2533 41012 2567
rect 40960 2524 41012 2533
rect 42432 2567 42484 2576
rect 42432 2533 42441 2567
rect 42441 2533 42475 2567
rect 42475 2533 42484 2567
rect 42432 2524 42484 2533
rect 43168 2524 43220 2576
rect 44548 2524 44600 2576
rect 46020 2524 46072 2576
rect 46296 2567 46348 2576
rect 46296 2533 46305 2567
rect 46305 2533 46339 2567
rect 46339 2533 46348 2567
rect 46296 2524 46348 2533
rect 46664 2524 46716 2576
rect 48320 2524 48372 2576
rect 48688 2524 48740 2576
rect 48872 2524 48924 2576
rect 49700 2567 49752 2576
rect 49700 2533 49709 2567
rect 49709 2533 49743 2567
rect 49743 2533 49752 2567
rect 49700 2524 49752 2533
rect 50068 2524 50120 2576
rect 50436 2567 50488 2576
rect 50436 2533 50445 2567
rect 50445 2533 50479 2567
rect 50479 2533 50488 2567
rect 50436 2524 50488 2533
rect 51632 2567 51684 2576
rect 51632 2533 51641 2567
rect 51641 2533 51675 2567
rect 51675 2533 51684 2567
rect 51632 2524 51684 2533
rect 32864 2388 32916 2440
rect 42708 2456 42760 2508
rect 49240 2456 49292 2508
rect 53472 2524 53524 2576
rect 53748 2524 53800 2576
rect 54484 2524 54536 2576
rect 55312 2524 55364 2576
rect 55864 2524 55916 2576
rect 56968 2567 57020 2576
rect 56968 2533 56977 2567
rect 56977 2533 57011 2567
rect 57011 2533 57020 2567
rect 56968 2524 57020 2533
rect 58164 2524 58216 2576
rect 52184 2499 52236 2508
rect 52184 2465 52193 2499
rect 52193 2465 52227 2499
rect 52227 2465 52236 2499
rect 52184 2456 52236 2465
rect 59360 2524 59412 2576
rect 59636 2567 59688 2576
rect 59636 2533 59645 2567
rect 59645 2533 59679 2567
rect 59679 2533 59688 2567
rect 59636 2524 59688 2533
rect 60556 2524 60608 2576
rect 61108 2567 61160 2576
rect 61108 2533 61117 2567
rect 61117 2533 61151 2567
rect 61151 2533 61160 2567
rect 61108 2524 61160 2533
rect 61844 2524 61896 2576
rect 63776 2567 63828 2576
rect 63776 2533 63785 2567
rect 63785 2533 63819 2567
rect 63819 2533 63828 2567
rect 63776 2524 63828 2533
rect 65248 2524 65300 2576
rect 65524 2524 65576 2576
rect 65800 2524 65852 2576
rect 67364 2524 67416 2576
rect 296 2320 348 2372
rect 6368 2320 6420 2372
rect 7288 2320 7340 2372
rect 15108 2363 15160 2372
rect 5908 2252 5960 2304
rect 6736 2252 6788 2304
rect 8116 2252 8168 2304
rect 13728 2252 13780 2304
rect 14096 2252 14148 2304
rect 15108 2329 15117 2363
rect 15117 2329 15151 2363
rect 15151 2329 15160 2363
rect 15108 2320 15160 2329
rect 33600 2363 33652 2372
rect 17592 2252 17644 2304
rect 19432 2252 19484 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 14246 2150 14298 2202
rect 14310 2150 14362 2202
rect 14374 2150 14426 2202
rect 14438 2150 14490 2202
rect 13912 2048 13964 2100
rect 17224 2048 17276 2100
rect 33600 2329 33609 2363
rect 33609 2329 33643 2363
rect 33643 2329 33652 2363
rect 33600 2320 33652 2329
rect 42432 2320 42484 2372
rect 46848 2363 46900 2372
rect 41604 2295 41656 2304
rect 22928 2159 22980 2168
rect 22928 2125 22937 2159
rect 22937 2125 22971 2159
rect 22971 2125 22980 2159
rect 22928 2116 22980 2125
rect 23204 2048 23256 2100
rect 41604 2261 41613 2295
rect 41613 2261 41647 2295
rect 41647 2261 41656 2295
rect 41604 2252 41656 2261
rect 42340 2295 42392 2304
rect 42340 2261 42349 2295
rect 42349 2261 42383 2295
rect 42383 2261 42392 2295
rect 42340 2252 42392 2261
rect 43536 2295 43588 2304
rect 43536 2261 43545 2295
rect 43545 2261 43579 2295
rect 43579 2261 43588 2295
rect 43536 2252 43588 2261
rect 43720 2252 43772 2304
rect 45100 2252 45152 2304
rect 46848 2329 46857 2363
rect 46857 2329 46891 2363
rect 46891 2329 46900 2363
rect 46848 2320 46900 2329
rect 49792 2388 49844 2440
rect 58532 2499 58584 2508
rect 58532 2465 58549 2499
rect 58549 2465 58583 2499
rect 58583 2465 58584 2499
rect 58532 2456 58584 2465
rect 61936 2456 61988 2508
rect 65156 2456 65208 2508
rect 58900 2388 58952 2440
rect 52092 2320 52144 2372
rect 57612 2363 57664 2372
rect 57612 2329 57621 2363
rect 57621 2329 57655 2363
rect 57655 2329 57664 2363
rect 57612 2320 57664 2329
rect 58072 2320 58124 2372
rect 60188 2320 60240 2372
rect 63408 2388 63460 2440
rect 61476 2320 61528 2372
rect 58440 2252 58492 2304
rect 58532 2252 58584 2304
rect 61568 2252 61620 2304
rect 68192 2320 68244 2372
rect 44246 2150 44298 2202
rect 44310 2150 44362 2202
rect 44374 2150 44426 2202
rect 44438 2150 44490 2202
rect 54246 2150 54298 2202
rect 54310 2150 54362 2202
rect 54374 2150 54426 2202
rect 54438 2150 54490 2202
rect 64246 2150 64298 2202
rect 64310 2150 64362 2202
rect 64374 2150 64426 2202
rect 64438 2150 64490 2202
rect 14096 1980 14148 2032
rect 21088 1980 21140 2032
rect 22836 1980 22888 2032
rect 23296 1980 23348 2032
rect 13728 1912 13780 1964
rect 21916 1912 21968 1964
rect 22100 1955 22152 1964
rect 22100 1921 22109 1955
rect 22109 1921 22143 1955
rect 22143 1921 22152 1955
rect 22100 1912 22152 1921
rect 32220 2048 32272 2100
rect 39672 2048 39724 2100
rect 39948 2048 40000 2100
rect 41052 2048 41104 2100
rect 46848 2048 46900 2100
rect 49332 2048 49384 2100
rect 51080 2048 51132 2100
rect 38568 1980 38620 2032
rect 45100 1980 45152 2032
rect 26332 1955 26384 1964
rect 26332 1921 26341 1955
rect 26341 1921 26375 1955
rect 26375 1921 26384 1955
rect 26332 1912 26384 1921
rect 26516 1955 26568 1964
rect 26516 1921 26525 1955
rect 26525 1921 26559 1955
rect 26559 1921 26568 1955
rect 26516 1912 26568 1921
rect 26608 1955 26660 1964
rect 26608 1921 26617 1955
rect 26617 1921 26651 1955
rect 26651 1921 26660 1955
rect 26884 1955 26936 1964
rect 26608 1912 26660 1921
rect 26884 1921 26893 1955
rect 26893 1921 26927 1955
rect 26927 1921 26936 1955
rect 26884 1912 26936 1921
rect 27160 1955 27212 1964
rect 27160 1921 27169 1955
rect 27169 1921 27203 1955
rect 27203 1921 27212 1955
rect 27160 1912 27212 1921
rect 27436 1955 27488 1964
rect 27436 1921 27445 1955
rect 27445 1921 27479 1955
rect 27479 1921 27488 1955
rect 27436 1912 27488 1921
rect 27620 1955 27672 1964
rect 27620 1921 27629 1955
rect 27629 1921 27663 1955
rect 27663 1921 27672 1955
rect 27620 1912 27672 1921
rect 27896 1955 27948 1964
rect 27896 1921 27905 1955
rect 27905 1921 27939 1955
rect 27939 1921 27948 1955
rect 27896 1912 27948 1921
rect 28724 1955 28776 1964
rect 28724 1921 28733 1955
rect 28733 1921 28767 1955
rect 28767 1921 28776 1955
rect 28724 1912 28776 1921
rect 29000 1955 29052 1964
rect 29000 1921 29009 1955
rect 29009 1921 29043 1955
rect 29043 1921 29052 1955
rect 29000 1912 29052 1921
rect 29184 1955 29236 1964
rect 29184 1921 29193 1955
rect 29193 1921 29227 1955
rect 29227 1921 29236 1955
rect 29184 1912 29236 1921
rect 29276 1912 29328 1964
rect 31760 1912 31812 1964
rect 34152 1955 34204 1964
rect 34152 1921 34161 1955
rect 34161 1921 34195 1955
rect 34195 1921 34204 1955
rect 34152 1912 34204 1921
rect 34428 1955 34480 1964
rect 34428 1921 34437 1955
rect 34437 1921 34471 1955
rect 34471 1921 34480 1955
rect 34428 1912 34480 1921
rect 41604 1912 41656 1964
rect 46848 1912 46900 1964
rect 47952 1912 48004 1964
rect 16580 1844 16632 1896
rect 19064 1844 19116 1896
rect 25320 1887 25372 1896
rect 25320 1853 25329 1887
rect 25329 1853 25363 1887
rect 25363 1853 25372 1887
rect 25320 1844 25372 1853
rect 25596 1887 25648 1896
rect 25596 1853 25605 1887
rect 25605 1853 25639 1887
rect 25639 1853 25648 1887
rect 25596 1844 25648 1853
rect 25780 1887 25832 1896
rect 25780 1853 25789 1887
rect 25789 1853 25823 1887
rect 25823 1853 25832 1887
rect 25780 1844 25832 1853
rect 25872 1887 25924 1896
rect 25872 1853 25881 1887
rect 25881 1853 25915 1887
rect 25915 1853 25924 1887
rect 26056 1887 26108 1896
rect 25872 1844 25924 1853
rect 26056 1853 26065 1887
rect 26065 1853 26099 1887
rect 26099 1853 26108 1887
rect 26056 1844 26108 1853
rect 26148 1844 26200 1896
rect 26792 1887 26844 1896
rect 26792 1853 26801 1887
rect 26801 1853 26835 1887
rect 26835 1853 26844 1887
rect 26792 1844 26844 1853
rect 27344 1887 27396 1896
rect 27344 1853 27353 1887
rect 27353 1853 27387 1887
rect 27387 1853 27396 1887
rect 27344 1844 27396 1853
rect 28448 1844 28500 1896
rect 31944 1844 31996 1896
rect 42340 1844 42392 1896
rect 44180 1844 44232 1896
rect 46940 1844 46992 1896
rect 12348 1776 12400 1828
rect 25504 1776 25556 1828
rect 13912 1708 13964 1760
rect 14648 1708 14700 1760
rect 17592 1708 17644 1760
rect 19248 1708 19300 1760
rect 22192 1708 22244 1760
rect 22652 1708 22704 1760
rect 25688 1708 25740 1760
rect 39948 1776 40000 1828
rect 43996 1776 44048 1828
rect 28632 1751 28684 1760
rect 28632 1717 28641 1751
rect 28641 1717 28675 1751
rect 28675 1717 28684 1751
rect 28632 1708 28684 1717
rect 29552 1751 29604 1760
rect 29552 1717 29561 1751
rect 29561 1717 29595 1751
rect 29595 1717 29604 1751
rect 29552 1708 29604 1717
rect 30012 1708 30064 1760
rect 43536 1708 43588 1760
rect 12348 1640 12400 1692
rect 13360 1640 13412 1692
rect 14280 1640 14332 1692
rect 14740 1640 14792 1692
rect 24492 1640 24544 1692
rect 31116 1683 31168 1692
rect 31116 1649 31125 1683
rect 31125 1649 31159 1683
rect 31159 1649 31168 1683
rect 31116 1640 31168 1649
rect 31300 1683 31352 1692
rect 31300 1649 31309 1683
rect 31309 1649 31343 1683
rect 31343 1649 31352 1683
rect 31300 1640 31352 1649
rect 31576 1683 31628 1692
rect 31576 1649 31585 1683
rect 31585 1649 31619 1683
rect 31619 1649 31628 1683
rect 31576 1640 31628 1649
rect 34244 1640 34296 1692
rect 43720 1640 43772 1692
rect 28356 1572 28408 1624
rect 8852 1504 8904 1556
rect 9312 1504 9364 1556
rect 13544 1504 13596 1556
rect 13728 1504 13780 1556
rect 29460 1547 29512 1556
rect 29460 1513 29469 1547
rect 29469 1513 29503 1547
rect 29503 1513 29512 1547
rect 29460 1504 29512 1513
rect 30288 1547 30340 1556
rect 30288 1513 30297 1547
rect 30297 1513 30331 1547
rect 30331 1513 30340 1547
rect 30288 1504 30340 1513
rect 30564 1547 30616 1556
rect 30564 1513 30573 1547
rect 30573 1513 30607 1547
rect 30607 1513 30616 1547
rect 30564 1504 30616 1513
rect 30840 1547 30892 1556
rect 30840 1513 30849 1547
rect 30849 1513 30883 1547
rect 30883 1513 30892 1547
rect 30840 1504 30892 1513
rect 31392 1504 31444 1556
rect 4344 1436 4396 1488
rect 4988 1436 5040 1488
rect 14740 1436 14792 1488
rect 15752 1436 15804 1488
rect 22468 1479 22520 1488
rect 22468 1445 22477 1479
rect 22477 1445 22511 1479
rect 22511 1445 22520 1479
rect 22468 1436 22520 1445
rect 24952 1436 25004 1488
rect 25228 1436 25280 1488
rect 27068 1436 27120 1488
rect 4252 1368 4304 1420
rect 4804 1368 4856 1420
rect 8392 1368 8444 1420
rect 8760 1368 8812 1420
rect 10508 1368 10560 1420
rect 16120 1368 16172 1420
rect 16580 1368 16632 1420
rect 17040 1368 17092 1420
rect 18236 1368 18288 1420
rect 19156 1368 19208 1420
rect 19892 1368 19944 1420
rect 20536 1368 20588 1420
rect 25688 1368 25740 1420
rect 29736 1368 29788 1420
rect 31668 1368 31720 1420
rect 32772 1368 32824 1420
rect 38108 1368 38160 1420
rect 38476 1368 38528 1420
rect 40040 1368 40092 1420
rect 41144 1368 41196 1420
rect 44456 1368 44508 1420
rect 48228 1368 48280 1420
rect 49700 1368 49752 1420
rect 50160 1368 50212 1420
rect 55220 1368 55272 1420
rect 55588 1368 55640 1420
rect 15016 1300 15068 1352
rect 15660 1300 15712 1352
rect 24952 1300 25004 1352
rect 30472 1343 30524 1352
rect 30472 1309 30481 1343
rect 30481 1309 30515 1343
rect 30515 1309 30524 1343
rect 30472 1300 30524 1309
rect 30748 1343 30800 1352
rect 30748 1309 30757 1343
rect 30757 1309 30791 1343
rect 30791 1309 30800 1343
rect 30748 1300 30800 1309
rect 32588 1300 32640 1352
rect 32956 1300 33008 1352
rect 58992 1300 59044 1352
rect 59176 1300 59228 1352
rect 4804 1232 4856 1284
rect 5172 1232 5224 1284
rect 33876 1232 33928 1284
rect 40592 1232 40644 1284
rect 40776 1232 40828 1284
rect 50160 1232 50212 1284
rect 50804 1232 50856 1284
rect 11428 1164 11480 1216
rect 12256 1164 12308 1216
rect 15660 1164 15712 1216
rect 16488 1164 16540 1216
rect 44640 1164 44692 1216
rect 45376 1164 45428 1216
rect 48320 1164 48372 1216
rect 52184 1164 52236 1216
rect 11060 1096 11112 1148
rect 12808 1096 12860 1148
rect 36084 1096 36136 1148
rect 33968 960 34020 1012
rect 61476 1368 61528 1420
rect 61936 1368 61988 1420
rect 63408 1368 63460 1420
rect 66812 1368 66864 1420
rect 67272 1368 67324 1420
rect 64420 1232 64472 1284
rect 64696 1232 64748 1284
rect 39764 1071 39816 1080
rect 39764 1037 39773 1071
rect 39773 1037 39807 1071
rect 39807 1037 39816 1071
rect 39764 1028 39816 1037
rect 59820 1028 59872 1080
rect 48688 960 48740 1012
rect 48964 960 49016 1012
rect 36084 892 36136 944
rect 53932 892 53984 944
rect 55036 892 55088 944
<< metal2 >>
rect 938 69200 994 70000
rect 2870 69200 2926 70000
rect 4802 69200 4858 70000
rect 6734 69200 6790 70000
rect 8666 69200 8722 70000
rect 10598 69200 10654 70000
rect 12530 69200 12586 70000
rect 14462 69200 14518 70000
rect 16486 69200 16542 70000
rect 18418 69200 18474 70000
rect 20350 69200 20406 70000
rect 22282 69200 22338 70000
rect 24214 69200 24270 70000
rect 26146 69200 26202 70000
rect 28078 69200 28134 70000
rect 30102 69200 30158 70000
rect 32034 69200 32090 70000
rect 33966 69200 34022 70000
rect 35898 69200 35954 70000
rect 37830 69200 37886 70000
rect 39762 69200 39818 70000
rect 41694 69200 41750 70000
rect 43718 69200 43774 70000
rect 45650 69200 45706 70000
rect 47582 69200 47638 70000
rect 49514 69200 49570 70000
rect 51446 69200 51502 70000
rect 53378 69200 53434 70000
rect 55310 69200 55366 70000
rect 57334 69200 57390 70000
rect 59266 69200 59322 70000
rect 61198 69200 61254 70000
rect 63130 69200 63186 70000
rect 65062 69200 65118 70000
rect 66994 69200 67050 70000
rect 67362 69320 67418 69329
rect 67362 69255 67418 69264
rect 952 67318 980 69200
rect 2778 67960 2834 67969
rect 2778 67895 2834 67904
rect 940 67312 992 67318
rect 940 67254 992 67260
rect 1768 66768 1820 66774
rect 1766 66736 1768 66745
rect 1820 66736 1822 66745
rect 2792 66706 2820 67895
rect 2884 67318 2912 69200
rect 4220 67484 4516 67504
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4298 67430 4300 67482
rect 4362 67430 4374 67482
rect 4436 67430 4438 67482
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4220 67408 4516 67428
rect 2872 67312 2924 67318
rect 2872 67254 2924 67260
rect 4816 67182 4844 69200
rect 8680 67318 8708 69200
rect 10612 67318 10640 69200
rect 8668 67312 8720 67318
rect 8668 67254 8720 67260
rect 10600 67312 10652 67318
rect 10600 67254 10652 67260
rect 12544 67182 12572 69200
rect 14220 67484 14516 67504
rect 14276 67482 14300 67484
rect 14356 67482 14380 67484
rect 14436 67482 14460 67484
rect 14298 67430 14300 67482
rect 14362 67430 14374 67482
rect 14436 67430 14438 67482
rect 14276 67428 14300 67430
rect 14356 67428 14380 67430
rect 14436 67428 14460 67430
rect 14220 67408 14516 67428
rect 16500 67386 16528 69200
rect 16488 67380 16540 67386
rect 16488 67322 16540 67328
rect 18432 67318 18460 69200
rect 18420 67312 18472 67318
rect 18420 67254 18472 67260
rect 20364 67182 20392 69200
rect 24228 67674 24256 69200
rect 24136 67646 24256 67674
rect 24136 67318 24164 67646
rect 24220 67484 24516 67504
rect 24276 67482 24300 67484
rect 24356 67482 24380 67484
rect 24436 67482 24460 67484
rect 24298 67430 24300 67482
rect 24362 67430 24374 67482
rect 24436 67430 24438 67482
rect 24276 67428 24300 67430
rect 24356 67428 24380 67430
rect 24436 67428 24460 67430
rect 24220 67408 24516 67428
rect 26160 67318 26188 69200
rect 24124 67312 24176 67318
rect 24124 67254 24176 67260
rect 26148 67312 26200 67318
rect 26148 67254 26200 67260
rect 28092 67182 28120 69200
rect 32048 67318 32076 69200
rect 33980 67318 34008 69200
rect 34220 67484 34516 67504
rect 34276 67482 34300 67484
rect 34356 67482 34380 67484
rect 34436 67482 34460 67484
rect 34298 67430 34300 67482
rect 34362 67430 34374 67482
rect 34436 67430 34438 67482
rect 34276 67428 34300 67430
rect 34356 67428 34380 67430
rect 34436 67428 34460 67430
rect 34220 67408 34516 67428
rect 32036 67312 32088 67318
rect 32036 67254 32088 67260
rect 33968 67312 34020 67318
rect 33968 67254 34020 67260
rect 35912 67182 35940 69200
rect 39776 67318 39804 69200
rect 41708 67318 41736 69200
rect 39764 67312 39816 67318
rect 39764 67254 39816 67260
rect 41696 67312 41748 67318
rect 41696 67254 41748 67260
rect 43732 67182 43760 69200
rect 44220 67484 44516 67504
rect 44276 67482 44300 67484
rect 44356 67482 44380 67484
rect 44436 67482 44460 67484
rect 44298 67430 44300 67482
rect 44362 67430 44374 67482
rect 44436 67430 44438 67482
rect 44276 67428 44300 67430
rect 44356 67428 44380 67430
rect 44436 67428 44460 67430
rect 44220 67408 44516 67428
rect 47596 67318 47624 69200
rect 49528 67318 49556 69200
rect 47584 67312 47636 67318
rect 47584 67254 47636 67260
rect 49516 67312 49568 67318
rect 49516 67254 49568 67260
rect 51460 67182 51488 69200
rect 54220 67484 54516 67504
rect 54276 67482 54300 67484
rect 54356 67482 54380 67484
rect 54436 67482 54460 67484
rect 54298 67430 54300 67482
rect 54362 67430 54374 67482
rect 54436 67430 54438 67482
rect 54276 67428 54300 67430
rect 54356 67428 54380 67430
rect 54436 67428 54460 67430
rect 54220 67408 54516 67428
rect 55324 67318 55352 69200
rect 57348 67318 57376 69200
rect 59280 67634 59308 69200
rect 59280 67606 59400 67634
rect 55312 67312 55364 67318
rect 55312 67254 55364 67260
rect 57336 67312 57388 67318
rect 57336 67254 57388 67260
rect 59372 67182 59400 67606
rect 63144 67318 63172 69200
rect 64220 67484 64516 67504
rect 64276 67482 64300 67484
rect 64356 67482 64380 67484
rect 64436 67482 64460 67484
rect 64298 67430 64300 67482
rect 64362 67430 64374 67482
rect 64436 67430 64438 67482
rect 64276 67428 64300 67430
rect 64356 67428 64380 67430
rect 64436 67428 64460 67430
rect 64220 67408 64516 67428
rect 65076 67318 65104 69200
rect 63132 67312 63184 67318
rect 63132 67254 63184 67260
rect 65064 67312 65116 67318
rect 65064 67254 65116 67260
rect 67008 67182 67036 69200
rect 67376 67318 67404 69255
rect 68926 69200 68982 70000
rect 67546 67960 67602 67969
rect 67546 67895 67602 67904
rect 67364 67312 67416 67318
rect 67364 67254 67416 67260
rect 4804 67176 4856 67182
rect 4804 67118 4856 67124
rect 12532 67176 12584 67182
rect 12532 67118 12584 67124
rect 20352 67176 20404 67182
rect 20352 67118 20404 67124
rect 26976 67176 27028 67182
rect 26976 67118 27028 67124
rect 28080 67176 28132 67182
rect 28080 67118 28132 67124
rect 35900 67176 35952 67182
rect 35900 67118 35952 67124
rect 43720 67176 43772 67182
rect 43720 67118 43772 67124
rect 51448 67176 51500 67182
rect 51448 67118 51500 67124
rect 59360 67176 59412 67182
rect 59360 67118 59412 67124
rect 64788 67176 64840 67182
rect 64788 67118 64840 67124
rect 66996 67176 67048 67182
rect 66996 67118 67048 67124
rect 3976 67108 4028 67114
rect 3976 67050 4028 67056
rect 11060 67108 11112 67114
rect 11060 67050 11112 67056
rect 16580 67108 16632 67114
rect 16580 67050 16632 67056
rect 3884 67040 3936 67046
rect 3884 66982 3936 66988
rect 1766 66671 1822 66680
rect 1952 66700 2004 66706
rect 1952 66642 2004 66648
rect 2780 66700 2832 66706
rect 2780 66642 2832 66648
rect 1964 66162 1992 66642
rect 3896 66638 3924 66982
rect 3884 66632 3936 66638
rect 3884 66574 3936 66580
rect 3988 66502 4016 67050
rect 9220 66940 9516 66960
rect 9276 66938 9300 66940
rect 9356 66938 9380 66940
rect 9436 66938 9460 66940
rect 9298 66886 9300 66938
rect 9362 66886 9374 66938
rect 9436 66886 9438 66938
rect 9276 66884 9300 66886
rect 9356 66884 9380 66886
rect 9436 66884 9460 66886
rect 9220 66864 9516 66884
rect 10140 66700 10192 66706
rect 10140 66642 10192 66648
rect 3976 66496 4028 66502
rect 3976 66438 4028 66444
rect 1952 66156 2004 66162
rect 1952 66098 2004 66104
rect 1860 65408 1912 65414
rect 1858 65376 1860 65385
rect 2688 65408 2740 65414
rect 1912 65376 1914 65385
rect 2688 65350 2740 65356
rect 1858 65311 1914 65320
rect 2228 64320 2280 64326
rect 2228 64262 2280 64268
rect 2240 64122 2268 64262
rect 2228 64116 2280 64122
rect 2228 64058 2280 64064
rect 2044 62960 2096 62966
rect 2044 62902 2096 62908
rect 1584 62824 1636 62830
rect 1582 62792 1584 62801
rect 1636 62792 1638 62801
rect 1582 62727 1638 62736
rect 1860 61600 1912 61606
rect 1858 61568 1860 61577
rect 1912 61568 1914 61577
rect 1858 61503 1914 61512
rect 1766 60208 1822 60217
rect 1766 60143 1768 60152
rect 1820 60143 1822 60152
rect 1860 60172 1912 60178
rect 1768 60114 1820 60120
rect 1860 60114 1912 60120
rect 1582 57624 1638 57633
rect 1582 57559 1638 57568
rect 1596 57390 1624 57559
rect 1584 57384 1636 57390
rect 1584 57326 1636 57332
rect 1766 56400 1822 56409
rect 1766 56335 1768 56344
rect 1820 56335 1822 56344
rect 1768 56306 1820 56312
rect 1872 55214 1900 60114
rect 1872 55186 1992 55214
rect 1860 55072 1912 55078
rect 1858 55040 1860 55049
rect 1912 55040 1914 55049
rect 1858 54975 1914 54984
rect 1584 52556 1636 52562
rect 1584 52498 1636 52504
rect 1596 52465 1624 52498
rect 1582 52456 1638 52465
rect 1582 52391 1638 52400
rect 1858 51096 1914 51105
rect 1858 51031 1860 51040
rect 1912 51031 1914 51040
rect 1860 51002 1912 51008
rect 1766 49872 1822 49881
rect 1766 49807 1768 49816
rect 1820 49807 1822 49816
rect 1768 49778 1820 49784
rect 1858 47288 1914 47297
rect 1858 47223 1914 47232
rect 1872 47190 1900 47223
rect 1860 47184 1912 47190
rect 1860 47126 1912 47132
rect 1872 46714 1900 47126
rect 1860 46708 1912 46714
rect 1860 46650 1912 46656
rect 1768 45960 1820 45966
rect 1766 45928 1768 45937
rect 1820 45928 1822 45937
rect 1766 45863 1822 45872
rect 1860 44736 1912 44742
rect 1858 44704 1860 44713
rect 1912 44704 1914 44713
rect 1858 44639 1914 44648
rect 1584 42152 1636 42158
rect 1582 42120 1584 42129
rect 1636 42120 1638 42129
rect 1582 42055 1638 42064
rect 1858 40760 1914 40769
rect 1858 40695 1860 40704
rect 1912 40695 1914 40704
rect 1860 40666 1912 40672
rect 1766 39536 1822 39545
rect 1766 39471 1768 39480
rect 1820 39471 1822 39480
rect 1768 39442 1820 39448
rect 1582 36952 1638 36961
rect 1582 36887 1638 36896
rect 1596 36718 1624 36887
rect 1584 36712 1636 36718
rect 1584 36654 1636 36660
rect 1768 35624 1820 35630
rect 1766 35592 1768 35601
rect 1820 35592 1822 35601
rect 1766 35527 1822 35536
rect 1308 35148 1360 35154
rect 1308 35090 1360 35096
rect 1320 6914 1348 35090
rect 1858 34232 1914 34241
rect 1858 34167 1860 34176
rect 1912 34167 1914 34176
rect 1860 34138 1912 34144
rect 1584 31884 1636 31890
rect 1584 31826 1636 31832
rect 1596 31657 1624 31826
rect 1582 31648 1638 31657
rect 1582 31583 1638 31592
rect 1766 30424 1822 30433
rect 1766 30359 1822 30368
rect 1780 30326 1808 30359
rect 1768 30320 1820 30326
rect 1768 30262 1820 30268
rect 1768 29096 1820 29102
rect 1766 29064 1768 29073
rect 1820 29064 1822 29073
rect 1766 28999 1822 29008
rect 1584 26920 1636 26926
rect 1584 26862 1636 26868
rect 1596 26489 1624 26862
rect 1582 26480 1638 26489
rect 1582 26415 1638 26424
rect 1964 26234 1992 55186
rect 2056 29102 2084 62902
rect 2320 61600 2372 61606
rect 2320 61542 2372 61548
rect 2136 60104 2188 60110
rect 2136 60046 2188 60052
rect 2148 45014 2176 60046
rect 2136 45008 2188 45014
rect 2136 44950 2188 44956
rect 2136 34060 2188 34066
rect 2136 34002 2188 34008
rect 2148 33862 2176 34002
rect 2136 33856 2188 33862
rect 2136 33798 2188 33804
rect 2044 29096 2096 29102
rect 2044 29038 2096 29044
rect 1872 26206 1992 26234
rect 1766 25256 1822 25265
rect 1766 25191 1768 25200
rect 1820 25191 1822 25200
rect 1768 25162 1820 25168
rect 1872 24206 1900 26206
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1858 23896 1914 23905
rect 1858 23831 1860 23840
rect 1912 23831 1914 23840
rect 1860 23802 1912 23808
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 21321 1440 21422
rect 1398 21312 1454 21321
rect 1398 21247 1454 21256
rect 1412 21146 1440 21247
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 1858 20088 1914 20097
rect 1858 20023 1860 20032
rect 1912 20023 1914 20032
rect 1860 19994 1912 20000
rect 1766 18728 1822 18737
rect 1766 18663 1768 18672
rect 1820 18663 1822 18672
rect 1768 18634 1820 18640
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1596 16046 1624 16079
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 2148 15570 2176 33798
rect 2228 30116 2280 30122
rect 2228 30058 2280 30064
rect 2240 29510 2268 30058
rect 2228 29504 2280 29510
rect 2228 29446 2280 29452
rect 2240 29306 2268 29446
rect 2228 29300 2280 29306
rect 2228 29242 2280 29248
rect 2332 28082 2360 61542
rect 2596 59968 2648 59974
rect 2596 59910 2648 59916
rect 2504 56160 2556 56166
rect 2504 56102 2556 56108
rect 2412 54324 2464 54330
rect 2412 54266 2464 54272
rect 2424 46170 2452 54266
rect 2516 51270 2544 56102
rect 2504 51264 2556 51270
rect 2504 51206 2556 51212
rect 2412 46164 2464 46170
rect 2412 46106 2464 46112
rect 2412 40588 2464 40594
rect 2412 40530 2464 40536
rect 2424 40390 2452 40530
rect 2412 40384 2464 40390
rect 2412 40326 2464 40332
rect 2424 35894 2452 40326
rect 2608 39642 2636 59910
rect 2700 58546 2728 65350
rect 3988 62898 4016 66438
rect 4220 66396 4516 66416
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4298 66342 4300 66394
rect 4362 66342 4374 66394
rect 4436 66342 4438 66394
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4220 66320 4516 66340
rect 4252 66088 4304 66094
rect 4252 66030 4304 66036
rect 4264 65550 4292 66030
rect 9220 65852 9516 65872
rect 9276 65850 9300 65852
rect 9356 65850 9380 65852
rect 9436 65850 9460 65852
rect 9298 65798 9300 65850
rect 9362 65798 9374 65850
rect 9436 65798 9438 65850
rect 9276 65796 9300 65798
rect 9356 65796 9380 65798
rect 9436 65796 9460 65798
rect 9220 65776 9516 65796
rect 4620 65612 4672 65618
rect 4620 65554 4672 65560
rect 4252 65544 4304 65550
rect 4252 65486 4304 65492
rect 4220 65308 4516 65328
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4298 65254 4300 65306
rect 4362 65254 4374 65306
rect 4436 65254 4438 65306
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4220 65232 4516 65252
rect 4220 64220 4516 64240
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4298 64166 4300 64218
rect 4362 64166 4374 64218
rect 4436 64166 4438 64218
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4220 64144 4516 64164
rect 4220 63132 4516 63152
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4298 63078 4300 63130
rect 4362 63078 4374 63130
rect 4436 63078 4438 63130
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4220 63056 4516 63076
rect 3976 62892 4028 62898
rect 3976 62834 4028 62840
rect 4220 62044 4516 62064
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4298 61990 4300 62042
rect 4362 61990 4374 62042
rect 4436 61990 4438 62042
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4220 61968 4516 61988
rect 4220 60956 4516 60976
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4298 60902 4300 60954
rect 4362 60902 4374 60954
rect 4436 60902 4438 60954
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4220 60880 4516 60900
rect 4220 59868 4516 59888
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4298 59814 4300 59866
rect 4362 59814 4374 59866
rect 4436 59814 4438 59866
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4220 59792 4516 59812
rect 4220 58780 4516 58800
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4298 58726 4300 58778
rect 4362 58726 4374 58778
rect 4436 58726 4438 58778
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4220 58704 4516 58724
rect 3884 58608 3936 58614
rect 3884 58550 3936 58556
rect 2688 58540 2740 58546
rect 2688 58482 2740 58488
rect 2688 55684 2740 55690
rect 2688 55626 2740 55632
rect 2700 55282 2728 55626
rect 2688 55276 2740 55282
rect 2688 55218 2740 55224
rect 2688 53236 2740 53242
rect 2688 53178 2740 53184
rect 2700 51066 2728 53178
rect 2688 51060 2740 51066
rect 2688 51002 2740 51008
rect 3148 50176 3200 50182
rect 3148 50118 3200 50124
rect 2596 39636 2648 39642
rect 2596 39578 2648 39584
rect 2688 39364 2740 39370
rect 2688 39306 2740 39312
rect 2424 35866 2636 35894
rect 2504 35216 2556 35222
rect 2504 35158 2556 35164
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2516 27826 2544 35158
rect 2240 27798 2544 27826
rect 2240 18970 2268 27798
rect 2608 26234 2636 35866
rect 2700 30326 2728 39306
rect 2872 36032 2924 36038
rect 2872 35974 2924 35980
rect 2688 30320 2740 30326
rect 2688 30262 2740 30268
rect 2424 26206 2636 26234
rect 2424 25974 2452 26206
rect 2412 25968 2464 25974
rect 2412 25910 2464 25916
rect 2596 25152 2648 25158
rect 2596 25094 2648 25100
rect 2608 24954 2636 25094
rect 2596 24948 2648 24954
rect 2596 24890 2648 24896
rect 2320 23588 2372 23594
rect 2320 23530 2372 23536
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 1860 14816 1912 14822
rect 1858 14784 1860 14793
rect 1912 14784 1914 14793
rect 1858 14719 1914 14728
rect 1858 13560 1914 13569
rect 1858 13495 1860 13504
rect 1912 13495 1914 13504
rect 1860 13466 1912 13472
rect 2332 13462 2360 23530
rect 2884 18698 2912 35974
rect 2964 29708 3016 29714
rect 2964 29650 3016 29656
rect 2872 18692 2924 18698
rect 2872 18634 2924 18640
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2332 12986 2360 13398
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1596 10985 1624 11154
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 2424 10266 2452 13398
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 1768 9648 1820 9654
rect 1766 9616 1768 9625
rect 1820 9616 1822 9625
rect 1766 9551 1822 9560
rect 2424 9518 2452 10202
rect 2608 9654 2636 14758
rect 2976 12434 3004 29650
rect 3160 23866 3188 50118
rect 3700 43308 3752 43314
rect 3700 43250 3752 43256
rect 3712 43110 3740 43250
rect 3700 43104 3752 43110
rect 3700 43046 3752 43052
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3712 22778 3740 43046
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 2792 12406 3004 12434
rect 2686 11112 2742 11121
rect 2686 11047 2742 11056
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1136 6886 1348 6914
rect 388 4140 440 4146
rect 388 4082 440 4088
rect 20 3528 72 3534
rect 20 3470 72 3476
rect 32 800 60 3470
rect 112 2848 164 2854
rect 112 2790 164 2796
rect 124 800 152 2790
rect 296 2372 348 2378
rect 296 2314 348 2320
rect 308 800 336 2314
rect 400 800 428 4082
rect 848 4072 900 4078
rect 848 4014 900 4020
rect 572 4004 624 4010
rect 572 3946 624 3952
rect 584 800 612 3946
rect 664 3460 716 3466
rect 664 3402 716 3408
rect 676 800 704 3402
rect 860 800 888 4014
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 952 800 980 3878
rect 1136 3534 1164 6886
rect 1412 6254 1440 8774
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 4026 1440 6190
rect 1504 5166 1532 7686
rect 1582 7032 1638 7041
rect 1582 6967 1638 6976
rect 1596 6866 1624 6967
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1688 6254 1716 8774
rect 1768 8424 1820 8430
rect 1766 8392 1768 8401
rect 1820 8392 1822 8401
rect 1766 8327 1822 8336
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1504 4146 1532 5102
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1596 4026 1624 5102
rect 1228 3998 1440 4026
rect 1504 3998 1624 4026
rect 1688 4010 1716 6190
rect 1768 5840 1820 5846
rect 1766 5808 1768 5817
rect 1820 5808 1822 5817
rect 1766 5743 1822 5752
rect 1872 4570 1900 7278
rect 1964 5166 1992 7686
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1780 4542 1900 4570
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1676 4004 1728 4010
rect 1124 3528 1176 3534
rect 1124 3470 1176 3476
rect 1124 2576 1176 2582
rect 1124 2518 1176 2524
rect 1136 800 1164 2518
rect 1228 800 1256 3998
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1412 800 1440 3470
rect 1504 800 1532 3998
rect 1676 3946 1728 3952
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1596 3233 1624 3538
rect 1582 3224 1638 3233
rect 1582 3159 1638 3168
rect 1688 3074 1716 3674
rect 1780 3466 1808 4542
rect 1860 4480 1912 4486
rect 1858 4448 1860 4457
rect 1912 4448 1914 4457
rect 1858 4383 1914 4392
rect 1964 3942 1992 4558
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 2056 3754 2084 5714
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1872 3726 2084 3754
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1872 3346 1900 3726
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1596 3046 1716 3074
rect 1780 3318 1900 3346
rect 1596 2854 1624 3046
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2514 1624 2790
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1688 800 1716 2926
rect 1780 1714 1808 3318
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 1873 1900 2790
rect 1858 1864 1914 1873
rect 1858 1799 1914 1808
rect 1780 1686 1900 1714
rect 1872 800 1900 1686
rect 1964 800 1992 3402
rect 2148 800 2176 4082
rect 2240 4078 2268 7142
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3618 2268 3878
rect 2332 3738 2360 5510
rect 2424 4078 2452 8842
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 7342 2544 8774
rect 2700 8650 2728 11047
rect 2792 9926 2820 12406
rect 3896 9926 3924 58550
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 2608 8622 2728 8650
rect 2608 8430 2636 8622
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2516 4690 2544 6666
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2240 3590 2360 3618
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2240 800 2268 2994
rect 2332 2922 2360 3590
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 2424 800 2452 3878
rect 2516 800 2544 4014
rect 2608 3602 2636 6598
rect 2700 5778 2728 8502
rect 2792 5846 2820 9862
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4026 2820 5102
rect 2700 3998 2820 4026
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2700 800 2728 3998
rect 2884 3194 2912 8230
rect 2976 6254 3004 8774
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2792 800 2820 3062
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 18 0 74 800
rect 110 0 166 800
rect 294 0 350 800
rect 386 0 442 800
rect 570 0 626 800
rect 662 0 718 800
rect 846 0 902 800
rect 938 0 994 800
rect 1122 0 1178 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 1950 0 2006 800
rect 2134 0 2190 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2884 649 2912 2790
rect 2976 800 3004 6190
rect 3068 5710 3096 8298
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3160 4078 3188 6598
rect 3252 4690 3280 7686
rect 3344 5778 3372 8298
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3332 5772 3384 5778
rect 3384 5732 3464 5760
rect 3332 5714 3384 5720
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3252 4146 3280 4626
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3148 4072 3200 4078
rect 3344 4026 3372 5102
rect 3148 4014 3200 4020
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 3252 3998 3372 4026
rect 3068 800 3096 3946
rect 3252 800 3280 3998
rect 3436 3942 3464 5732
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3344 800 3372 3130
rect 3528 800 3556 4014
rect 3620 3602 3648 6054
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3712 2990 3740 9862
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3976 8832 4028 8838
rect 4172 8820 4200 9454
rect 3976 8774 4028 8780
rect 4080 8792 4200 8820
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 4078 3832 6598
rect 3896 5166 3924 7686
rect 3988 5273 4016 8774
rect 4080 8548 4108 8792
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4632 8634 4660 65554
rect 9220 64764 9516 64784
rect 9276 64762 9300 64764
rect 9356 64762 9380 64764
rect 9436 64762 9460 64764
rect 9298 64710 9300 64762
rect 9362 64710 9374 64762
rect 9436 64710 9438 64762
rect 9276 64708 9300 64710
rect 9356 64708 9380 64710
rect 9436 64708 9460 64710
rect 9220 64688 9516 64708
rect 6736 64320 6788 64326
rect 6736 64262 6788 64268
rect 4712 57996 4764 58002
rect 4712 57938 4764 57944
rect 4724 57798 4752 57938
rect 6368 57928 6420 57934
rect 6368 57870 6420 57876
rect 4712 57792 4764 57798
rect 4712 57734 4764 57740
rect 4724 14890 4752 57734
rect 6380 57254 6408 57870
rect 6368 57248 6420 57254
rect 6368 57190 6420 57196
rect 5724 38004 5776 38010
rect 5724 37946 5776 37952
rect 4896 37800 4948 37806
rect 4896 37742 4948 37748
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4816 12434 4844 29038
rect 4724 12406 4844 12434
rect 4724 9926 4752 12406
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4080 8520 4200 8548
rect 4172 7834 4200 8520
rect 4080 7806 4200 7834
rect 4080 7546 4108 7806
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4632 7410 4660 8570
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3974 5264 4030 5273
rect 4080 5234 4108 7142
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 3974 5199 4030 5208
rect 4068 5228 4120 5234
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3988 4758 4016 5199
rect 4068 5170 4120 5176
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 4172 4570 4200 5102
rect 4632 4690 4660 6054
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4080 4542 4200 4570
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3896 3670 3924 4422
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 800 3740 2790
rect 3804 800 3832 3402
rect 3988 800 4016 4082
rect 4080 2922 4108 4542
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4632 4146 4660 4626
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4172 2774 4200 2994
rect 4080 2746 4200 2774
rect 4080 800 4108 2746
rect 4632 2530 4660 3946
rect 4724 3738 4752 9862
rect 4816 9518 4844 10610
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4908 8294 4936 37742
rect 5356 35692 5408 35698
rect 5356 35634 5408 35640
rect 4988 29028 5040 29034
rect 4988 28970 5040 28976
rect 5000 9382 5028 28970
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 9654 5120 19654
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4816 5302 4844 7686
rect 4908 5778 4936 7686
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6322 5120 6598
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4816 3584 4844 5102
rect 4724 3556 4844 3584
rect 4724 3058 4752 3556
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4632 2502 4752 2530
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4526 2000 4582 2009
rect 4526 1935 4582 1944
rect 4344 1488 4396 1494
rect 4344 1430 4396 1436
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 4264 800 4292 1362
rect 4356 800 4384 1430
rect 4540 800 4568 1935
rect 4724 1306 4752 2502
rect 4816 1426 4844 3402
rect 4804 1420 4856 1426
rect 4804 1362 4856 1368
rect 4632 1278 4752 1306
rect 4804 1284 4856 1290
rect 4632 800 4660 1278
rect 4804 1226 4856 1232
rect 4816 800 4844 1226
rect 4908 800 4936 5714
rect 5000 4690 5028 6054
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5000 1494 5028 4626
rect 5092 4146 5120 6122
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5184 4078 5212 9862
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4988 1488 5040 1494
rect 4988 1430 5040 1436
rect 5092 800 5120 3334
rect 5184 1290 5212 3674
rect 5276 2922 5304 9318
rect 5368 8838 5396 35634
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5460 9926 5488 23802
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5644 9518 5672 14486
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5262 2816 5318 2825
rect 5262 2751 5318 2760
rect 5172 1284 5224 1290
rect 5172 1226 5224 1232
rect 5276 898 5304 2751
rect 5368 2582 5396 8774
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 5302 5488 7142
rect 5552 5778 5580 7686
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5448 5160 5500 5166
rect 5446 5128 5448 5137
rect 5500 5128 5502 5137
rect 5446 5063 5502 5072
rect 5552 4128 5580 5714
rect 5460 4100 5580 4128
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 5460 898 5488 4100
rect 5644 3670 5672 9318
rect 5736 8362 5764 37946
rect 6092 34944 6144 34950
rect 6092 34886 6144 34892
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5724 7200 5776 7206
rect 5722 7168 5724 7177
rect 5776 7168 5778 7177
rect 5722 7103 5778 7112
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 4690 5764 6054
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5736 3738 5764 4626
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5184 870 5304 898
rect 5368 870 5488 898
rect 5184 800 5212 870
rect 5368 800 5396 870
rect 5552 800 5580 2926
rect 5644 800 5672 3470
rect 5828 3058 5856 9454
rect 6104 8838 6132 34886
rect 6748 16574 6776 64262
rect 9220 63676 9516 63696
rect 9276 63674 9300 63676
rect 9356 63674 9380 63676
rect 9436 63674 9460 63676
rect 9298 63622 9300 63674
rect 9362 63622 9374 63674
rect 9436 63622 9438 63674
rect 9276 63620 9300 63622
rect 9356 63620 9380 63622
rect 9436 63620 9460 63622
rect 9220 63600 9516 63620
rect 9772 62824 9824 62830
rect 9772 62766 9824 62772
rect 9220 62588 9516 62608
rect 9276 62586 9300 62588
rect 9356 62586 9380 62588
rect 9436 62586 9460 62588
rect 9298 62534 9300 62586
rect 9362 62534 9374 62586
rect 9436 62534 9438 62586
rect 9276 62532 9300 62534
rect 9356 62532 9380 62534
rect 9436 62532 9460 62534
rect 9220 62512 9516 62532
rect 9784 62490 9812 62766
rect 9772 62484 9824 62490
rect 9772 62426 9824 62432
rect 9220 61500 9516 61520
rect 9276 61498 9300 61500
rect 9356 61498 9380 61500
rect 9436 61498 9460 61500
rect 9298 61446 9300 61498
rect 9362 61446 9374 61498
rect 9436 61446 9438 61498
rect 9276 61444 9300 61446
rect 9356 61444 9380 61446
rect 9436 61444 9460 61446
rect 9220 61424 9516 61444
rect 9220 60412 9516 60432
rect 9276 60410 9300 60412
rect 9356 60410 9380 60412
rect 9436 60410 9460 60412
rect 9298 60358 9300 60410
rect 9362 60358 9374 60410
rect 9436 60358 9438 60410
rect 9276 60356 9300 60358
rect 9356 60356 9380 60358
rect 9436 60356 9460 60358
rect 9220 60336 9516 60356
rect 9220 59324 9516 59344
rect 9276 59322 9300 59324
rect 9356 59322 9380 59324
rect 9436 59322 9460 59324
rect 9298 59270 9300 59322
rect 9362 59270 9374 59322
rect 9436 59270 9438 59322
rect 9276 59268 9300 59270
rect 9356 59268 9380 59270
rect 9436 59268 9460 59270
rect 9220 59248 9516 59268
rect 8208 58676 8260 58682
rect 8208 58618 8260 58624
rect 8220 58138 8248 58618
rect 9220 58236 9516 58256
rect 9276 58234 9300 58236
rect 9356 58234 9380 58236
rect 9436 58234 9460 58236
rect 9298 58182 9300 58234
rect 9362 58182 9374 58234
rect 9436 58182 9438 58234
rect 9276 58180 9300 58182
rect 9356 58180 9380 58182
rect 9436 58180 9460 58182
rect 9220 58160 9516 58180
rect 6920 58132 6972 58138
rect 6920 58074 6972 58080
rect 8208 58132 8260 58138
rect 8208 58074 8260 58080
rect 6932 58002 6960 58074
rect 6920 57996 6972 58002
rect 6920 57938 6972 57944
rect 8208 57792 8260 57798
rect 8208 57734 8260 57740
rect 8220 57594 8248 57734
rect 8208 57588 8260 57594
rect 8208 57530 8260 57536
rect 8852 57452 8904 57458
rect 8852 57394 8904 57400
rect 6920 49768 6972 49774
rect 6920 49710 6972 49716
rect 6656 16546 6776 16574
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5828 800 5856 2790
rect 5920 2582 5948 8774
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 6012 4690 6040 6666
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6104 5166 6132 6598
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 2825 6040 4626
rect 6196 3924 6224 8298
rect 6288 8090 6316 8842
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6288 7274 6316 8026
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 4078 6316 5510
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6196 3896 6316 3924
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5998 2816 6054 2825
rect 5998 2751 6054 2760
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5920 800 5948 2246
rect 6104 800 6132 3470
rect 6196 800 6224 3674
rect 6288 2774 6316 3896
rect 6380 3670 6408 9862
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6288 2746 6408 2774
rect 6380 2514 6408 2746
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6380 800 6408 2314
rect 6472 800 6500 4014
rect 6564 2922 6592 9658
rect 6656 9382 6684 16546
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6748 9926 6776 14418
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6840 7546 6868 9454
rect 6932 8634 6960 49710
rect 7288 44804 7340 44810
rect 7288 44746 7340 44752
rect 7012 44736 7064 44742
rect 7012 44678 7064 44684
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6932 7342 6960 8570
rect 7024 7546 7052 44678
rect 7196 35624 7248 35630
rect 7196 35566 7248 35572
rect 7104 34740 7156 34746
rect 7104 34682 7156 34688
rect 7116 8838 7144 34682
rect 7208 32473 7236 35566
rect 7194 32464 7250 32473
rect 7194 32399 7250 32408
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 7208 9926 7236 27270
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6656 800 6684 5102
rect 6748 3602 6776 6054
rect 6828 4208 6880 4214
rect 6826 4176 6828 4185
rect 6880 4176 6882 4185
rect 6826 4111 6882 4120
rect 6932 4078 6960 6598
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 4826 7052 6258
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6748 800 6776 2246
rect 6932 800 6960 3402
rect 7024 2854 7052 4626
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7116 2582 7144 8774
rect 7208 2990 7236 9862
rect 7300 8906 7328 44746
rect 7840 42560 7892 42566
rect 7840 42502 7892 42508
rect 7380 29504 7432 29510
rect 7380 29446 7432 29452
rect 7392 21457 7420 29446
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7378 21448 7434 21457
rect 7378 21383 7434 21392
rect 7484 9178 7512 24074
rect 7852 9382 7880 42502
rect 8392 35012 8444 35018
rect 8392 34954 8444 34960
rect 8404 34746 8432 34954
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8484 27940 8536 27946
rect 8484 27882 8536 27888
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7944 24886 7972 25094
rect 7932 24880 7984 24886
rect 7932 24822 7984 24828
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 9382 8432 18566
rect 8496 12434 8524 27882
rect 8576 22432 8628 22438
rect 8576 22374 8628 22380
rect 8588 22234 8616 22374
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8496 12406 8616 12434
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7300 2774 7328 5102
rect 7392 4690 7420 7686
rect 7484 7342 7512 9114
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7576 5166 7604 8298
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7208 2746 7328 2774
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7208 1442 7236 2746
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7116 1414 7236 1442
rect 7116 800 7144 1414
rect 7300 1170 7328 2314
rect 7208 1142 7328 1170
rect 7208 800 7236 1142
rect 7392 800 7420 4014
rect 7484 800 7512 5034
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7576 3738 7604 4626
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7668 3602 7696 6598
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7760 5098 7788 5510
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7760 3738 7788 4762
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7852 2582 7880 9318
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7944 4690 7972 7686
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7668 800 7696 2450
rect 7944 1578 7972 4014
rect 8036 3602 8064 7142
rect 8128 5166 8156 8298
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8220 4128 8248 6598
rect 8312 5778 8340 8774
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8128 4100 8248 4128
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7760 1550 7972 1578
rect 7760 800 7788 1550
rect 8036 1442 8064 3334
rect 8128 3126 8156 4100
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8128 2990 8156 3062
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 7944 1414 8064 1442
rect 7944 800 7972 1414
rect 8128 1170 8156 2246
rect 8036 1142 8156 1170
rect 8036 800 8064 1142
rect 8220 800 8248 3946
rect 8312 800 8340 5714
rect 8404 4078 8432 7686
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8404 1426 8432 3674
rect 8496 3058 8524 10474
rect 8588 9926 8616 12406
rect 8864 10470 8892 57394
rect 9220 57148 9516 57168
rect 9276 57146 9300 57148
rect 9356 57146 9380 57148
rect 9436 57146 9460 57148
rect 9298 57094 9300 57146
rect 9362 57094 9374 57146
rect 9436 57094 9438 57146
rect 9276 57092 9300 57094
rect 9356 57092 9380 57094
rect 9436 57092 9460 57094
rect 9220 57072 9516 57092
rect 9220 56060 9516 56080
rect 9276 56058 9300 56060
rect 9356 56058 9380 56060
rect 9436 56058 9460 56060
rect 9298 56006 9300 56058
rect 9362 56006 9374 56058
rect 9436 56006 9438 56058
rect 9276 56004 9300 56006
rect 9356 56004 9380 56006
rect 9436 56004 9460 56006
rect 9220 55984 9516 56004
rect 9956 55820 10008 55826
rect 9956 55762 10008 55768
rect 9968 55350 9996 55762
rect 9956 55344 10008 55350
rect 9956 55286 10008 55292
rect 9220 54972 9516 54992
rect 9276 54970 9300 54972
rect 9356 54970 9380 54972
rect 9436 54970 9460 54972
rect 9298 54918 9300 54970
rect 9362 54918 9374 54970
rect 9436 54918 9438 54970
rect 9276 54916 9300 54918
rect 9356 54916 9380 54918
rect 9436 54916 9460 54918
rect 9220 54896 9516 54916
rect 9220 53884 9516 53904
rect 9276 53882 9300 53884
rect 9356 53882 9380 53884
rect 9436 53882 9460 53884
rect 9298 53830 9300 53882
rect 9362 53830 9374 53882
rect 9436 53830 9438 53882
rect 9276 53828 9300 53830
rect 9356 53828 9380 53830
rect 9436 53828 9460 53830
rect 9220 53808 9516 53828
rect 9220 52796 9516 52816
rect 9276 52794 9300 52796
rect 9356 52794 9380 52796
rect 9436 52794 9460 52796
rect 9298 52742 9300 52794
rect 9362 52742 9374 52794
rect 9436 52742 9438 52794
rect 9276 52740 9300 52742
rect 9356 52740 9380 52742
rect 9436 52740 9460 52742
rect 9220 52720 9516 52740
rect 9220 51708 9516 51728
rect 9276 51706 9300 51708
rect 9356 51706 9380 51708
rect 9436 51706 9460 51708
rect 9298 51654 9300 51706
rect 9362 51654 9374 51706
rect 9436 51654 9438 51706
rect 9276 51652 9300 51654
rect 9356 51652 9380 51654
rect 9436 51652 9460 51654
rect 9220 51632 9516 51652
rect 9220 50620 9516 50640
rect 9276 50618 9300 50620
rect 9356 50618 9380 50620
rect 9436 50618 9460 50620
rect 9298 50566 9300 50618
rect 9362 50566 9374 50618
rect 9436 50566 9438 50618
rect 9276 50564 9300 50566
rect 9356 50564 9380 50566
rect 9436 50564 9460 50566
rect 9220 50544 9516 50564
rect 9220 49532 9516 49552
rect 9276 49530 9300 49532
rect 9356 49530 9380 49532
rect 9436 49530 9460 49532
rect 9298 49478 9300 49530
rect 9362 49478 9374 49530
rect 9436 49478 9438 49530
rect 9276 49476 9300 49478
rect 9356 49476 9380 49478
rect 9436 49476 9460 49478
rect 9220 49456 9516 49476
rect 9220 48444 9516 48464
rect 9276 48442 9300 48444
rect 9356 48442 9380 48444
rect 9436 48442 9460 48444
rect 9298 48390 9300 48442
rect 9362 48390 9374 48442
rect 9436 48390 9438 48442
rect 9276 48388 9300 48390
rect 9356 48388 9380 48390
rect 9436 48388 9460 48390
rect 9220 48368 9516 48388
rect 9220 47356 9516 47376
rect 9276 47354 9300 47356
rect 9356 47354 9380 47356
rect 9436 47354 9460 47356
rect 9298 47302 9300 47354
rect 9362 47302 9374 47354
rect 9436 47302 9438 47354
rect 9276 47300 9300 47302
rect 9356 47300 9380 47302
rect 9436 47300 9460 47302
rect 9220 47280 9516 47300
rect 9220 46268 9516 46288
rect 9276 46266 9300 46268
rect 9356 46266 9380 46268
rect 9436 46266 9460 46268
rect 9298 46214 9300 46266
rect 9362 46214 9374 46266
rect 9436 46214 9438 46266
rect 9276 46212 9300 46214
rect 9356 46212 9380 46214
rect 9436 46212 9460 46214
rect 9220 46192 9516 46212
rect 9220 45180 9516 45200
rect 9276 45178 9300 45180
rect 9356 45178 9380 45180
rect 9436 45178 9460 45180
rect 9298 45126 9300 45178
rect 9362 45126 9374 45178
rect 9436 45126 9438 45178
rect 9276 45124 9300 45126
rect 9356 45124 9380 45126
rect 9436 45124 9460 45126
rect 9220 45104 9516 45124
rect 9220 44092 9516 44112
rect 9276 44090 9300 44092
rect 9356 44090 9380 44092
rect 9436 44090 9460 44092
rect 9298 44038 9300 44090
rect 9362 44038 9374 44090
rect 9436 44038 9438 44090
rect 9276 44036 9300 44038
rect 9356 44036 9380 44038
rect 9436 44036 9460 44038
rect 9220 44016 9516 44036
rect 9220 43004 9516 43024
rect 9276 43002 9300 43004
rect 9356 43002 9380 43004
rect 9436 43002 9460 43004
rect 9298 42950 9300 43002
rect 9362 42950 9374 43002
rect 9436 42950 9438 43002
rect 9276 42948 9300 42950
rect 9356 42948 9380 42950
rect 9436 42948 9460 42950
rect 9220 42928 9516 42948
rect 9220 41916 9516 41936
rect 9276 41914 9300 41916
rect 9356 41914 9380 41916
rect 9436 41914 9460 41916
rect 9298 41862 9300 41914
rect 9362 41862 9374 41914
rect 9436 41862 9438 41914
rect 9276 41860 9300 41862
rect 9356 41860 9380 41862
rect 9436 41860 9460 41862
rect 9220 41840 9516 41860
rect 9220 40828 9516 40848
rect 9276 40826 9300 40828
rect 9356 40826 9380 40828
rect 9436 40826 9460 40828
rect 9298 40774 9300 40826
rect 9362 40774 9374 40826
rect 9436 40774 9438 40826
rect 9276 40772 9300 40774
rect 9356 40772 9380 40774
rect 9436 40772 9460 40774
rect 9220 40752 9516 40772
rect 9220 39740 9516 39760
rect 9276 39738 9300 39740
rect 9356 39738 9380 39740
rect 9436 39738 9460 39740
rect 9298 39686 9300 39738
rect 9362 39686 9374 39738
rect 9436 39686 9438 39738
rect 9276 39684 9300 39686
rect 9356 39684 9380 39686
rect 9436 39684 9460 39686
rect 9220 39664 9516 39684
rect 9772 39432 9824 39438
rect 9772 39374 9824 39380
rect 9220 38652 9516 38672
rect 9276 38650 9300 38652
rect 9356 38650 9380 38652
rect 9436 38650 9460 38652
rect 9298 38598 9300 38650
rect 9362 38598 9374 38650
rect 9436 38598 9438 38650
rect 9276 38596 9300 38598
rect 9356 38596 9380 38598
rect 9436 38596 9460 38598
rect 9220 38576 9516 38596
rect 9220 37564 9516 37584
rect 9276 37562 9300 37564
rect 9356 37562 9380 37564
rect 9436 37562 9460 37564
rect 9298 37510 9300 37562
rect 9362 37510 9374 37562
rect 9436 37510 9438 37562
rect 9276 37508 9300 37510
rect 9356 37508 9380 37510
rect 9436 37508 9460 37510
rect 9220 37488 9516 37508
rect 9220 36476 9516 36496
rect 9276 36474 9300 36476
rect 9356 36474 9380 36476
rect 9436 36474 9460 36476
rect 9298 36422 9300 36474
rect 9362 36422 9374 36474
rect 9436 36422 9438 36474
rect 9276 36420 9300 36422
rect 9356 36420 9380 36422
rect 9436 36420 9460 36422
rect 9220 36400 9516 36420
rect 9220 35388 9516 35408
rect 9276 35386 9300 35388
rect 9356 35386 9380 35388
rect 9436 35386 9460 35388
rect 9298 35334 9300 35386
rect 9362 35334 9374 35386
rect 9436 35334 9438 35386
rect 9276 35332 9300 35334
rect 9356 35332 9380 35334
rect 9436 35332 9460 35334
rect 9220 35312 9516 35332
rect 9036 35080 9088 35086
rect 9036 35022 9088 35028
rect 9048 34746 9076 35022
rect 9036 34740 9088 34746
rect 9036 34682 9088 34688
rect 9048 34610 9076 34682
rect 9036 34604 9088 34610
rect 9036 34546 9088 34552
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 9220 34300 9516 34320
rect 9276 34298 9300 34300
rect 9356 34298 9380 34300
rect 9436 34298 9460 34300
rect 9298 34246 9300 34298
rect 9362 34246 9374 34298
rect 9436 34246 9438 34298
rect 9276 34244 9300 34246
rect 9356 34244 9380 34246
rect 9436 34244 9460 34246
rect 9220 34224 9516 34244
rect 9220 33212 9516 33232
rect 9276 33210 9300 33212
rect 9356 33210 9380 33212
rect 9436 33210 9460 33212
rect 9298 33158 9300 33210
rect 9362 33158 9374 33210
rect 9436 33158 9438 33210
rect 9276 33156 9300 33158
rect 9356 33156 9380 33158
rect 9436 33156 9460 33158
rect 9220 33136 9516 33156
rect 9220 32124 9516 32144
rect 9276 32122 9300 32124
rect 9356 32122 9380 32124
rect 9436 32122 9460 32124
rect 9298 32070 9300 32122
rect 9362 32070 9374 32122
rect 9436 32070 9438 32122
rect 9276 32068 9300 32070
rect 9356 32068 9380 32070
rect 9436 32068 9460 32070
rect 9220 32048 9516 32068
rect 9220 31036 9516 31056
rect 9276 31034 9300 31036
rect 9356 31034 9380 31036
rect 9436 31034 9460 31036
rect 9298 30982 9300 31034
rect 9362 30982 9374 31034
rect 9436 30982 9438 31034
rect 9276 30980 9300 30982
rect 9356 30980 9380 30982
rect 9436 30980 9460 30982
rect 9220 30960 9516 30980
rect 9220 29948 9516 29968
rect 9276 29946 9300 29948
rect 9356 29946 9380 29948
rect 9436 29946 9460 29948
rect 9298 29894 9300 29946
rect 9362 29894 9374 29946
rect 9436 29894 9438 29946
rect 9276 29892 9300 29894
rect 9356 29892 9380 29894
rect 9436 29892 9460 29894
rect 9220 29872 9516 29892
rect 9220 28860 9516 28880
rect 9276 28858 9300 28860
rect 9356 28858 9380 28860
rect 9436 28858 9460 28860
rect 9298 28806 9300 28858
rect 9362 28806 9374 28858
rect 9436 28806 9438 28858
rect 9276 28804 9300 28806
rect 9356 28804 9380 28806
rect 9436 28804 9460 28806
rect 9220 28784 9516 28804
rect 9220 27772 9516 27792
rect 9276 27770 9300 27772
rect 9356 27770 9380 27772
rect 9436 27770 9460 27772
rect 9298 27718 9300 27770
rect 9362 27718 9374 27770
rect 9436 27718 9438 27770
rect 9276 27716 9300 27718
rect 9356 27716 9380 27718
rect 9436 27716 9460 27718
rect 9220 27696 9516 27716
rect 9220 26684 9516 26704
rect 9276 26682 9300 26684
rect 9356 26682 9380 26684
rect 9436 26682 9460 26684
rect 9298 26630 9300 26682
rect 9362 26630 9374 26682
rect 9436 26630 9438 26682
rect 9276 26628 9300 26630
rect 9356 26628 9380 26630
rect 9436 26628 9460 26630
rect 9220 26608 9516 26628
rect 9600 26246 9628 34478
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 9220 25596 9516 25616
rect 9276 25594 9300 25596
rect 9356 25594 9380 25596
rect 9436 25594 9460 25596
rect 9298 25542 9300 25594
rect 9362 25542 9374 25594
rect 9436 25542 9438 25594
rect 9276 25540 9300 25542
rect 9356 25540 9380 25542
rect 9436 25540 9460 25542
rect 9220 25520 9516 25540
rect 9220 24508 9516 24528
rect 9276 24506 9300 24508
rect 9356 24506 9380 24508
rect 9436 24506 9460 24508
rect 9298 24454 9300 24506
rect 9362 24454 9374 24506
rect 9436 24454 9438 24506
rect 9276 24452 9300 24454
rect 9356 24452 9380 24454
rect 9436 24452 9460 24454
rect 9220 24432 9516 24452
rect 9220 23420 9516 23440
rect 9276 23418 9300 23420
rect 9356 23418 9380 23420
rect 9436 23418 9460 23420
rect 9298 23366 9300 23418
rect 9362 23366 9374 23418
rect 9436 23366 9438 23418
rect 9276 23364 9300 23366
rect 9356 23364 9380 23366
rect 9436 23364 9460 23366
rect 9220 23344 9516 23364
rect 9220 23248 9272 23254
rect 9220 23190 9272 23196
rect 9232 22710 9260 23190
rect 9220 22704 9272 22710
rect 9220 22646 9272 22652
rect 9220 22332 9516 22352
rect 9276 22330 9300 22332
rect 9356 22330 9380 22332
rect 9436 22330 9460 22332
rect 9298 22278 9300 22330
rect 9362 22278 9374 22330
rect 9436 22278 9438 22330
rect 9276 22276 9300 22278
rect 9356 22276 9380 22278
rect 9436 22276 9460 22278
rect 9220 22256 9516 22276
rect 9220 21244 9516 21264
rect 9276 21242 9300 21244
rect 9356 21242 9380 21244
rect 9436 21242 9460 21244
rect 9298 21190 9300 21242
rect 9362 21190 9374 21242
rect 9436 21190 9438 21242
rect 9276 21188 9300 21190
rect 9356 21188 9380 21190
rect 9436 21188 9460 21190
rect 9220 21168 9516 21188
rect 9220 20156 9516 20176
rect 9276 20154 9300 20156
rect 9356 20154 9380 20156
rect 9436 20154 9460 20156
rect 9298 20102 9300 20154
rect 9362 20102 9374 20154
rect 9436 20102 9438 20154
rect 9276 20100 9300 20102
rect 9356 20100 9380 20102
rect 9436 20100 9460 20102
rect 9220 20080 9516 20100
rect 9220 19068 9516 19088
rect 9276 19066 9300 19068
rect 9356 19066 9380 19068
rect 9436 19066 9460 19068
rect 9298 19014 9300 19066
rect 9362 19014 9374 19066
rect 9436 19014 9438 19066
rect 9276 19012 9300 19014
rect 9356 19012 9380 19014
rect 9436 19012 9460 19014
rect 9220 18992 9516 19012
rect 9220 17980 9516 18000
rect 9276 17978 9300 17980
rect 9356 17978 9380 17980
rect 9436 17978 9460 17980
rect 9298 17926 9300 17978
rect 9362 17926 9374 17978
rect 9436 17926 9438 17978
rect 9276 17924 9300 17926
rect 9356 17924 9380 17926
rect 9436 17924 9460 17926
rect 9220 17904 9516 17924
rect 9220 16892 9516 16912
rect 9276 16890 9300 16892
rect 9356 16890 9380 16892
rect 9436 16890 9460 16892
rect 9298 16838 9300 16890
rect 9362 16838 9374 16890
rect 9436 16838 9438 16890
rect 9276 16836 9300 16838
rect 9356 16836 9380 16838
rect 9436 16836 9460 16838
rect 9220 16816 9516 16836
rect 9220 15804 9516 15824
rect 9276 15802 9300 15804
rect 9356 15802 9380 15804
rect 9436 15802 9460 15804
rect 9298 15750 9300 15802
rect 9362 15750 9374 15802
rect 9436 15750 9438 15802
rect 9276 15748 9300 15750
rect 9356 15748 9380 15750
rect 9436 15748 9460 15750
rect 9220 15728 9516 15748
rect 9784 15162 9812 39374
rect 10152 34066 10180 66642
rect 11072 66502 11100 67050
rect 11704 67040 11756 67046
rect 11704 66982 11756 66988
rect 11060 66496 11112 66502
rect 11060 66438 11112 66444
rect 11072 66298 11100 66438
rect 11060 66292 11112 66298
rect 11060 66234 11112 66240
rect 11716 57526 11744 66982
rect 13544 66836 13596 66842
rect 13544 66778 13596 66784
rect 12900 63776 12952 63782
rect 12900 63718 12952 63724
rect 12912 63578 12940 63718
rect 12900 63572 12952 63578
rect 12900 63514 12952 63520
rect 12716 63436 12768 63442
rect 12716 63378 12768 63384
rect 12728 63238 12756 63378
rect 13176 63368 13228 63374
rect 13176 63310 13228 63316
rect 13188 63238 13216 63310
rect 12716 63232 12768 63238
rect 12716 63174 12768 63180
rect 13176 63232 13228 63238
rect 13176 63174 13228 63180
rect 12728 63034 12756 63174
rect 12716 63028 12768 63034
rect 12716 62970 12768 62976
rect 11704 57520 11756 57526
rect 11704 57462 11756 57468
rect 12624 56704 12676 56710
rect 12624 56646 12676 56652
rect 11060 55616 11112 55622
rect 11060 55558 11112 55564
rect 11072 55418 11100 55558
rect 11060 55412 11112 55418
rect 11060 55354 11112 55360
rect 12164 53440 12216 53446
rect 12164 53382 12216 53388
rect 11244 52556 11296 52562
rect 11244 52498 11296 52504
rect 10692 44328 10744 44334
rect 10692 44270 10744 44276
rect 10324 35488 10376 35494
rect 10324 35430 10376 35436
rect 10140 34060 10192 34066
rect 10140 34002 10192 34008
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9220 14716 9516 14736
rect 9276 14714 9300 14716
rect 9356 14714 9380 14716
rect 9436 14714 9460 14716
rect 9298 14662 9300 14714
rect 9362 14662 9374 14714
rect 9436 14662 9438 14714
rect 9276 14660 9300 14662
rect 9356 14660 9380 14662
rect 9436 14660 9460 14662
rect 9220 14640 9516 14660
rect 9220 13628 9516 13648
rect 9276 13626 9300 13628
rect 9356 13626 9380 13628
rect 9436 13626 9460 13628
rect 9298 13574 9300 13626
rect 9362 13574 9374 13626
rect 9436 13574 9438 13626
rect 9276 13572 9300 13574
rect 9356 13572 9380 13574
rect 9436 13572 9460 13574
rect 9220 13552 9516 13572
rect 9220 12540 9516 12560
rect 9276 12538 9300 12540
rect 9356 12538 9380 12540
rect 9436 12538 9460 12540
rect 9298 12486 9300 12538
rect 9362 12486 9374 12538
rect 9436 12486 9438 12538
rect 9276 12484 9300 12486
rect 9356 12484 9380 12486
rect 9436 12484 9460 12486
rect 9220 12464 9516 12484
rect 9680 12436 9732 12442
rect 10244 12434 10272 17206
rect 10336 16574 10364 35430
rect 10336 16546 10548 16574
rect 10520 12714 10548 16546
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 9680 12378 9732 12384
rect 10152 12406 10272 12434
rect 9220 11452 9516 11472
rect 9276 11450 9300 11452
rect 9356 11450 9380 11452
rect 9436 11450 9460 11452
rect 9298 11398 9300 11450
rect 9362 11398 9374 11450
rect 9436 11398 9438 11450
rect 9276 11396 9300 11398
rect 9356 11396 9380 11398
rect 9436 11396 9460 11398
rect 9220 11376 9516 11396
rect 9692 11257 9720 12378
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9678 11248 9734 11257
rect 9678 11183 9680 11192
rect 9732 11183 9734 11192
rect 9680 11154 9732 11160
rect 9968 10713 9996 11562
rect 10152 11558 10180 12406
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9954 10704 10010 10713
rect 9954 10639 10010 10648
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8496 800 8524 2858
rect 8588 2582 8616 9862
rect 8680 2990 8708 10406
rect 9220 10364 9516 10384
rect 9276 10362 9300 10364
rect 9356 10362 9380 10364
rect 9436 10362 9460 10364
rect 9298 10310 9300 10362
rect 9362 10310 9374 10362
rect 9436 10310 9438 10362
rect 9276 10308 9300 10310
rect 9356 10308 9380 10310
rect 9436 10308 9460 10310
rect 9220 10288 9516 10308
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 8772 9178 8800 9318
rect 9220 9276 9516 9296
rect 9276 9274 9300 9276
rect 9356 9274 9380 9276
rect 9436 9274 9460 9276
rect 9298 9222 9300 9274
rect 9362 9222 9374 9274
rect 9436 9222 9438 9274
rect 9276 9220 9300 9222
rect 9356 9220 9380 9222
rect 9436 9220 9460 9222
rect 9220 9200 9516 9220
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 4690 8800 8230
rect 8864 5166 8892 8774
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8772 2774 8800 4082
rect 8864 3398 8892 5102
rect 8956 4078 8984 7686
rect 9048 5302 9076 8298
rect 9220 8188 9516 8208
rect 9276 8186 9300 8188
rect 9356 8186 9380 8188
rect 9436 8186 9460 8188
rect 9298 8134 9300 8186
rect 9362 8134 9374 8186
rect 9436 8134 9438 8186
rect 9276 8132 9300 8134
rect 9356 8132 9380 8134
rect 9436 8132 9460 8134
rect 9220 8112 9516 8132
rect 9220 7100 9516 7120
rect 9276 7098 9300 7100
rect 9356 7098 9380 7100
rect 9436 7098 9460 7100
rect 9298 7046 9300 7098
rect 9362 7046 9374 7098
rect 9436 7046 9438 7098
rect 9276 7044 9300 7046
rect 9356 7044 9380 7046
rect 9436 7044 9460 7046
rect 9220 7024 9516 7044
rect 9600 6254 9628 9318
rect 9692 8634 9720 9454
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8942 3904 8998 3913
rect 8942 3839 8998 3848
rect 8956 3466 8984 3839
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8680 2746 8800 2774
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8680 1442 8708 2746
rect 8864 1562 8892 2926
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 8852 1556 8904 1562
rect 8852 1498 8904 1504
rect 8588 1414 8708 1442
rect 8760 1420 8812 1426
rect 8588 800 8616 1414
rect 8760 1362 8812 1368
rect 8772 800 8800 1362
rect 8956 800 8984 2858
rect 9048 800 9076 5238
rect 9140 1442 9168 6190
rect 9220 6012 9516 6032
rect 9276 6010 9300 6012
rect 9356 6010 9380 6012
rect 9436 6010 9460 6012
rect 9298 5958 9300 6010
rect 9362 5958 9374 6010
rect 9436 5958 9438 6010
rect 9276 5956 9300 5958
rect 9356 5956 9380 5958
rect 9436 5956 9460 5958
rect 9220 5936 9516 5956
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5302 9444 5510
rect 9404 5296 9456 5302
rect 9692 5250 9720 7686
rect 9784 6254 9812 9862
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9404 5238 9456 5244
rect 9600 5222 9720 5250
rect 9220 4924 9516 4944
rect 9276 4922 9300 4924
rect 9356 4922 9380 4924
rect 9436 4922 9460 4924
rect 9298 4870 9300 4922
rect 9362 4870 9374 4922
rect 9436 4870 9438 4922
rect 9276 4868 9300 4870
rect 9356 4868 9380 4870
rect 9436 4868 9460 4870
rect 9220 4848 9516 4868
rect 9600 4690 9628 5222
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9232 4049 9260 4626
rect 9600 4298 9628 4626
rect 9508 4270 9628 4298
rect 9508 4146 9536 4270
rect 9496 4140 9548 4146
rect 9692 4128 9720 5102
rect 9496 4082 9548 4088
rect 9600 4100 9720 4128
rect 9218 4040 9274 4049
rect 9218 3975 9274 3984
rect 9220 3836 9516 3856
rect 9276 3834 9300 3836
rect 9356 3834 9380 3836
rect 9436 3834 9460 3836
rect 9298 3782 9300 3834
rect 9362 3782 9374 3834
rect 9436 3782 9438 3834
rect 9276 3780 9300 3782
rect 9356 3780 9380 3782
rect 9436 3780 9460 3782
rect 9220 3760 9516 3780
rect 9220 2748 9516 2768
rect 9276 2746 9300 2748
rect 9356 2746 9380 2748
rect 9436 2746 9460 2748
rect 9298 2694 9300 2746
rect 9362 2694 9374 2746
rect 9436 2694 9438 2746
rect 9276 2692 9300 2694
rect 9356 2692 9380 2694
rect 9436 2692 9460 2694
rect 9220 2672 9516 2692
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9140 1414 9260 1442
rect 9232 800 9260 1414
rect 9324 800 9352 1498
rect 9600 1442 9628 4100
rect 9784 3924 9812 6190
rect 9876 5166 9904 8298
rect 9968 5794 9996 10639
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 5914 10088 8774
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9968 5766 10088 5794
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9508 1414 9628 1442
rect 9692 3896 9812 3924
rect 9508 800 9536 1414
rect 9692 1306 9720 3896
rect 9770 3768 9826 3777
rect 9770 3703 9826 3712
rect 9784 2922 9812 3703
rect 9876 3505 9904 4966
rect 9862 3496 9918 3505
rect 9862 3431 9918 3440
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9770 2816 9826 2825
rect 9770 2751 9826 2760
rect 9784 2582 9812 2751
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9876 1578 9904 3334
rect 9600 1278 9720 1306
rect 9784 1550 9904 1578
rect 9600 800 9628 1278
rect 9784 800 9812 1550
rect 9968 1442 9996 5578
rect 10060 3641 10088 5766
rect 10046 3632 10102 3641
rect 10152 3602 10180 11494
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 6866 10272 9862
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10046 3567 10102 3576
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10244 3482 10272 6802
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 9876 1414 9996 1442
rect 10060 3454 10272 3482
rect 9876 800 9904 1414
rect 10060 800 10088 3454
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10152 800 10180 2994
rect 10244 2514 10272 3334
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10336 800 10364 5714
rect 10428 800 10456 7278
rect 10520 3738 10548 12650
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10506 3632 10562 3641
rect 10506 3567 10562 3576
rect 10520 3074 10548 3567
rect 10612 3398 10640 11018
rect 10704 10538 10732 44270
rect 10876 30660 10928 30666
rect 10876 30602 10928 30608
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 5778 10732 8774
rect 10796 8634 10824 15506
rect 10888 11082 10916 30602
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11072 26246 11100 27066
rect 11060 26240 11112 26246
rect 11060 26182 11112 26188
rect 11072 22438 11100 26182
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10796 4826 10824 8298
rect 10888 7342 10916 9862
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10796 4690 10824 4762
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10888 4078 10916 6054
rect 10980 5030 11008 11086
rect 11164 10470 11192 17546
rect 11256 15706 11284 52498
rect 11796 49836 11848 49842
rect 11796 49778 11848 49784
rect 11704 44396 11756 44402
rect 11704 44338 11756 44344
rect 11612 34944 11664 34950
rect 11612 34886 11664 34892
rect 11624 34610 11652 34886
rect 11612 34604 11664 34610
rect 11612 34546 11664 34552
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11716 12434 11744 44338
rect 11808 22098 11836 49778
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11900 15366 11928 22374
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11624 12406 11744 12434
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 6254 11100 8774
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10704 3194 10732 4014
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10520 3046 10732 3074
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10520 1426 10548 2926
rect 10508 1420 10560 1426
rect 10508 1362 10560 1368
rect 10612 800 10640 2926
rect 10704 2582 10732 3046
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10796 800 10824 3946
rect 10980 3584 11008 4150
rect 11072 4010 11100 6190
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11058 3904 11114 3913
rect 11058 3839 11114 3848
rect 11072 3670 11100 3839
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11164 3602 11192 10406
rect 11256 7954 11284 10406
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 10888 3556 11008 3584
rect 11152 3596 11204 3602
rect 10888 2922 10916 3556
rect 11152 3538 11204 3544
rect 11256 3482 11284 7890
rect 11348 7342 11376 10474
rect 11440 7449 11468 12038
rect 11624 10062 11652 12406
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11612 10056 11664 10062
rect 11610 10024 11612 10033
rect 11664 10024 11666 10033
rect 11610 9959 11666 9968
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11426 7440 11482 7449
rect 11426 7375 11482 7384
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 10980 3454 11284 3482
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10980 2774 11008 3454
rect 11060 3392 11112 3398
rect 11112 3352 11192 3380
rect 11060 3334 11112 3340
rect 10888 2746 11008 2774
rect 10888 800 10916 2746
rect 11060 1148 11112 1154
rect 11060 1090 11112 1096
rect 11072 800 11100 1090
rect 11164 800 11192 3352
rect 11348 800 11376 7278
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11440 4690 11468 7210
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11440 4282 11468 4626
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11440 3618 11468 4082
rect 11532 4078 11560 7686
rect 11624 6866 11652 9862
rect 11716 7954 11744 11018
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11532 3777 11560 4014
rect 11518 3768 11574 3777
rect 11518 3703 11574 3712
rect 11440 3590 11560 3618
rect 11532 3126 11560 3590
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11428 1216 11480 1222
rect 11428 1158 11480 1164
rect 11440 800 11468 1158
rect 11624 800 11652 6802
rect 11716 800 11744 7890
rect 11808 2922 11836 12038
rect 11992 11558 12020 21422
rect 12084 14482 12112 30126
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12176 12646 12204 53382
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12360 23730 12388 24006
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 13530 12296 15302
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 4690 11928 7142
rect 11992 6798 12020 9454
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11992 4570 12020 6734
rect 12084 5778 12112 9318
rect 12176 7002 12204 12582
rect 12268 10674 12296 13466
rect 12636 12374 12664 56646
rect 13084 55616 13136 55622
rect 13084 55558 13136 55564
rect 12992 45416 13044 45422
rect 12992 45358 13044 45364
rect 13004 45082 13032 45358
rect 12992 45076 13044 45082
rect 12992 45018 13044 45024
rect 12992 43240 13044 43246
rect 12992 43182 13044 43188
rect 12808 42560 12860 42566
rect 12808 42502 12860 42508
rect 12820 42362 12848 42502
rect 12808 42356 12860 42362
rect 12808 42298 12860 42304
rect 12808 37936 12860 37942
rect 12808 37878 12860 37884
rect 12820 16574 12848 37878
rect 13004 35018 13032 43182
rect 12992 35012 13044 35018
rect 12992 34954 13044 34960
rect 13004 30394 13032 34954
rect 12992 30388 13044 30394
rect 12992 30330 13044 30336
rect 12728 16546 12848 16574
rect 12728 12646 12756 16546
rect 13096 14074 13124 55558
rect 13188 25838 13216 63174
rect 13452 58880 13504 58886
rect 13452 58822 13504 58828
rect 13360 43104 13412 43110
rect 13360 43046 13412 43052
rect 13372 42906 13400 43046
rect 13360 42900 13412 42906
rect 13360 42842 13412 42848
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 13188 25498 13216 25774
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13188 22710 13216 23258
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13372 12646 13400 13330
rect 12716 12640 12768 12646
rect 13360 12640 13412 12646
rect 12716 12582 12768 12588
rect 13358 12608 13360 12617
rect 13412 12608 13414 12617
rect 12728 12434 12756 12582
rect 13358 12543 13414 12552
rect 13464 12434 13492 58822
rect 13556 28218 13584 66778
rect 14220 66396 14516 66416
rect 14276 66394 14300 66396
rect 14356 66394 14380 66396
rect 14436 66394 14460 66396
rect 14298 66342 14300 66394
rect 14362 66342 14374 66394
rect 14436 66342 14438 66394
rect 14276 66340 14300 66342
rect 14356 66340 14380 66342
rect 14436 66340 14460 66342
rect 14220 66320 14516 66340
rect 14556 66088 14608 66094
rect 14556 66030 14608 66036
rect 14220 65308 14516 65328
rect 14276 65306 14300 65308
rect 14356 65306 14380 65308
rect 14436 65306 14460 65308
rect 14298 65254 14300 65306
rect 14362 65254 14374 65306
rect 14436 65254 14438 65306
rect 14276 65252 14300 65254
rect 14356 65252 14380 65254
rect 14436 65252 14460 65254
rect 14220 65232 14516 65252
rect 14220 64220 14516 64240
rect 14276 64218 14300 64220
rect 14356 64218 14380 64220
rect 14436 64218 14460 64220
rect 14298 64166 14300 64218
rect 14362 64166 14374 64218
rect 14436 64166 14438 64218
rect 14276 64164 14300 64166
rect 14356 64164 14380 64166
rect 14436 64164 14460 64166
rect 14220 64144 14516 64164
rect 14004 63912 14056 63918
rect 14004 63854 14056 63860
rect 13636 45008 13688 45014
rect 13636 44950 13688 44956
rect 13544 28212 13596 28218
rect 13544 28154 13596 28160
rect 13648 16574 13676 44950
rect 13820 41064 13872 41070
rect 13820 41006 13872 41012
rect 13556 16546 13676 16574
rect 13556 13190 13584 16546
rect 13544 13184 13596 13190
rect 13542 13152 13544 13161
rect 13596 13152 13598 13161
rect 13542 13087 13598 13096
rect 12728 12406 12848 12434
rect 12624 12368 12676 12374
rect 12544 12328 12624 12356
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 8537 12296 10610
rect 12254 8528 12310 8537
rect 12254 8463 12310 8472
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12162 6896 12218 6905
rect 12162 6831 12218 6840
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11900 4542 12020 4570
rect 11900 4146 11928 4542
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11900 800 11928 3946
rect 11992 800 12020 4082
rect 12084 3777 12112 5714
rect 12176 5370 12204 6831
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12176 4214 12204 5306
rect 12268 4690 12296 8230
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12254 4040 12310 4049
rect 12070 3768 12126 3777
rect 12070 3703 12126 3712
rect 12176 3074 12204 4014
rect 12254 3975 12256 3984
rect 12308 3975 12310 3984
rect 12256 3946 12308 3952
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12084 3046 12204 3074
rect 12084 2836 12112 3046
rect 12084 2808 12204 2836
rect 12176 800 12204 2808
rect 12268 1222 12296 3470
rect 12360 2582 12388 11494
rect 12544 10130 12572 12328
rect 12624 12310 12676 12316
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 6866 12480 9862
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12452 4146 12480 6802
rect 12544 6798 12572 9930
rect 12636 7954 12664 11494
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12438 3768 12494 3777
rect 12438 3703 12494 3712
rect 12452 3398 12480 3703
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12452 2394 12480 3334
rect 12360 2366 12480 2394
rect 12360 1834 12388 2366
rect 12348 1828 12400 1834
rect 12348 1770 12400 1776
rect 12348 1692 12400 1698
rect 12348 1634 12400 1640
rect 12256 1216 12308 1222
rect 12256 1158 12308 1164
rect 12360 800 12388 1634
rect 12544 1442 12572 6734
rect 12452 1414 12572 1442
rect 12452 800 12480 1414
rect 12636 800 12664 7890
rect 12728 7886 12756 11018
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12728 4146 12756 7822
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12728 800 12756 3946
rect 12820 2990 12848 12406
rect 13372 12406 13492 12434
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 7342 12940 10406
rect 13004 8430 13032 11494
rect 13372 11286 13400 12406
rect 13832 12238 13860 41006
rect 14016 26858 14044 63854
rect 14220 63132 14516 63152
rect 14276 63130 14300 63132
rect 14356 63130 14380 63132
rect 14436 63130 14460 63132
rect 14298 63078 14300 63130
rect 14362 63078 14374 63130
rect 14436 63078 14438 63130
rect 14276 63076 14300 63078
rect 14356 63076 14380 63078
rect 14436 63076 14460 63078
rect 14220 63056 14516 63076
rect 14220 62044 14516 62064
rect 14276 62042 14300 62044
rect 14356 62042 14380 62044
rect 14436 62042 14460 62044
rect 14298 61990 14300 62042
rect 14362 61990 14374 62042
rect 14436 61990 14438 62042
rect 14276 61988 14300 61990
rect 14356 61988 14380 61990
rect 14436 61988 14460 61990
rect 14220 61968 14516 61988
rect 14220 60956 14516 60976
rect 14276 60954 14300 60956
rect 14356 60954 14380 60956
rect 14436 60954 14460 60956
rect 14298 60902 14300 60954
rect 14362 60902 14374 60954
rect 14436 60902 14438 60954
rect 14276 60900 14300 60902
rect 14356 60900 14380 60902
rect 14436 60900 14460 60902
rect 14220 60880 14516 60900
rect 14220 59868 14516 59888
rect 14276 59866 14300 59868
rect 14356 59866 14380 59868
rect 14436 59866 14460 59868
rect 14298 59814 14300 59866
rect 14362 59814 14374 59866
rect 14436 59814 14438 59866
rect 14276 59812 14300 59814
rect 14356 59812 14380 59814
rect 14436 59812 14460 59814
rect 14220 59792 14516 59812
rect 14220 58780 14516 58800
rect 14276 58778 14300 58780
rect 14356 58778 14380 58780
rect 14436 58778 14460 58780
rect 14298 58726 14300 58778
rect 14362 58726 14374 58778
rect 14436 58726 14438 58778
rect 14276 58724 14300 58726
rect 14356 58724 14380 58726
rect 14436 58724 14460 58726
rect 14220 58704 14516 58724
rect 14220 57692 14516 57712
rect 14276 57690 14300 57692
rect 14356 57690 14380 57692
rect 14436 57690 14460 57692
rect 14298 57638 14300 57690
rect 14362 57638 14374 57690
rect 14436 57638 14438 57690
rect 14276 57636 14300 57638
rect 14356 57636 14380 57638
rect 14436 57636 14460 57638
rect 14220 57616 14516 57636
rect 14220 56604 14516 56624
rect 14276 56602 14300 56604
rect 14356 56602 14380 56604
rect 14436 56602 14460 56604
rect 14298 56550 14300 56602
rect 14362 56550 14374 56602
rect 14436 56550 14438 56602
rect 14276 56548 14300 56550
rect 14356 56548 14380 56550
rect 14436 56548 14460 56550
rect 14220 56528 14516 56548
rect 14220 55516 14516 55536
rect 14276 55514 14300 55516
rect 14356 55514 14380 55516
rect 14436 55514 14460 55516
rect 14298 55462 14300 55514
rect 14362 55462 14374 55514
rect 14436 55462 14438 55514
rect 14276 55460 14300 55462
rect 14356 55460 14380 55462
rect 14436 55460 14460 55462
rect 14220 55440 14516 55460
rect 14220 54428 14516 54448
rect 14276 54426 14300 54428
rect 14356 54426 14380 54428
rect 14436 54426 14460 54428
rect 14298 54374 14300 54426
rect 14362 54374 14374 54426
rect 14436 54374 14438 54426
rect 14276 54372 14300 54374
rect 14356 54372 14380 54374
rect 14436 54372 14460 54374
rect 14220 54352 14516 54372
rect 14220 53340 14516 53360
rect 14276 53338 14300 53340
rect 14356 53338 14380 53340
rect 14436 53338 14460 53340
rect 14298 53286 14300 53338
rect 14362 53286 14374 53338
rect 14436 53286 14438 53338
rect 14276 53284 14300 53286
rect 14356 53284 14380 53286
rect 14436 53284 14460 53286
rect 14220 53264 14516 53284
rect 14220 52252 14516 52272
rect 14276 52250 14300 52252
rect 14356 52250 14380 52252
rect 14436 52250 14460 52252
rect 14298 52198 14300 52250
rect 14362 52198 14374 52250
rect 14436 52198 14438 52250
rect 14276 52196 14300 52198
rect 14356 52196 14380 52198
rect 14436 52196 14460 52198
rect 14220 52176 14516 52196
rect 14220 51164 14516 51184
rect 14276 51162 14300 51164
rect 14356 51162 14380 51164
rect 14436 51162 14460 51164
rect 14298 51110 14300 51162
rect 14362 51110 14374 51162
rect 14436 51110 14438 51162
rect 14276 51108 14300 51110
rect 14356 51108 14380 51110
rect 14436 51108 14460 51110
rect 14220 51088 14516 51108
rect 14220 50076 14516 50096
rect 14276 50074 14300 50076
rect 14356 50074 14380 50076
rect 14436 50074 14460 50076
rect 14298 50022 14300 50074
rect 14362 50022 14374 50074
rect 14436 50022 14438 50074
rect 14276 50020 14300 50022
rect 14356 50020 14380 50022
rect 14436 50020 14460 50022
rect 14220 50000 14516 50020
rect 14220 48988 14516 49008
rect 14276 48986 14300 48988
rect 14356 48986 14380 48988
rect 14436 48986 14460 48988
rect 14298 48934 14300 48986
rect 14362 48934 14374 48986
rect 14436 48934 14438 48986
rect 14276 48932 14300 48934
rect 14356 48932 14380 48934
rect 14436 48932 14460 48934
rect 14220 48912 14516 48932
rect 14220 47900 14516 47920
rect 14276 47898 14300 47900
rect 14356 47898 14380 47900
rect 14436 47898 14460 47900
rect 14298 47846 14300 47898
rect 14362 47846 14374 47898
rect 14436 47846 14438 47898
rect 14276 47844 14300 47846
rect 14356 47844 14380 47846
rect 14436 47844 14460 47846
rect 14220 47824 14516 47844
rect 14220 46812 14516 46832
rect 14276 46810 14300 46812
rect 14356 46810 14380 46812
rect 14436 46810 14460 46812
rect 14298 46758 14300 46810
rect 14362 46758 14374 46810
rect 14436 46758 14438 46810
rect 14276 46756 14300 46758
rect 14356 46756 14380 46758
rect 14436 46756 14460 46758
rect 14220 46736 14516 46756
rect 14220 45724 14516 45744
rect 14276 45722 14300 45724
rect 14356 45722 14380 45724
rect 14436 45722 14460 45724
rect 14298 45670 14300 45722
rect 14362 45670 14374 45722
rect 14436 45670 14438 45722
rect 14276 45668 14300 45670
rect 14356 45668 14380 45670
rect 14436 45668 14460 45670
rect 14220 45648 14516 45668
rect 14220 44636 14516 44656
rect 14276 44634 14300 44636
rect 14356 44634 14380 44636
rect 14436 44634 14460 44636
rect 14298 44582 14300 44634
rect 14362 44582 14374 44634
rect 14436 44582 14438 44634
rect 14276 44580 14300 44582
rect 14356 44580 14380 44582
rect 14436 44580 14460 44582
rect 14220 44560 14516 44580
rect 14220 43548 14516 43568
rect 14276 43546 14300 43548
rect 14356 43546 14380 43548
rect 14436 43546 14460 43548
rect 14298 43494 14300 43546
rect 14362 43494 14374 43546
rect 14436 43494 14438 43546
rect 14276 43492 14300 43494
rect 14356 43492 14380 43494
rect 14436 43492 14460 43494
rect 14220 43472 14516 43492
rect 14220 42460 14516 42480
rect 14276 42458 14300 42460
rect 14356 42458 14380 42460
rect 14436 42458 14460 42460
rect 14298 42406 14300 42458
rect 14362 42406 14374 42458
rect 14436 42406 14438 42458
rect 14276 42404 14300 42406
rect 14356 42404 14380 42406
rect 14436 42404 14460 42406
rect 14220 42384 14516 42404
rect 14220 41372 14516 41392
rect 14276 41370 14300 41372
rect 14356 41370 14380 41372
rect 14436 41370 14460 41372
rect 14298 41318 14300 41370
rect 14362 41318 14374 41370
rect 14436 41318 14438 41370
rect 14276 41316 14300 41318
rect 14356 41316 14380 41318
rect 14436 41316 14460 41318
rect 14220 41296 14516 41316
rect 14220 40284 14516 40304
rect 14276 40282 14300 40284
rect 14356 40282 14380 40284
rect 14436 40282 14460 40284
rect 14298 40230 14300 40282
rect 14362 40230 14374 40282
rect 14436 40230 14438 40282
rect 14276 40228 14300 40230
rect 14356 40228 14380 40230
rect 14436 40228 14460 40230
rect 14220 40208 14516 40228
rect 14220 39196 14516 39216
rect 14276 39194 14300 39196
rect 14356 39194 14380 39196
rect 14436 39194 14460 39196
rect 14298 39142 14300 39194
rect 14362 39142 14374 39194
rect 14436 39142 14438 39194
rect 14276 39140 14300 39142
rect 14356 39140 14380 39142
rect 14436 39140 14460 39142
rect 14220 39120 14516 39140
rect 14220 38108 14516 38128
rect 14276 38106 14300 38108
rect 14356 38106 14380 38108
rect 14436 38106 14460 38108
rect 14298 38054 14300 38106
rect 14362 38054 14374 38106
rect 14436 38054 14438 38106
rect 14276 38052 14300 38054
rect 14356 38052 14380 38054
rect 14436 38052 14460 38054
rect 14220 38032 14516 38052
rect 14220 37020 14516 37040
rect 14276 37018 14300 37020
rect 14356 37018 14380 37020
rect 14436 37018 14460 37020
rect 14298 36966 14300 37018
rect 14362 36966 14374 37018
rect 14436 36966 14438 37018
rect 14276 36964 14300 36966
rect 14356 36964 14380 36966
rect 14436 36964 14460 36966
rect 14220 36944 14516 36964
rect 14220 35932 14516 35952
rect 14276 35930 14300 35932
rect 14356 35930 14380 35932
rect 14436 35930 14460 35932
rect 14298 35878 14300 35930
rect 14362 35878 14374 35930
rect 14436 35878 14438 35930
rect 14276 35876 14300 35878
rect 14356 35876 14380 35878
rect 14436 35876 14460 35878
rect 14220 35856 14516 35876
rect 14220 34844 14516 34864
rect 14276 34842 14300 34844
rect 14356 34842 14380 34844
rect 14436 34842 14460 34844
rect 14298 34790 14300 34842
rect 14362 34790 14374 34842
rect 14436 34790 14438 34842
rect 14276 34788 14300 34790
rect 14356 34788 14380 34790
rect 14436 34788 14460 34790
rect 14220 34768 14516 34788
rect 14220 33756 14516 33776
rect 14276 33754 14300 33756
rect 14356 33754 14380 33756
rect 14436 33754 14460 33756
rect 14298 33702 14300 33754
rect 14362 33702 14374 33754
rect 14436 33702 14438 33754
rect 14276 33700 14300 33702
rect 14356 33700 14380 33702
rect 14436 33700 14460 33702
rect 14220 33680 14516 33700
rect 14220 32668 14516 32688
rect 14276 32666 14300 32668
rect 14356 32666 14380 32668
rect 14436 32666 14460 32668
rect 14298 32614 14300 32666
rect 14362 32614 14374 32666
rect 14436 32614 14438 32666
rect 14276 32612 14300 32614
rect 14356 32612 14380 32614
rect 14436 32612 14460 32614
rect 14220 32592 14516 32612
rect 14220 31580 14516 31600
rect 14276 31578 14300 31580
rect 14356 31578 14380 31580
rect 14436 31578 14460 31580
rect 14298 31526 14300 31578
rect 14362 31526 14374 31578
rect 14436 31526 14438 31578
rect 14276 31524 14300 31526
rect 14356 31524 14380 31526
rect 14436 31524 14460 31526
rect 14220 31504 14516 31524
rect 14220 30492 14516 30512
rect 14276 30490 14300 30492
rect 14356 30490 14380 30492
rect 14436 30490 14460 30492
rect 14298 30438 14300 30490
rect 14362 30438 14374 30490
rect 14436 30438 14438 30490
rect 14276 30436 14300 30438
rect 14356 30436 14380 30438
rect 14436 30436 14460 30438
rect 14220 30416 14516 30436
rect 14220 29404 14516 29424
rect 14276 29402 14300 29404
rect 14356 29402 14380 29404
rect 14436 29402 14460 29404
rect 14298 29350 14300 29402
rect 14362 29350 14374 29402
rect 14436 29350 14438 29402
rect 14276 29348 14300 29350
rect 14356 29348 14380 29350
rect 14436 29348 14460 29350
rect 14220 29328 14516 29348
rect 14220 28316 14516 28336
rect 14276 28314 14300 28316
rect 14356 28314 14380 28316
rect 14436 28314 14460 28316
rect 14298 28262 14300 28314
rect 14362 28262 14374 28314
rect 14436 28262 14438 28314
rect 14276 28260 14300 28262
rect 14356 28260 14380 28262
rect 14436 28260 14460 28262
rect 14220 28240 14516 28260
rect 14220 27228 14516 27248
rect 14276 27226 14300 27228
rect 14356 27226 14380 27228
rect 14436 27226 14460 27228
rect 14298 27174 14300 27226
rect 14362 27174 14374 27226
rect 14436 27174 14438 27226
rect 14276 27172 14300 27174
rect 14356 27172 14380 27174
rect 14436 27172 14460 27174
rect 14220 27152 14516 27172
rect 14004 26852 14056 26858
rect 14004 26794 14056 26800
rect 14220 26140 14516 26160
rect 14276 26138 14300 26140
rect 14356 26138 14380 26140
rect 14436 26138 14460 26140
rect 14298 26086 14300 26138
rect 14362 26086 14374 26138
rect 14436 26086 14438 26138
rect 14276 26084 14300 26086
rect 14356 26084 14380 26086
rect 14436 26084 14460 26086
rect 14220 26064 14516 26084
rect 14220 25052 14516 25072
rect 14276 25050 14300 25052
rect 14356 25050 14380 25052
rect 14436 25050 14460 25052
rect 14298 24998 14300 25050
rect 14362 24998 14374 25050
rect 14436 24998 14438 25050
rect 14276 24996 14300 24998
rect 14356 24996 14380 24998
rect 14436 24996 14460 24998
rect 14220 24976 14516 24996
rect 14220 23964 14516 23984
rect 14276 23962 14300 23964
rect 14356 23962 14380 23964
rect 14436 23962 14460 23964
rect 14298 23910 14300 23962
rect 14362 23910 14374 23962
rect 14436 23910 14438 23962
rect 14276 23908 14300 23910
rect 14356 23908 14380 23910
rect 14436 23908 14460 23910
rect 14220 23888 14516 23908
rect 14220 22876 14516 22896
rect 14276 22874 14300 22876
rect 14356 22874 14380 22876
rect 14436 22874 14460 22876
rect 14298 22822 14300 22874
rect 14362 22822 14374 22874
rect 14436 22822 14438 22874
rect 14276 22820 14300 22822
rect 14356 22820 14380 22822
rect 14436 22820 14460 22822
rect 14220 22800 14516 22820
rect 14220 21788 14516 21808
rect 14276 21786 14300 21788
rect 14356 21786 14380 21788
rect 14436 21786 14460 21788
rect 14298 21734 14300 21786
rect 14362 21734 14374 21786
rect 14436 21734 14438 21786
rect 14276 21732 14300 21734
rect 14356 21732 14380 21734
rect 14436 21732 14460 21734
rect 14220 21712 14516 21732
rect 14220 20700 14516 20720
rect 14276 20698 14300 20700
rect 14356 20698 14380 20700
rect 14436 20698 14460 20700
rect 14298 20646 14300 20698
rect 14362 20646 14374 20698
rect 14436 20646 14438 20698
rect 14276 20644 14300 20646
rect 14356 20644 14380 20646
rect 14436 20644 14460 20646
rect 14220 20624 14516 20644
rect 14220 19612 14516 19632
rect 14276 19610 14300 19612
rect 14356 19610 14380 19612
rect 14436 19610 14460 19612
rect 14298 19558 14300 19610
rect 14362 19558 14374 19610
rect 14436 19558 14438 19610
rect 14276 19556 14300 19558
rect 14356 19556 14380 19558
rect 14436 19556 14460 19558
rect 14220 19536 14516 19556
rect 14568 19334 14596 66030
rect 14832 59628 14884 59634
rect 14832 59570 14884 59576
rect 14844 59430 14872 59570
rect 14832 59424 14884 59430
rect 14832 59366 14884 59372
rect 14844 19922 14872 59366
rect 15844 51944 15896 51950
rect 15844 51886 15896 51892
rect 15200 30388 15252 30394
rect 15200 30330 15252 30336
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14568 19306 14688 19334
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13924 16574 13952 18770
rect 14220 18524 14516 18544
rect 14276 18522 14300 18524
rect 14356 18522 14380 18524
rect 14436 18522 14460 18524
rect 14298 18470 14300 18522
rect 14362 18470 14374 18522
rect 14436 18470 14438 18522
rect 14276 18468 14300 18470
rect 14356 18468 14380 18470
rect 14436 18468 14460 18470
rect 14220 18448 14516 18468
rect 14220 17436 14516 17456
rect 14276 17434 14300 17436
rect 14356 17434 14380 17436
rect 14436 17434 14460 17436
rect 14298 17382 14300 17434
rect 14362 17382 14374 17434
rect 14436 17382 14438 17434
rect 14276 17380 14300 17382
rect 14356 17380 14380 17382
rect 14436 17380 14460 17382
rect 14220 17360 14516 17380
rect 13924 16546 14044 16574
rect 14016 13954 14044 16546
rect 14220 16348 14516 16368
rect 14276 16346 14300 16348
rect 14356 16346 14380 16348
rect 14436 16346 14460 16348
rect 14298 16294 14300 16346
rect 14362 16294 14374 16346
rect 14436 16294 14438 16346
rect 14276 16292 14300 16294
rect 14356 16292 14380 16294
rect 14436 16292 14460 16294
rect 14220 16272 14516 16292
rect 14220 15260 14516 15280
rect 14276 15258 14300 15260
rect 14356 15258 14380 15260
rect 14436 15258 14460 15260
rect 14298 15206 14300 15258
rect 14362 15206 14374 15258
rect 14436 15206 14438 15258
rect 14276 15204 14300 15206
rect 14356 15204 14380 15206
rect 14436 15204 14460 15206
rect 14220 15184 14516 15204
rect 14220 14172 14516 14192
rect 14276 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14298 14118 14300 14170
rect 14362 14118 14374 14170
rect 14436 14118 14438 14170
rect 14276 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14220 14096 14516 14116
rect 14660 14006 14688 19306
rect 15028 16574 15056 21558
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 14844 16546 15056 16574
rect 14648 14000 14700 14006
rect 14016 13926 14596 13954
rect 14648 13942 14700 13948
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14108 13734 14136 13806
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 12434 14136 13670
rect 14220 13084 14516 13104
rect 14276 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14298 13030 14300 13082
rect 14362 13030 14374 13082
rect 14436 13030 14438 13082
rect 14276 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14220 13008 14516 13028
rect 14016 12406 14136 12434
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13910 12200 13966 12209
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 9722 13124 10474
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12820 1154 12848 2790
rect 12808 1148 12860 1154
rect 12808 1090 12860 1096
rect 12912 800 12940 7278
rect 13004 800 13032 8366
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13096 3670 13124 6938
rect 13188 6254 13216 9318
rect 13280 7342 13308 11018
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13188 5953 13216 6190
rect 13174 5944 13230 5953
rect 13174 5879 13230 5888
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13082 2680 13138 2689
rect 13082 2615 13138 2624
rect 13096 2582 13124 2615
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 13188 800 13216 3946
rect 13280 800 13308 7278
rect 13372 5914 13400 9318
rect 13464 9042 13492 12038
rect 13832 11393 13860 12174
rect 13910 12135 13966 12144
rect 13818 11384 13874 11393
rect 13818 11319 13874 11328
rect 13924 11234 13952 12135
rect 13832 11206 13952 11234
rect 13832 10554 13860 11206
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13740 10526 13860 10554
rect 13740 9738 13768 10526
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13648 9710 13768 9738
rect 13648 9450 13676 9710
rect 13832 9602 13860 10406
rect 13740 9574 13860 9602
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13372 4622 13400 5102
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13358 3768 13414 3777
rect 13358 3703 13414 3712
rect 13372 3670 13400 3703
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 1698 13400 3334
rect 13360 1692 13412 1698
rect 13360 1634 13412 1640
rect 13464 800 13492 8978
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 5166 13584 8774
rect 13648 7721 13676 9386
rect 13634 7712 13690 7721
rect 13634 7647 13690 7656
rect 13740 6866 13768 9574
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 5817 13676 6122
rect 13634 5808 13690 5817
rect 13740 5778 13768 6598
rect 13634 5743 13690 5752
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13556 3913 13584 4626
rect 13648 4214 13676 4694
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13636 3936 13688 3942
rect 13542 3904 13598 3913
rect 13636 3878 13688 3884
rect 13542 3839 13598 3848
rect 13556 3670 13584 3839
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13556 1562 13584 3130
rect 13544 1556 13596 1562
rect 13544 1498 13596 1504
rect 13648 1442 13676 3878
rect 13740 2961 13768 5714
rect 13726 2952 13782 2961
rect 13726 2887 13782 2896
rect 13832 2774 13860 9454
rect 13924 7954 13952 11018
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13740 2746 13860 2774
rect 13924 2774 13952 7890
rect 14016 4010 14044 12406
rect 14568 12322 14596 13926
rect 14108 12294 14596 12322
rect 14108 10266 14136 12294
rect 14220 11996 14516 12016
rect 14276 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14298 11942 14300 11994
rect 14362 11942 14374 11994
rect 14436 11942 14438 11994
rect 14276 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14220 11920 14516 11940
rect 14220 10908 14516 10928
rect 14276 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14298 10854 14300 10906
rect 14362 10854 14374 10906
rect 14436 10854 14438 10906
rect 14276 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14220 10832 14516 10852
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14476 10577 14504 10678
rect 14462 10568 14518 10577
rect 14462 10503 14518 10512
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14108 9081 14136 10202
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14476 9908 14504 10066
rect 14568 10033 14596 10406
rect 14554 10024 14610 10033
rect 14554 9959 14610 9968
rect 14476 9880 14596 9908
rect 14220 9820 14516 9840
rect 14276 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14298 9766 14300 9818
rect 14362 9766 14374 9818
rect 14436 9766 14438 9818
rect 14276 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14220 9744 14516 9764
rect 14370 9688 14426 9697
rect 14370 9623 14426 9632
rect 14094 9072 14150 9081
rect 14094 9007 14150 9016
rect 14096 8968 14148 8974
rect 14384 8945 14412 9623
rect 14096 8910 14148 8916
rect 14370 8936 14426 8945
rect 14108 6186 14136 8910
rect 14370 8871 14426 8880
rect 14220 8732 14516 8752
rect 14276 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14298 8678 14300 8730
rect 14362 8678 14374 8730
rect 14436 8678 14438 8730
rect 14276 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14220 8656 14516 8676
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14476 7834 14504 8434
rect 14568 8090 14596 9880
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14476 7806 14596 7834
rect 14220 7644 14516 7664
rect 14276 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14298 7590 14300 7642
rect 14362 7590 14374 7642
rect 14436 7590 14438 7642
rect 14276 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14220 7568 14516 7588
rect 14220 6556 14516 6576
rect 14276 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14298 6502 14300 6554
rect 14362 6502 14374 6554
rect 14436 6502 14438 6554
rect 14276 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14220 6480 14516 6500
rect 14462 6352 14518 6361
rect 14462 6287 14518 6296
rect 14476 6254 14504 6287
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14476 5642 14504 6190
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14220 5468 14516 5488
rect 14276 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14298 5414 14300 5466
rect 14362 5414 14374 5466
rect 14436 5414 14438 5466
rect 14276 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14220 5392 14516 5412
rect 14568 5234 14596 7806
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14660 5098 14688 13942
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 10169 14780 12038
rect 14844 11665 14872 16546
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14830 11656 14886 11665
rect 14830 11591 14886 11600
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14844 10305 14872 11494
rect 14830 10296 14886 10305
rect 14830 10231 14886 10240
rect 14738 10160 14794 10169
rect 14738 10095 14794 10104
rect 14832 9716 14884 9722
rect 14738 9688 14794 9697
rect 14832 9658 14884 9664
rect 14738 9623 14794 9632
rect 14752 9042 14780 9623
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 14004 4004 14056 4010
rect 14004 3946 14056 3952
rect 14002 3904 14058 3913
rect 14002 3839 14058 3848
rect 14016 2990 14044 3839
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13924 2746 14044 2774
rect 13740 2394 13768 2746
rect 13818 2680 13874 2689
rect 13818 2615 13874 2624
rect 13832 2582 13860 2615
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 13740 2366 13860 2394
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13740 1970 13768 2246
rect 13728 1964 13780 1970
rect 13728 1906 13780 1912
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13556 1414 13676 1442
rect 13556 800 13584 1414
rect 13740 800 13768 1498
rect 13832 800 13860 2366
rect 13924 2106 13952 2450
rect 13912 2100 13964 2106
rect 13912 2042 13964 2048
rect 13912 1760 13964 1766
rect 13912 1702 13964 1708
rect 13924 1306 13952 1702
rect 14016 1442 14044 2746
rect 14108 2514 14136 4626
rect 14476 4570 14504 5034
rect 14476 4542 14596 4570
rect 14220 4380 14516 4400
rect 14276 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14298 4326 14300 4378
rect 14362 4326 14374 4378
rect 14436 4326 14438 4378
rect 14276 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14220 4304 14516 4324
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14462 4040 14518 4049
rect 14384 3913 14412 4014
rect 14462 3975 14464 3984
rect 14516 3975 14518 3984
rect 14464 3946 14516 3952
rect 14370 3904 14426 3913
rect 14370 3839 14426 3848
rect 14220 3292 14516 3312
rect 14276 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14298 3238 14300 3290
rect 14362 3238 14374 3290
rect 14436 3238 14438 3290
rect 14276 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14220 3216 14516 3236
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 2038 14136 2246
rect 14220 2204 14516 2224
rect 14276 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14298 2150 14300 2202
rect 14362 2150 14374 2202
rect 14436 2150 14438 2202
rect 14276 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14220 2128 14516 2148
rect 14096 2032 14148 2038
rect 14096 1974 14148 1980
rect 14280 1692 14332 1698
rect 14280 1634 14332 1640
rect 14016 1414 14228 1442
rect 13924 1278 14044 1306
rect 14016 800 14044 1278
rect 14200 800 14228 1414
rect 14292 800 14320 1634
rect 14568 1442 14596 4542
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14660 1766 14688 4490
rect 14648 1760 14700 1766
rect 14648 1702 14700 1708
rect 14752 1698 14780 8978
rect 14844 8362 14872 9658
rect 14936 9518 14964 11494
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14922 9344 14978 9353
rect 14922 9279 14978 9288
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14740 1692 14792 1698
rect 14740 1634 14792 1640
rect 14844 1578 14872 8298
rect 14936 8242 14964 9279
rect 15028 8430 15056 12038
rect 15120 11218 15148 18906
rect 15212 12102 15240 30330
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15304 25294 15332 25842
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15304 16574 15332 25230
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15304 16546 15516 16574
rect 15488 12986 15516 16546
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15672 13274 15700 13806
rect 15580 13258 15700 13274
rect 15568 13252 15700 13258
rect 15620 13246 15700 13252
rect 15568 13194 15620 13200
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15488 12646 15516 12922
rect 15672 12730 15700 13246
rect 15764 12918 15792 18566
rect 15856 17338 15884 51886
rect 16592 50930 16620 67050
rect 19064 67040 19116 67046
rect 19064 66982 19116 66988
rect 25596 67040 25648 67046
rect 25596 66982 25648 66988
rect 18052 66632 18104 66638
rect 18052 66574 18104 66580
rect 16672 65748 16724 65754
rect 16672 65690 16724 65696
rect 16684 64054 16712 65690
rect 17132 65000 17184 65006
rect 17132 64942 17184 64948
rect 16672 64048 16724 64054
rect 16672 63990 16724 63996
rect 16684 59566 16712 63990
rect 16672 59560 16724 59566
rect 16672 59502 16724 59508
rect 16580 50924 16632 50930
rect 16580 50866 16632 50872
rect 16948 41472 17000 41478
rect 16948 41414 17000 41420
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16684 27402 16712 29242
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16396 18896 16448 18902
rect 16396 18838 16448 18844
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15844 13864 15896 13870
rect 15842 13832 15844 13841
rect 15896 13832 15898 13841
rect 15842 13767 15898 13776
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15672 12702 15792 12730
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15120 8498 15148 11154
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15212 10130 15240 10474
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15198 10024 15254 10033
rect 15198 9959 15254 9968
rect 15212 9722 15240 9959
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15212 8294 15240 9454
rect 15304 8498 15332 10202
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15396 8378 15424 11018
rect 15488 9518 15516 11018
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15304 8350 15424 8378
rect 15200 8288 15252 8294
rect 14936 8214 15148 8242
rect 15200 8230 15252 8236
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14936 2825 14964 5170
rect 15028 2990 15056 8026
rect 15120 3602 15148 8214
rect 15304 7818 15332 8350
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15212 4690 15240 7754
rect 15304 7342 15332 7754
rect 15396 7342 15424 8230
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 6458 15424 6802
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15488 6089 15516 9318
rect 15580 6254 15608 9862
rect 15672 9042 15700 11494
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15290 6080 15346 6089
rect 15290 6015 15346 6024
rect 15474 6080 15530 6089
rect 15474 6015 15530 6024
rect 15304 5846 15332 6015
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 14922 2816 14978 2825
rect 15212 2774 15240 4490
rect 15396 3738 15424 5714
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15488 3777 15516 5646
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15474 3768 15530 3777
rect 15384 3732 15436 3738
rect 15580 3754 15608 5102
rect 15672 3890 15700 8978
rect 15764 4078 15792 12702
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 7041 15884 10406
rect 15842 7032 15898 7041
rect 15842 6967 15898 6976
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15672 3862 15792 3890
rect 15580 3726 15700 3754
rect 15474 3703 15530 3712
rect 15384 3674 15436 3680
rect 15396 3618 15424 3674
rect 14922 2751 14978 2760
rect 14476 1414 14596 1442
rect 14660 1550 14872 1578
rect 15028 2746 15240 2774
rect 15304 3590 15424 3618
rect 14476 800 14504 1414
rect 14660 1306 14688 1550
rect 14740 1488 14792 1494
rect 15028 1442 15056 2746
rect 15198 2680 15254 2689
rect 15198 2615 15254 2624
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 14740 1430 14792 1436
rect 14568 1278 14688 1306
rect 14568 800 14596 1278
rect 14752 800 14780 1430
rect 14844 1414 15056 1442
rect 14844 800 14872 1414
rect 15016 1352 15068 1358
rect 15016 1294 15068 1300
rect 15028 800 15056 1294
rect 15120 800 15148 2314
rect 15212 1306 15240 2615
rect 15304 1442 15332 3590
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 2582 15424 3470
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 15304 1414 15424 1442
rect 15212 1278 15332 1306
rect 15304 800 15332 1278
rect 15396 800 15424 1414
rect 15488 1170 15516 2790
rect 15672 1358 15700 3726
rect 15764 1494 15792 3862
rect 15752 1488 15804 1494
rect 15752 1430 15804 1436
rect 15660 1352 15712 1358
rect 15660 1294 15712 1300
rect 15660 1216 15712 1222
rect 15488 1142 15608 1170
rect 15660 1158 15712 1164
rect 15580 800 15608 1142
rect 15672 800 15700 1158
rect 15856 800 15884 6802
rect 15948 3534 15976 13126
rect 16040 4758 16068 14554
rect 16304 13864 16356 13870
rect 16302 13832 16304 13841
rect 16356 13832 16358 13841
rect 16302 13767 16358 13776
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 12850 16344 13194
rect 16408 13190 16436 18838
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16132 12238 16160 12650
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 12073 16160 12174
rect 16118 12064 16174 12073
rect 16118 11999 16174 12008
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 6866 16160 10406
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16224 9489 16252 10134
rect 16210 9480 16266 9489
rect 16210 9415 16266 9424
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16118 6760 16174 6769
rect 16118 6695 16174 6704
rect 16132 6322 16160 6695
rect 16224 6338 16252 9318
rect 16316 8566 16344 12786
rect 16500 12434 16528 14214
rect 16408 12406 16528 12434
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16302 8392 16358 8401
rect 16302 8327 16358 8336
rect 16316 6458 16344 8327
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16120 6316 16172 6322
rect 16224 6310 16344 6338
rect 16120 6258 16172 6264
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15934 3088 15990 3097
rect 15934 3023 15990 3032
rect 15948 2990 15976 3023
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16040 800 16068 3946
rect 16132 2854 16160 6258
rect 16316 6254 16344 6310
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16224 4865 16252 6190
rect 16210 4856 16266 4865
rect 16210 4791 16266 4800
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16210 4040 16266 4049
rect 16210 3975 16266 3984
rect 16224 2990 16252 3975
rect 16316 2990 16344 4626
rect 16408 3670 16436 12406
rect 16592 12374 16620 24890
rect 16776 13190 16804 32370
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 8022 16528 11494
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 5778 16528 7686
rect 16592 6866 16620 9862
rect 16684 7410 16712 11018
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16592 5710 16620 6054
rect 16580 5704 16632 5710
rect 16578 5672 16580 5681
rect 16632 5672 16634 5681
rect 16578 5607 16634 5616
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16500 4185 16528 4762
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16684 4282 16712 4558
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16486 4176 16542 4185
rect 16486 4111 16542 4120
rect 16592 4060 16620 4218
rect 16500 4032 16620 4060
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16210 2816 16266 2825
rect 16210 2751 16266 2760
rect 16224 1442 16252 2751
rect 16316 2650 16344 2926
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16120 1420 16172 1426
rect 16224 1414 16344 1442
rect 16120 1362 16172 1368
rect 16132 800 16160 1362
rect 16316 800 16344 1414
rect 16408 800 16436 2858
rect 16500 1222 16528 4032
rect 16578 3632 16634 3641
rect 16578 3567 16634 3576
rect 16672 3596 16724 3602
rect 16592 1902 16620 3567
rect 16672 3538 16724 3544
rect 16580 1896 16632 1902
rect 16580 1838 16632 1844
rect 16580 1420 16632 1426
rect 16580 1362 16632 1368
rect 16488 1216 16540 1222
rect 16488 1158 16540 1164
rect 16592 800 16620 1362
rect 16684 800 16712 3538
rect 16776 2582 16804 13126
rect 16960 12306 16988 41414
rect 17040 38752 17092 38758
rect 17040 38694 17092 38700
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 6322 16896 8774
rect 16960 7886 16988 11494
rect 17052 8634 17080 38694
rect 17144 14618 17172 64942
rect 17776 62688 17828 62694
rect 17776 62630 17828 62636
rect 17224 59560 17276 59566
rect 17224 59502 17276 59508
rect 17236 59430 17264 59502
rect 17224 59424 17276 59430
rect 17224 59366 17276 59372
rect 17236 44946 17264 59366
rect 17224 44940 17276 44946
rect 17224 44882 17276 44888
rect 17684 44940 17736 44946
rect 17684 44882 17736 44888
rect 17696 41682 17724 44882
rect 17684 41676 17736 41682
rect 17684 41618 17736 41624
rect 17500 40928 17552 40934
rect 17500 40870 17552 40876
rect 17512 40730 17540 40870
rect 17500 40724 17552 40730
rect 17500 40666 17552 40672
rect 17512 26234 17540 40666
rect 17684 32360 17736 32366
rect 17684 32302 17736 32308
rect 17420 26206 17540 26234
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17144 13870 17172 14418
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17052 7698 17080 8026
rect 17144 7954 17172 11018
rect 17236 10606 17264 17614
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 14618 17356 15846
rect 17420 15570 17448 26206
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 9081 17264 10542
rect 17222 9072 17278 9081
rect 17222 9007 17278 9016
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17236 8090 17264 8910
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 16960 7670 17080 7698
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16960 6202 16988 7670
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16868 6174 16988 6202
rect 16868 4672 16896 6174
rect 17052 5778 17080 6598
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16868 4644 16988 4672
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 16868 800 16896 4490
rect 16960 800 16988 4644
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 17052 1426 17080 4490
rect 17040 1420 17092 1426
rect 17040 1362 17092 1368
rect 17144 800 17172 7890
rect 17222 5264 17278 5273
rect 17222 5199 17278 5208
rect 17236 4758 17264 5199
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17236 3670 17264 4490
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17328 3602 17356 14554
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17420 4078 17448 14282
rect 17696 14278 17724 32302
rect 17788 17882 17816 62630
rect 17868 50788 17920 50794
rect 17868 50730 17920 50736
rect 17880 44946 17908 50730
rect 17868 44940 17920 44946
rect 17868 44882 17920 44888
rect 17868 44736 17920 44742
rect 17868 44678 17920 44684
rect 17880 43654 17908 44678
rect 17868 43648 17920 43654
rect 17868 43590 17920 43596
rect 17880 43314 17908 43590
rect 17868 43308 17920 43314
rect 17868 43250 17920 43256
rect 17960 41676 18012 41682
rect 17960 41618 18012 41624
rect 17972 40730 18000 41618
rect 17960 40724 18012 40730
rect 17960 40666 18012 40672
rect 17868 30116 17920 30122
rect 17868 30058 17920 30064
rect 17880 29306 17908 30058
rect 17868 29300 17920 29306
rect 17868 29242 17920 29248
rect 17868 25764 17920 25770
rect 17868 25706 17920 25712
rect 17880 24954 17908 25706
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17880 17746 17908 18090
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 18064 16250 18092 66574
rect 19076 65482 19104 66982
rect 19220 66940 19516 66960
rect 19276 66938 19300 66940
rect 19356 66938 19380 66940
rect 19436 66938 19460 66940
rect 19298 66886 19300 66938
rect 19362 66886 19374 66938
rect 19436 66886 19438 66938
rect 19276 66884 19300 66886
rect 19356 66884 19380 66886
rect 19436 66884 19460 66886
rect 19220 66864 19516 66884
rect 24220 66396 24516 66416
rect 24276 66394 24300 66396
rect 24356 66394 24380 66396
rect 24436 66394 24460 66396
rect 24298 66342 24300 66394
rect 24362 66342 24374 66394
rect 24436 66342 24438 66394
rect 24276 66340 24300 66342
rect 24356 66340 24380 66342
rect 24436 66340 24460 66342
rect 24220 66320 24516 66340
rect 19220 65852 19516 65872
rect 19276 65850 19300 65852
rect 19356 65850 19380 65852
rect 19436 65850 19460 65852
rect 19298 65798 19300 65850
rect 19362 65798 19374 65850
rect 19436 65798 19438 65850
rect 19276 65796 19300 65798
rect 19356 65796 19380 65798
rect 19436 65796 19460 65798
rect 19220 65776 19516 65796
rect 19064 65476 19116 65482
rect 19064 65418 19116 65424
rect 23020 65408 23072 65414
rect 23020 65350 23072 65356
rect 23032 65142 23060 65350
rect 24220 65308 24516 65328
rect 24276 65306 24300 65308
rect 24356 65306 24380 65308
rect 24436 65306 24460 65308
rect 24298 65254 24300 65306
rect 24362 65254 24374 65306
rect 24436 65254 24438 65306
rect 24276 65252 24300 65254
rect 24356 65252 24380 65254
rect 24436 65252 24460 65254
rect 24220 65232 24516 65252
rect 23020 65136 23072 65142
rect 23020 65078 23072 65084
rect 19220 64764 19516 64784
rect 19276 64762 19300 64764
rect 19356 64762 19380 64764
rect 19436 64762 19460 64764
rect 19298 64710 19300 64762
rect 19362 64710 19374 64762
rect 19436 64710 19438 64762
rect 19276 64708 19300 64710
rect 19356 64708 19380 64710
rect 19436 64708 19460 64710
rect 19220 64688 19516 64708
rect 24220 64220 24516 64240
rect 24276 64218 24300 64220
rect 24356 64218 24380 64220
rect 24436 64218 24460 64220
rect 24298 64166 24300 64218
rect 24362 64166 24374 64218
rect 24436 64166 24438 64218
rect 24276 64164 24300 64166
rect 24356 64164 24380 64166
rect 24436 64164 24460 64166
rect 24220 64144 24516 64164
rect 19220 63676 19516 63696
rect 19276 63674 19300 63676
rect 19356 63674 19380 63676
rect 19436 63674 19460 63676
rect 19298 63622 19300 63674
rect 19362 63622 19374 63674
rect 19436 63622 19438 63674
rect 19276 63620 19300 63622
rect 19356 63620 19380 63622
rect 19436 63620 19460 63622
rect 19220 63600 19516 63620
rect 24220 63132 24516 63152
rect 24276 63130 24300 63132
rect 24356 63130 24380 63132
rect 24436 63130 24460 63132
rect 24298 63078 24300 63130
rect 24362 63078 24374 63130
rect 24436 63078 24438 63130
rect 24276 63076 24300 63078
rect 24356 63076 24380 63078
rect 24436 63076 24460 63078
rect 24220 63056 24516 63076
rect 19984 63028 20036 63034
rect 19984 62970 20036 62976
rect 19220 62588 19516 62608
rect 19276 62586 19300 62588
rect 19356 62586 19380 62588
rect 19436 62586 19460 62588
rect 19298 62534 19300 62586
rect 19362 62534 19374 62586
rect 19436 62534 19438 62586
rect 19276 62532 19300 62534
rect 19356 62532 19380 62534
rect 19436 62532 19460 62534
rect 19220 62512 19516 62532
rect 19220 61500 19516 61520
rect 19276 61498 19300 61500
rect 19356 61498 19380 61500
rect 19436 61498 19460 61500
rect 19298 61446 19300 61498
rect 19362 61446 19374 61498
rect 19436 61446 19438 61498
rect 19276 61444 19300 61446
rect 19356 61444 19380 61446
rect 19436 61444 19460 61446
rect 19220 61424 19516 61444
rect 19220 60412 19516 60432
rect 19276 60410 19300 60412
rect 19356 60410 19380 60412
rect 19436 60410 19460 60412
rect 19298 60358 19300 60410
rect 19362 60358 19374 60410
rect 19436 60358 19438 60410
rect 19276 60356 19300 60358
rect 19356 60356 19380 60358
rect 19436 60356 19460 60358
rect 19220 60336 19516 60356
rect 19220 59324 19516 59344
rect 19276 59322 19300 59324
rect 19356 59322 19380 59324
rect 19436 59322 19460 59324
rect 19298 59270 19300 59322
rect 19362 59270 19374 59322
rect 19436 59270 19438 59322
rect 19276 59268 19300 59270
rect 19356 59268 19380 59270
rect 19436 59268 19460 59270
rect 19220 59248 19516 59268
rect 19220 58236 19516 58256
rect 19276 58234 19300 58236
rect 19356 58234 19380 58236
rect 19436 58234 19460 58236
rect 19298 58182 19300 58234
rect 19362 58182 19374 58234
rect 19436 58182 19438 58234
rect 19276 58180 19300 58182
rect 19356 58180 19380 58182
rect 19436 58180 19460 58182
rect 19220 58160 19516 58180
rect 18328 57248 18380 57254
rect 18328 57190 18380 57196
rect 18340 42294 18368 57190
rect 19220 57148 19516 57168
rect 19276 57146 19300 57148
rect 19356 57146 19380 57148
rect 19436 57146 19460 57148
rect 19298 57094 19300 57146
rect 19362 57094 19374 57146
rect 19436 57094 19438 57146
rect 19276 57092 19300 57094
rect 19356 57092 19380 57094
rect 19436 57092 19460 57094
rect 19220 57072 19516 57092
rect 19220 56060 19516 56080
rect 19276 56058 19300 56060
rect 19356 56058 19380 56060
rect 19436 56058 19460 56060
rect 19298 56006 19300 56058
rect 19362 56006 19374 56058
rect 19436 56006 19438 56058
rect 19276 56004 19300 56006
rect 19356 56004 19380 56006
rect 19436 56004 19460 56006
rect 19220 55984 19516 56004
rect 19220 54972 19516 54992
rect 19276 54970 19300 54972
rect 19356 54970 19380 54972
rect 19436 54970 19460 54972
rect 19298 54918 19300 54970
rect 19362 54918 19374 54970
rect 19436 54918 19438 54970
rect 19276 54916 19300 54918
rect 19356 54916 19380 54918
rect 19436 54916 19460 54918
rect 19220 54896 19516 54916
rect 19220 53884 19516 53904
rect 19276 53882 19300 53884
rect 19356 53882 19380 53884
rect 19436 53882 19460 53884
rect 19298 53830 19300 53882
rect 19362 53830 19374 53882
rect 19436 53830 19438 53882
rect 19276 53828 19300 53830
rect 19356 53828 19380 53830
rect 19436 53828 19460 53830
rect 19220 53808 19516 53828
rect 19996 53446 20024 62970
rect 24220 62044 24516 62064
rect 24276 62042 24300 62044
rect 24356 62042 24380 62044
rect 24436 62042 24460 62044
rect 24298 61990 24300 62042
rect 24362 61990 24374 62042
rect 24436 61990 24438 62042
rect 24276 61988 24300 61990
rect 24356 61988 24380 61990
rect 24436 61988 24460 61990
rect 24220 61968 24516 61988
rect 24220 60956 24516 60976
rect 24276 60954 24300 60956
rect 24356 60954 24380 60956
rect 24436 60954 24460 60956
rect 24298 60902 24300 60954
rect 24362 60902 24374 60954
rect 24436 60902 24438 60954
rect 24276 60900 24300 60902
rect 24356 60900 24380 60902
rect 24436 60900 24460 60902
rect 24220 60880 24516 60900
rect 24220 59868 24516 59888
rect 24276 59866 24300 59868
rect 24356 59866 24380 59868
rect 24436 59866 24460 59868
rect 24298 59814 24300 59866
rect 24362 59814 24374 59866
rect 24436 59814 24438 59866
rect 24276 59812 24300 59814
rect 24356 59812 24380 59814
rect 24436 59812 24460 59814
rect 24220 59792 24516 59812
rect 24220 58780 24516 58800
rect 24276 58778 24300 58780
rect 24356 58778 24380 58780
rect 24436 58778 24460 58780
rect 24298 58726 24300 58778
rect 24362 58726 24374 58778
rect 24436 58726 24438 58778
rect 24276 58724 24300 58726
rect 24356 58724 24380 58726
rect 24436 58724 24460 58726
rect 24220 58704 24516 58724
rect 24220 57692 24516 57712
rect 24276 57690 24300 57692
rect 24356 57690 24380 57692
rect 24436 57690 24460 57692
rect 24298 57638 24300 57690
rect 24362 57638 24374 57690
rect 24436 57638 24438 57690
rect 24276 57636 24300 57638
rect 24356 57636 24380 57638
rect 24436 57636 24460 57638
rect 24220 57616 24516 57636
rect 25504 57384 25556 57390
rect 25504 57326 25556 57332
rect 24220 56604 24516 56624
rect 24276 56602 24300 56604
rect 24356 56602 24380 56604
rect 24436 56602 24460 56604
rect 24298 56550 24300 56602
rect 24362 56550 24374 56602
rect 24436 56550 24438 56602
rect 24276 56548 24300 56550
rect 24356 56548 24380 56550
rect 24436 56548 24460 56550
rect 24220 56528 24516 56548
rect 25516 55690 25544 57326
rect 25504 55684 25556 55690
rect 25504 55626 25556 55632
rect 24220 55516 24516 55536
rect 24276 55514 24300 55516
rect 24356 55514 24380 55516
rect 24436 55514 24460 55516
rect 24298 55462 24300 55514
rect 24362 55462 24374 55514
rect 24436 55462 24438 55514
rect 24276 55460 24300 55462
rect 24356 55460 24380 55462
rect 24436 55460 24460 55462
rect 24220 55440 24516 55460
rect 24220 54428 24516 54448
rect 24276 54426 24300 54428
rect 24356 54426 24380 54428
rect 24436 54426 24460 54428
rect 24298 54374 24300 54426
rect 24362 54374 24374 54426
rect 24436 54374 24438 54426
rect 24276 54372 24300 54374
rect 24356 54372 24380 54374
rect 24436 54372 24460 54374
rect 24220 54352 24516 54372
rect 19984 53440 20036 53446
rect 19984 53382 20036 53388
rect 19220 52796 19516 52816
rect 19276 52794 19300 52796
rect 19356 52794 19380 52796
rect 19436 52794 19460 52796
rect 19298 52742 19300 52794
rect 19362 52742 19374 52794
rect 19436 52742 19438 52794
rect 19276 52740 19300 52742
rect 19356 52740 19380 52742
rect 19436 52740 19460 52742
rect 19220 52720 19516 52740
rect 19996 52494 20024 53382
rect 24220 53340 24516 53360
rect 24276 53338 24300 53340
rect 24356 53338 24380 53340
rect 24436 53338 24460 53340
rect 24298 53286 24300 53338
rect 24362 53286 24374 53338
rect 24436 53286 24438 53338
rect 24276 53284 24300 53286
rect 24356 53284 24380 53286
rect 24436 53284 24460 53286
rect 24220 53264 24516 53284
rect 19984 52488 20036 52494
rect 19984 52430 20036 52436
rect 20628 52488 20680 52494
rect 20628 52430 20680 52436
rect 19220 51708 19516 51728
rect 19276 51706 19300 51708
rect 19356 51706 19380 51708
rect 19436 51706 19460 51708
rect 19298 51654 19300 51706
rect 19362 51654 19374 51706
rect 19436 51654 19438 51706
rect 19276 51652 19300 51654
rect 19356 51652 19380 51654
rect 19436 51652 19460 51654
rect 19220 51632 19516 51652
rect 19220 50620 19516 50640
rect 19276 50618 19300 50620
rect 19356 50618 19380 50620
rect 19436 50618 19460 50620
rect 19298 50566 19300 50618
rect 19362 50566 19374 50618
rect 19436 50566 19438 50618
rect 19276 50564 19300 50566
rect 19356 50564 19380 50566
rect 19436 50564 19460 50566
rect 19220 50544 19516 50564
rect 19220 49532 19516 49552
rect 19276 49530 19300 49532
rect 19356 49530 19380 49532
rect 19436 49530 19460 49532
rect 19298 49478 19300 49530
rect 19362 49478 19374 49530
rect 19436 49478 19438 49530
rect 19276 49476 19300 49478
rect 19356 49476 19380 49478
rect 19436 49476 19460 49478
rect 19220 49456 19516 49476
rect 19220 48444 19516 48464
rect 19276 48442 19300 48444
rect 19356 48442 19380 48444
rect 19436 48442 19460 48444
rect 19298 48390 19300 48442
rect 19362 48390 19374 48442
rect 19436 48390 19438 48442
rect 19276 48388 19300 48390
rect 19356 48388 19380 48390
rect 19436 48388 19460 48390
rect 19220 48368 19516 48388
rect 19220 47356 19516 47376
rect 19276 47354 19300 47356
rect 19356 47354 19380 47356
rect 19436 47354 19460 47356
rect 19298 47302 19300 47354
rect 19362 47302 19374 47354
rect 19436 47302 19438 47354
rect 19276 47300 19300 47302
rect 19356 47300 19380 47302
rect 19436 47300 19460 47302
rect 19220 47280 19516 47300
rect 19220 46268 19516 46288
rect 19276 46266 19300 46268
rect 19356 46266 19380 46268
rect 19436 46266 19460 46268
rect 19298 46214 19300 46266
rect 19362 46214 19374 46266
rect 19436 46214 19438 46266
rect 19276 46212 19300 46214
rect 19356 46212 19380 46214
rect 19436 46212 19460 46214
rect 19220 46192 19516 46212
rect 19220 45180 19516 45200
rect 19276 45178 19300 45180
rect 19356 45178 19380 45180
rect 19436 45178 19460 45180
rect 19298 45126 19300 45178
rect 19362 45126 19374 45178
rect 19436 45126 19438 45178
rect 19276 45124 19300 45126
rect 19356 45124 19380 45126
rect 19436 45124 19460 45126
rect 19220 45104 19516 45124
rect 19220 44092 19516 44112
rect 19276 44090 19300 44092
rect 19356 44090 19380 44092
rect 19436 44090 19460 44092
rect 19298 44038 19300 44090
rect 19362 44038 19374 44090
rect 19436 44038 19438 44090
rect 19276 44036 19300 44038
rect 19356 44036 19380 44038
rect 19436 44036 19460 44038
rect 19220 44016 19516 44036
rect 19220 43004 19516 43024
rect 19276 43002 19300 43004
rect 19356 43002 19380 43004
rect 19436 43002 19460 43004
rect 19298 42950 19300 43002
rect 19362 42950 19374 43002
rect 19436 42950 19438 43002
rect 19276 42948 19300 42950
rect 19356 42948 19380 42950
rect 19436 42948 19460 42950
rect 19220 42928 19516 42948
rect 18328 42288 18380 42294
rect 18328 42230 18380 42236
rect 18340 41834 18368 42230
rect 19220 41916 19516 41936
rect 19276 41914 19300 41916
rect 19356 41914 19380 41916
rect 19436 41914 19460 41916
rect 19298 41862 19300 41914
rect 19362 41862 19374 41914
rect 19436 41862 19438 41914
rect 19276 41860 19300 41862
rect 19356 41860 19380 41862
rect 19436 41860 19460 41862
rect 19220 41840 19516 41860
rect 18156 41806 18368 41834
rect 18156 41682 18184 41806
rect 18144 41676 18196 41682
rect 18144 41618 18196 41624
rect 18604 41676 18656 41682
rect 18604 41618 18656 41624
rect 18616 40934 18644 41618
rect 18604 40928 18656 40934
rect 18604 40870 18656 40876
rect 19220 40828 19516 40848
rect 19276 40826 19300 40828
rect 19356 40826 19380 40828
rect 19436 40826 19460 40828
rect 19298 40774 19300 40826
rect 19362 40774 19374 40826
rect 19436 40774 19438 40826
rect 19276 40772 19300 40774
rect 19356 40772 19380 40774
rect 19436 40772 19460 40774
rect 19220 40752 19516 40772
rect 19220 39740 19516 39760
rect 19276 39738 19300 39740
rect 19356 39738 19380 39740
rect 19436 39738 19460 39740
rect 19298 39686 19300 39738
rect 19362 39686 19374 39738
rect 19436 39686 19438 39738
rect 19276 39684 19300 39686
rect 19356 39684 19380 39686
rect 19436 39684 19460 39686
rect 19220 39664 19516 39684
rect 19220 38652 19516 38672
rect 19276 38650 19300 38652
rect 19356 38650 19380 38652
rect 19436 38650 19460 38652
rect 19298 38598 19300 38650
rect 19362 38598 19374 38650
rect 19436 38598 19438 38650
rect 19276 38596 19300 38598
rect 19356 38596 19380 38598
rect 19436 38596 19460 38598
rect 19220 38576 19516 38596
rect 19220 37564 19516 37584
rect 19276 37562 19300 37564
rect 19356 37562 19380 37564
rect 19436 37562 19460 37564
rect 19298 37510 19300 37562
rect 19362 37510 19374 37562
rect 19436 37510 19438 37562
rect 19276 37508 19300 37510
rect 19356 37508 19380 37510
rect 19436 37508 19460 37510
rect 19220 37488 19516 37508
rect 19220 36476 19516 36496
rect 19276 36474 19300 36476
rect 19356 36474 19380 36476
rect 19436 36474 19460 36476
rect 19298 36422 19300 36474
rect 19362 36422 19374 36474
rect 19436 36422 19438 36474
rect 19276 36420 19300 36422
rect 19356 36420 19380 36422
rect 19436 36420 19460 36422
rect 19220 36400 19516 36420
rect 19220 35388 19516 35408
rect 19276 35386 19300 35388
rect 19356 35386 19380 35388
rect 19436 35386 19460 35388
rect 19298 35334 19300 35386
rect 19362 35334 19374 35386
rect 19436 35334 19438 35386
rect 19276 35332 19300 35334
rect 19356 35332 19380 35334
rect 19436 35332 19460 35334
rect 19220 35312 19516 35332
rect 19220 34300 19516 34320
rect 19276 34298 19300 34300
rect 19356 34298 19380 34300
rect 19436 34298 19460 34300
rect 19298 34246 19300 34298
rect 19362 34246 19374 34298
rect 19436 34246 19438 34298
rect 19276 34244 19300 34246
rect 19356 34244 19380 34246
rect 19436 34244 19460 34246
rect 19220 34224 19516 34244
rect 19220 33212 19516 33232
rect 19276 33210 19300 33212
rect 19356 33210 19380 33212
rect 19436 33210 19460 33212
rect 19298 33158 19300 33210
rect 19362 33158 19374 33210
rect 19436 33158 19438 33210
rect 19276 33156 19300 33158
rect 19356 33156 19380 33158
rect 19436 33156 19460 33158
rect 19220 33136 19516 33156
rect 19220 32124 19516 32144
rect 19276 32122 19300 32124
rect 19356 32122 19380 32124
rect 19436 32122 19460 32124
rect 19298 32070 19300 32122
rect 19362 32070 19374 32122
rect 19436 32070 19438 32122
rect 19276 32068 19300 32070
rect 19356 32068 19380 32070
rect 19436 32068 19460 32070
rect 19220 32048 19516 32068
rect 19220 31036 19516 31056
rect 19276 31034 19300 31036
rect 19356 31034 19380 31036
rect 19436 31034 19460 31036
rect 19298 30982 19300 31034
rect 19362 30982 19374 31034
rect 19436 30982 19438 31034
rect 19276 30980 19300 30982
rect 19356 30980 19380 30982
rect 19436 30980 19460 30982
rect 19220 30960 19516 30980
rect 19220 29948 19516 29968
rect 19276 29946 19300 29948
rect 19356 29946 19380 29948
rect 19436 29946 19460 29948
rect 19298 29894 19300 29946
rect 19362 29894 19374 29946
rect 19436 29894 19438 29946
rect 19276 29892 19300 29894
rect 19356 29892 19380 29894
rect 19436 29892 19460 29894
rect 19220 29872 19516 29892
rect 19220 28860 19516 28880
rect 19276 28858 19300 28860
rect 19356 28858 19380 28860
rect 19436 28858 19460 28860
rect 19298 28806 19300 28858
rect 19362 28806 19374 28858
rect 19436 28806 19438 28858
rect 19276 28804 19300 28806
rect 19356 28804 19380 28806
rect 19436 28804 19460 28806
rect 19220 28784 19516 28804
rect 19220 27772 19516 27792
rect 19276 27770 19300 27772
rect 19356 27770 19380 27772
rect 19436 27770 19460 27772
rect 19298 27718 19300 27770
rect 19362 27718 19374 27770
rect 19436 27718 19438 27770
rect 19276 27716 19300 27718
rect 19356 27716 19380 27718
rect 19436 27716 19460 27718
rect 19220 27696 19516 27716
rect 18236 27532 18288 27538
rect 18236 27474 18288 27480
rect 18248 26790 18276 27474
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18236 26784 18288 26790
rect 18236 26726 18288 26732
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18248 18426 18276 19450
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18248 17814 18276 18362
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17604 13870 17632 14010
rect 17972 13954 18000 14214
rect 18064 14074 18092 14486
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17972 13926 18092 13954
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17498 12336 17554 12345
rect 17498 12271 17554 12280
rect 17512 10810 17540 12271
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17512 8922 17540 9454
rect 17604 9042 17632 12582
rect 18064 12434 18092 13926
rect 18156 12986 18184 17478
rect 18340 16574 18368 18702
rect 18340 16546 18460 16574
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17972 12406 18092 12434
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17512 8894 17632 8922
rect 17498 8800 17554 8809
rect 17498 8735 17554 8744
rect 17512 6610 17540 8735
rect 17604 6866 17632 8894
rect 17696 8362 17724 11494
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17696 7154 17724 7414
rect 17788 7274 17816 11018
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17696 7126 17816 7154
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 6730 17632 6802
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17512 6582 17632 6610
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17512 3890 17540 4966
rect 17604 4554 17632 6582
rect 17684 5092 17736 5098
rect 17684 5034 17736 5040
rect 17592 4548 17644 4554
rect 17592 4490 17644 4496
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17420 3862 17540 3890
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17224 2100 17276 2106
rect 17224 2042 17276 2048
rect 17236 800 17264 2042
rect 17420 800 17448 3862
rect 17498 3496 17554 3505
rect 17498 3431 17554 3440
rect 17512 2990 17540 3431
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 1170 17540 2790
rect 17604 2310 17632 4014
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17604 1766 17632 2246
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 17512 1142 17632 1170
rect 17604 800 17632 1142
rect 17696 800 17724 5034
rect 17788 2774 17816 7126
rect 17880 5166 17908 9114
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17972 3670 18000 12406
rect 18156 12322 18184 12922
rect 18064 12294 18184 12322
rect 18248 12306 18276 15302
rect 18432 13190 18460 16546
rect 18524 14890 18552 27270
rect 18800 27130 18828 27406
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 19220 26684 19516 26704
rect 19276 26682 19300 26684
rect 19356 26682 19380 26684
rect 19436 26682 19460 26684
rect 19298 26630 19300 26682
rect 19362 26630 19374 26682
rect 19436 26630 19438 26682
rect 19276 26628 19300 26630
rect 19356 26628 19380 26630
rect 19436 26628 19460 26630
rect 19220 26608 19516 26628
rect 19220 25596 19516 25616
rect 19276 25594 19300 25596
rect 19356 25594 19380 25596
rect 19436 25594 19460 25596
rect 19298 25542 19300 25594
rect 19362 25542 19374 25594
rect 19436 25542 19438 25594
rect 19276 25540 19300 25542
rect 19356 25540 19380 25542
rect 19436 25540 19460 25542
rect 19220 25520 19516 25540
rect 19220 24508 19516 24528
rect 19276 24506 19300 24508
rect 19356 24506 19380 24508
rect 19436 24506 19460 24508
rect 19298 24454 19300 24506
rect 19362 24454 19374 24506
rect 19436 24454 19438 24506
rect 19276 24452 19300 24454
rect 19356 24452 19380 24454
rect 19436 24452 19460 24454
rect 19220 24432 19516 24452
rect 20640 24274 20668 52430
rect 24220 52252 24516 52272
rect 24276 52250 24300 52252
rect 24356 52250 24380 52252
rect 24436 52250 24460 52252
rect 24298 52198 24300 52250
rect 24362 52198 24374 52250
rect 24436 52198 24438 52250
rect 24276 52196 24300 52198
rect 24356 52196 24380 52198
rect 24436 52196 24460 52198
rect 24220 52176 24516 52196
rect 24220 51164 24516 51184
rect 24276 51162 24300 51164
rect 24356 51162 24380 51164
rect 24436 51162 24460 51164
rect 24298 51110 24300 51162
rect 24362 51110 24374 51162
rect 24436 51110 24438 51162
rect 24276 51108 24300 51110
rect 24356 51108 24380 51110
rect 24436 51108 24460 51110
rect 24220 51088 24516 51108
rect 23296 50176 23348 50182
rect 23296 50118 23348 50124
rect 23308 49978 23336 50118
rect 24220 50076 24516 50096
rect 24276 50074 24300 50076
rect 24356 50074 24380 50076
rect 24436 50074 24460 50076
rect 24298 50022 24300 50074
rect 24362 50022 24374 50074
rect 24436 50022 24438 50074
rect 24276 50020 24300 50022
rect 24356 50020 24380 50022
rect 24436 50020 24460 50022
rect 24220 50000 24516 50020
rect 23296 49972 23348 49978
rect 23296 49914 23348 49920
rect 24220 48988 24516 49008
rect 24276 48986 24300 48988
rect 24356 48986 24380 48988
rect 24436 48986 24460 48988
rect 24298 48934 24300 48986
rect 24362 48934 24374 48986
rect 24436 48934 24438 48986
rect 24276 48932 24300 48934
rect 24356 48932 24380 48934
rect 24436 48932 24460 48934
rect 24220 48912 24516 48932
rect 24220 47900 24516 47920
rect 24276 47898 24300 47900
rect 24356 47898 24380 47900
rect 24436 47898 24460 47900
rect 24298 47846 24300 47898
rect 24362 47846 24374 47898
rect 24436 47846 24438 47898
rect 24276 47844 24300 47846
rect 24356 47844 24380 47846
rect 24436 47844 24460 47846
rect 24220 47824 24516 47844
rect 24220 46812 24516 46832
rect 24276 46810 24300 46812
rect 24356 46810 24380 46812
rect 24436 46810 24460 46812
rect 24298 46758 24300 46810
rect 24362 46758 24374 46810
rect 24436 46758 24438 46810
rect 24276 46756 24300 46758
rect 24356 46756 24380 46758
rect 24436 46756 24460 46758
rect 24220 46736 24516 46756
rect 24220 45724 24516 45744
rect 24276 45722 24300 45724
rect 24356 45722 24380 45724
rect 24436 45722 24460 45724
rect 24298 45670 24300 45722
rect 24362 45670 24374 45722
rect 24436 45670 24438 45722
rect 24276 45668 24300 45670
rect 24356 45668 24380 45670
rect 24436 45668 24460 45670
rect 24220 45648 24516 45668
rect 21364 45008 21416 45014
rect 21364 44950 21416 44956
rect 21376 44402 21404 44950
rect 24220 44636 24516 44656
rect 24276 44634 24300 44636
rect 24356 44634 24380 44636
rect 24436 44634 24460 44636
rect 24298 44582 24300 44634
rect 24362 44582 24374 44634
rect 24436 44582 24438 44634
rect 24276 44580 24300 44582
rect 24356 44580 24380 44582
rect 24436 44580 24460 44582
rect 24220 44560 24516 44580
rect 21364 44396 21416 44402
rect 21364 44338 21416 44344
rect 24220 43548 24516 43568
rect 24276 43546 24300 43548
rect 24356 43546 24380 43548
rect 24436 43546 24460 43548
rect 24298 43494 24300 43546
rect 24362 43494 24374 43546
rect 24436 43494 24438 43546
rect 24276 43492 24300 43494
rect 24356 43492 24380 43494
rect 24436 43492 24460 43494
rect 24220 43472 24516 43492
rect 24220 42460 24516 42480
rect 24276 42458 24300 42460
rect 24356 42458 24380 42460
rect 24436 42458 24460 42460
rect 24298 42406 24300 42458
rect 24362 42406 24374 42458
rect 24436 42406 24438 42458
rect 24276 42404 24300 42406
rect 24356 42404 24380 42406
rect 24436 42404 24460 42406
rect 24220 42384 24516 42404
rect 22928 42288 22980 42294
rect 22928 42230 22980 42236
rect 22940 42090 22968 42230
rect 22928 42084 22980 42090
rect 22928 42026 22980 42032
rect 21364 42016 21416 42022
rect 21364 41958 21416 41964
rect 21376 41750 21404 41958
rect 21364 41744 21416 41750
rect 21364 41686 21416 41692
rect 22940 40594 22968 42026
rect 24220 41372 24516 41392
rect 24276 41370 24300 41372
rect 24356 41370 24380 41372
rect 24436 41370 24460 41372
rect 24298 41318 24300 41370
rect 24362 41318 24374 41370
rect 24436 41318 24438 41370
rect 24276 41316 24300 41318
rect 24356 41316 24380 41318
rect 24436 41316 24460 41318
rect 24220 41296 24516 41316
rect 22928 40588 22980 40594
rect 22928 40530 22980 40536
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 21008 29306 21036 29446
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 19220 23420 19516 23440
rect 19276 23418 19300 23420
rect 19356 23418 19380 23420
rect 19436 23418 19460 23420
rect 19298 23366 19300 23418
rect 19362 23366 19374 23418
rect 19436 23366 19438 23418
rect 19276 23364 19300 23366
rect 19356 23364 19380 23366
rect 19436 23364 19460 23366
rect 19220 23344 19516 23364
rect 19220 22332 19516 22352
rect 19276 22330 19300 22332
rect 19356 22330 19380 22332
rect 19436 22330 19460 22332
rect 19298 22278 19300 22330
rect 19362 22278 19374 22330
rect 19436 22278 19438 22330
rect 19276 22276 19300 22278
rect 19356 22276 19380 22278
rect 19436 22276 19460 22278
rect 19220 22256 19516 22276
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18236 12300 18288 12306
rect 18064 12238 18092 12294
rect 18236 12242 18288 12248
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 8430 18092 11494
rect 18326 11248 18382 11257
rect 18326 11183 18382 11192
rect 18234 10840 18290 10849
rect 18234 10775 18236 10784
rect 18288 10775 18290 10784
rect 18236 10746 18288 10752
rect 18340 10130 18368 11183
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17880 2922 17908 3538
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 2990 18000 3334
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 18064 2774 18092 8366
rect 18156 6866 18184 9862
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 7954 18276 9318
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18236 7336 18288 7342
rect 18340 7324 18368 9930
rect 18288 7296 18368 7324
rect 18236 7278 18288 7284
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 4146 18184 5510
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18248 3738 18276 7278
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 17788 2746 17908 2774
rect 17880 800 17908 2746
rect 17972 2746 18092 2774
rect 17972 800 18000 2746
rect 18156 800 18184 3674
rect 18340 2825 18368 4218
rect 18326 2816 18382 2825
rect 18326 2751 18382 2760
rect 18326 2680 18382 2689
rect 18326 2615 18382 2624
rect 18340 1442 18368 2615
rect 18432 2582 18460 13126
rect 18524 4622 18552 14826
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18616 3890 18644 13806
rect 18708 4078 18736 14418
rect 18800 6361 18828 14758
rect 18892 9654 18920 22034
rect 19220 21244 19516 21264
rect 19276 21242 19300 21244
rect 19356 21242 19380 21244
rect 19436 21242 19460 21244
rect 19298 21190 19300 21242
rect 19362 21190 19374 21242
rect 19436 21190 19438 21242
rect 19276 21188 19300 21190
rect 19356 21188 19380 21190
rect 19436 21188 19460 21190
rect 19220 21168 19516 21188
rect 19220 20156 19516 20176
rect 19276 20154 19300 20156
rect 19356 20154 19380 20156
rect 19436 20154 19460 20156
rect 19298 20102 19300 20154
rect 19362 20102 19374 20154
rect 19436 20102 19438 20154
rect 19276 20100 19300 20102
rect 19356 20100 19380 20102
rect 19436 20100 19460 20102
rect 19220 20080 19516 20100
rect 19996 12782 20024 24210
rect 22940 23186 22968 40530
rect 23020 40384 23072 40390
rect 23020 40326 23072 40332
rect 23032 28762 23060 40326
rect 24220 40284 24516 40304
rect 24276 40282 24300 40284
rect 24356 40282 24380 40284
rect 24436 40282 24460 40284
rect 24298 40230 24300 40282
rect 24362 40230 24374 40282
rect 24436 40230 24438 40282
rect 24276 40228 24300 40230
rect 24356 40228 24380 40230
rect 24436 40228 24460 40230
rect 24220 40208 24516 40228
rect 24220 39196 24516 39216
rect 24276 39194 24300 39196
rect 24356 39194 24380 39196
rect 24436 39194 24460 39196
rect 24298 39142 24300 39194
rect 24362 39142 24374 39194
rect 24436 39142 24438 39194
rect 24276 39140 24300 39142
rect 24356 39140 24380 39142
rect 24436 39140 24460 39142
rect 24220 39120 24516 39140
rect 24220 38108 24516 38128
rect 24276 38106 24300 38108
rect 24356 38106 24380 38108
rect 24436 38106 24460 38108
rect 24298 38054 24300 38106
rect 24362 38054 24374 38106
rect 24436 38054 24438 38106
rect 24276 38052 24300 38054
rect 24356 38052 24380 38054
rect 24436 38052 24460 38054
rect 24220 38032 24516 38052
rect 24220 37020 24516 37040
rect 24276 37018 24300 37020
rect 24356 37018 24380 37020
rect 24436 37018 24460 37020
rect 24298 36966 24300 37018
rect 24362 36966 24374 37018
rect 24436 36966 24438 37018
rect 24276 36964 24300 36966
rect 24356 36964 24380 36966
rect 24436 36964 24460 36966
rect 24220 36944 24516 36964
rect 24220 35932 24516 35952
rect 24276 35930 24300 35932
rect 24356 35930 24380 35932
rect 24436 35930 24460 35932
rect 24298 35878 24300 35930
rect 24362 35878 24374 35930
rect 24436 35878 24438 35930
rect 24276 35876 24300 35878
rect 24356 35876 24380 35878
rect 24436 35876 24460 35878
rect 24220 35856 24516 35876
rect 24220 34844 24516 34864
rect 24276 34842 24300 34844
rect 24356 34842 24380 34844
rect 24436 34842 24460 34844
rect 24298 34790 24300 34842
rect 24362 34790 24374 34842
rect 24436 34790 24438 34842
rect 24276 34788 24300 34790
rect 24356 34788 24380 34790
rect 24436 34788 24460 34790
rect 24220 34768 24516 34788
rect 24220 33756 24516 33776
rect 24276 33754 24300 33756
rect 24356 33754 24380 33756
rect 24436 33754 24460 33756
rect 24298 33702 24300 33754
rect 24362 33702 24374 33754
rect 24436 33702 24438 33754
rect 24276 33700 24300 33702
rect 24356 33700 24380 33702
rect 24436 33700 24460 33702
rect 24220 33680 24516 33700
rect 24220 32668 24516 32688
rect 24276 32666 24300 32668
rect 24356 32666 24380 32668
rect 24436 32666 24460 32668
rect 24298 32614 24300 32666
rect 24362 32614 24374 32666
rect 24436 32614 24438 32666
rect 24276 32612 24300 32614
rect 24356 32612 24380 32614
rect 24436 32612 24460 32614
rect 24220 32592 24516 32612
rect 24220 31580 24516 31600
rect 24276 31578 24300 31580
rect 24356 31578 24380 31580
rect 24436 31578 24460 31580
rect 24298 31526 24300 31578
rect 24362 31526 24374 31578
rect 24436 31526 24438 31578
rect 24276 31524 24300 31526
rect 24356 31524 24380 31526
rect 24436 31524 24460 31526
rect 24220 31504 24516 31524
rect 25228 30592 25280 30598
rect 25228 30534 25280 30540
rect 24220 30492 24516 30512
rect 24276 30490 24300 30492
rect 24356 30490 24380 30492
rect 24436 30490 24460 30492
rect 24298 30438 24300 30490
rect 24362 30438 24374 30490
rect 24436 30438 24438 30490
rect 24276 30436 24300 30438
rect 24356 30436 24380 30438
rect 24436 30436 24460 30438
rect 24220 30416 24516 30436
rect 24220 29404 24516 29424
rect 24276 29402 24300 29404
rect 24356 29402 24380 29404
rect 24436 29402 24460 29404
rect 24298 29350 24300 29402
rect 24362 29350 24374 29402
rect 24436 29350 24438 29402
rect 24276 29348 24300 29350
rect 24356 29348 24380 29350
rect 24436 29348 24460 29350
rect 24220 29328 24516 29348
rect 23020 28756 23072 28762
rect 23020 28698 23072 28704
rect 24220 28316 24516 28336
rect 24276 28314 24300 28316
rect 24356 28314 24380 28316
rect 24436 28314 24460 28316
rect 24298 28262 24300 28314
rect 24362 28262 24374 28314
rect 24436 28262 24438 28314
rect 24276 28260 24300 28262
rect 24356 28260 24380 28262
rect 24436 28260 24460 28262
rect 24220 28240 24516 28260
rect 24220 27228 24516 27248
rect 24276 27226 24300 27228
rect 24356 27226 24380 27228
rect 24436 27226 24460 27228
rect 24298 27174 24300 27226
rect 24362 27174 24374 27226
rect 24436 27174 24438 27226
rect 24276 27172 24300 27174
rect 24356 27172 24380 27174
rect 24436 27172 24460 27174
rect 24220 27152 24516 27172
rect 25240 27130 25268 30534
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 24220 26140 24516 26160
rect 24276 26138 24300 26140
rect 24356 26138 24380 26140
rect 24436 26138 24460 26140
rect 24298 26086 24300 26138
rect 24362 26086 24374 26138
rect 24436 26086 24438 26138
rect 24276 26084 24300 26086
rect 24356 26084 24380 26086
rect 24436 26084 24460 26086
rect 24220 26064 24516 26084
rect 24220 25052 24516 25072
rect 24276 25050 24300 25052
rect 24356 25050 24380 25052
rect 24436 25050 24460 25052
rect 24298 24998 24300 25050
rect 24362 24998 24374 25050
rect 24436 24998 24438 25050
rect 24276 24996 24300 24998
rect 24356 24996 24380 24998
rect 24436 24996 24460 24998
rect 24220 24976 24516 24996
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23492 24410 23520 24754
rect 23480 24404 23532 24410
rect 23480 24346 23532 24352
rect 24220 23964 24516 23984
rect 24276 23962 24300 23964
rect 24356 23962 24380 23964
rect 24436 23962 24460 23964
rect 24298 23910 24300 23962
rect 24362 23910 24374 23962
rect 24436 23910 24438 23962
rect 24276 23908 24300 23910
rect 24356 23908 24380 23910
rect 24436 23908 24460 23910
rect 24220 23888 24516 23908
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22940 22094 22968 23122
rect 24220 22876 24516 22896
rect 24276 22874 24300 22876
rect 24356 22874 24380 22876
rect 24436 22874 24460 22876
rect 24298 22822 24300 22874
rect 24362 22822 24374 22874
rect 24436 22822 24438 22874
rect 24276 22820 24300 22822
rect 24356 22820 24380 22822
rect 24436 22820 24460 22822
rect 24220 22800 24516 22820
rect 22940 22066 23336 22094
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22112 17241 22140 21830
rect 22098 17232 22154 17241
rect 22098 17167 22154 17176
rect 23308 12850 23336 22066
rect 24220 21788 24516 21808
rect 24276 21786 24300 21788
rect 24356 21786 24380 21788
rect 24436 21786 24460 21788
rect 24298 21734 24300 21786
rect 24362 21734 24374 21786
rect 24436 21734 24438 21786
rect 24276 21732 24300 21734
rect 24356 21732 24380 21734
rect 24436 21732 24460 21734
rect 24220 21712 24516 21732
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 23952 12442 23980 21490
rect 25608 21486 25636 66982
rect 26884 66632 26936 66638
rect 26884 66574 26936 66580
rect 26332 48204 26384 48210
rect 26332 48146 26384 48152
rect 26344 29510 26372 48146
rect 26896 31890 26924 66574
rect 26988 57866 27016 67118
rect 34152 67108 34204 67114
rect 34152 67050 34204 67056
rect 41512 67108 41564 67114
rect 41512 67050 41564 67056
rect 47768 67108 47820 67114
rect 47768 67050 47820 67056
rect 57796 67108 57848 67114
rect 57796 67050 57848 67056
rect 33232 67040 33284 67046
rect 33232 66982 33284 66988
rect 29220 66940 29516 66960
rect 29276 66938 29300 66940
rect 29356 66938 29380 66940
rect 29436 66938 29460 66940
rect 29298 66886 29300 66938
rect 29362 66886 29374 66938
rect 29436 66886 29438 66938
rect 29276 66884 29300 66886
rect 29356 66884 29380 66886
rect 29436 66884 29460 66886
rect 29220 66864 29516 66884
rect 30472 66496 30524 66502
rect 30472 66438 30524 66444
rect 30288 66088 30340 66094
rect 30288 66030 30340 66036
rect 30196 65952 30248 65958
rect 30196 65894 30248 65900
rect 29220 65852 29516 65872
rect 29276 65850 29300 65852
rect 29356 65850 29380 65852
rect 29436 65850 29460 65852
rect 29298 65798 29300 65850
rect 29362 65798 29374 65850
rect 29436 65798 29438 65850
rect 29276 65796 29300 65798
rect 29356 65796 29380 65798
rect 29436 65796 29460 65798
rect 29220 65776 29516 65796
rect 30208 65754 30236 65894
rect 30300 65754 30328 66030
rect 30196 65748 30248 65754
rect 30196 65690 30248 65696
rect 30288 65748 30340 65754
rect 30288 65690 30340 65696
rect 29220 64764 29516 64784
rect 29276 64762 29300 64764
rect 29356 64762 29380 64764
rect 29436 64762 29460 64764
rect 29298 64710 29300 64762
rect 29362 64710 29374 64762
rect 29436 64710 29438 64762
rect 29276 64708 29300 64710
rect 29356 64708 29380 64710
rect 29436 64708 29460 64710
rect 29220 64688 29516 64708
rect 27528 64388 27580 64394
rect 27528 64330 27580 64336
rect 27540 63578 27568 64330
rect 29220 63676 29516 63696
rect 29276 63674 29300 63676
rect 29356 63674 29380 63676
rect 29436 63674 29460 63676
rect 29298 63622 29300 63674
rect 29362 63622 29374 63674
rect 29436 63622 29438 63674
rect 29276 63620 29300 63622
rect 29356 63620 29380 63622
rect 29436 63620 29460 63622
rect 29220 63600 29516 63620
rect 27528 63572 27580 63578
rect 27528 63514 27580 63520
rect 26976 57860 27028 57866
rect 26976 57802 27028 57808
rect 27540 48210 27568 63514
rect 29220 62588 29516 62608
rect 29276 62586 29300 62588
rect 29356 62586 29380 62588
rect 29436 62586 29460 62588
rect 29298 62534 29300 62586
rect 29362 62534 29374 62586
rect 29436 62534 29438 62586
rect 29276 62532 29300 62534
rect 29356 62532 29380 62534
rect 29436 62532 29460 62534
rect 29220 62512 29516 62532
rect 29220 61500 29516 61520
rect 29276 61498 29300 61500
rect 29356 61498 29380 61500
rect 29436 61498 29460 61500
rect 29298 61446 29300 61498
rect 29362 61446 29374 61498
rect 29436 61446 29438 61498
rect 29276 61444 29300 61446
rect 29356 61444 29380 61446
rect 29436 61444 29460 61446
rect 29220 61424 29516 61444
rect 29220 60412 29516 60432
rect 29276 60410 29300 60412
rect 29356 60410 29380 60412
rect 29436 60410 29460 60412
rect 29298 60358 29300 60410
rect 29362 60358 29374 60410
rect 29436 60358 29438 60410
rect 29276 60356 29300 60358
rect 29356 60356 29380 60358
rect 29436 60356 29460 60358
rect 29220 60336 29516 60356
rect 30288 60036 30340 60042
rect 30288 59978 30340 59984
rect 29220 59324 29516 59344
rect 29276 59322 29300 59324
rect 29356 59322 29380 59324
rect 29436 59322 29460 59324
rect 29298 59270 29300 59322
rect 29362 59270 29374 59322
rect 29436 59270 29438 59322
rect 29276 59268 29300 59270
rect 29356 59268 29380 59270
rect 29436 59268 29460 59270
rect 29220 59248 29516 59268
rect 30300 58682 30328 59978
rect 29092 58676 29144 58682
rect 29092 58618 29144 58624
rect 30288 58676 30340 58682
rect 30288 58618 30340 58624
rect 27988 58472 28040 58478
rect 27988 58414 28040 58420
rect 28000 58002 28028 58414
rect 27988 57996 28040 58002
rect 27988 57938 28040 57944
rect 27804 57792 27856 57798
rect 27804 57734 27856 57740
rect 27528 48204 27580 48210
rect 27528 48146 27580 48152
rect 27540 47258 27568 48146
rect 27528 47252 27580 47258
rect 27528 47194 27580 47200
rect 27252 42900 27304 42906
rect 27252 42842 27304 42848
rect 26884 31884 26936 31890
rect 26884 31826 26936 31832
rect 26884 29708 26936 29714
rect 26884 29650 26936 29656
rect 26332 29504 26384 29510
rect 26332 29446 26384 29452
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26160 22642 26188 27066
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 24220 20700 24516 20720
rect 24276 20698 24300 20700
rect 24356 20698 24380 20700
rect 24436 20698 24460 20700
rect 24298 20646 24300 20698
rect 24362 20646 24374 20698
rect 24436 20646 24438 20698
rect 24276 20644 24300 20646
rect 24356 20644 24380 20646
rect 24436 20644 24460 20646
rect 24220 20624 24516 20644
rect 24220 19612 24516 19632
rect 24276 19610 24300 19612
rect 24356 19610 24380 19612
rect 24436 19610 24460 19612
rect 24298 19558 24300 19610
rect 24362 19558 24374 19610
rect 24436 19558 24438 19610
rect 24276 19556 24300 19558
rect 24356 19556 24380 19558
rect 24436 19556 24460 19558
rect 24220 19536 24516 19556
rect 26344 18970 26372 29446
rect 26896 29238 26924 29650
rect 26884 29232 26936 29238
rect 26884 29174 26936 29180
rect 27264 20058 27292 42842
rect 27620 30184 27672 30190
rect 27620 30126 27672 30132
rect 27344 27056 27396 27062
rect 27344 26998 27396 27004
rect 27356 26314 27384 26998
rect 27344 26308 27396 26314
rect 27344 26250 27396 26256
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 27632 16590 27660 30126
rect 27816 20602 27844 57734
rect 29104 53582 29132 58618
rect 29220 58236 29516 58256
rect 29276 58234 29300 58236
rect 29356 58234 29380 58236
rect 29436 58234 29460 58236
rect 29298 58182 29300 58234
rect 29362 58182 29374 58234
rect 29436 58182 29438 58234
rect 29276 58180 29300 58182
rect 29356 58180 29380 58182
rect 29436 58180 29460 58182
rect 29220 58160 29516 58180
rect 29220 57148 29516 57168
rect 29276 57146 29300 57148
rect 29356 57146 29380 57148
rect 29436 57146 29460 57148
rect 29298 57094 29300 57146
rect 29362 57094 29374 57146
rect 29436 57094 29438 57146
rect 29276 57092 29300 57094
rect 29356 57092 29380 57094
rect 29436 57092 29460 57094
rect 29220 57072 29516 57092
rect 30288 56296 30340 56302
rect 30288 56238 30340 56244
rect 29220 56060 29516 56080
rect 29276 56058 29300 56060
rect 29356 56058 29380 56060
rect 29436 56058 29460 56060
rect 29298 56006 29300 56058
rect 29362 56006 29374 56058
rect 29436 56006 29438 56058
rect 29276 56004 29300 56006
rect 29356 56004 29380 56006
rect 29436 56004 29460 56006
rect 29220 55984 29516 56004
rect 29220 54972 29516 54992
rect 29276 54970 29300 54972
rect 29356 54970 29380 54972
rect 29436 54970 29460 54972
rect 29298 54918 29300 54970
rect 29362 54918 29374 54970
rect 29436 54918 29438 54970
rect 29276 54916 29300 54918
rect 29356 54916 29380 54918
rect 29436 54916 29460 54918
rect 29220 54896 29516 54916
rect 29220 53884 29516 53904
rect 29276 53882 29300 53884
rect 29356 53882 29380 53884
rect 29436 53882 29460 53884
rect 29298 53830 29300 53882
rect 29362 53830 29374 53882
rect 29436 53830 29438 53882
rect 29276 53828 29300 53830
rect 29356 53828 29380 53830
rect 29436 53828 29460 53830
rect 29220 53808 29516 53828
rect 29092 53576 29144 53582
rect 29092 53518 29144 53524
rect 29552 53576 29604 53582
rect 29552 53518 29604 53524
rect 29220 52796 29516 52816
rect 29276 52794 29300 52796
rect 29356 52794 29380 52796
rect 29436 52794 29460 52796
rect 29298 52742 29300 52794
rect 29362 52742 29374 52794
rect 29436 52742 29438 52794
rect 29276 52740 29300 52742
rect 29356 52740 29380 52742
rect 29436 52740 29460 52742
rect 29220 52720 29516 52740
rect 29220 51708 29516 51728
rect 29276 51706 29300 51708
rect 29356 51706 29380 51708
rect 29436 51706 29460 51708
rect 29298 51654 29300 51706
rect 29362 51654 29374 51706
rect 29436 51654 29438 51706
rect 29276 51652 29300 51654
rect 29356 51652 29380 51654
rect 29436 51652 29460 51654
rect 29220 51632 29516 51652
rect 29220 50620 29516 50640
rect 29276 50618 29300 50620
rect 29356 50618 29380 50620
rect 29436 50618 29460 50620
rect 29298 50566 29300 50618
rect 29362 50566 29374 50618
rect 29436 50566 29438 50618
rect 29276 50564 29300 50566
rect 29356 50564 29380 50566
rect 29436 50564 29460 50566
rect 29220 50544 29516 50564
rect 28264 49632 28316 49638
rect 28264 49574 28316 49580
rect 28276 41546 28304 49574
rect 29220 49532 29516 49552
rect 29276 49530 29300 49532
rect 29356 49530 29380 49532
rect 29436 49530 29460 49532
rect 29298 49478 29300 49530
rect 29362 49478 29374 49530
rect 29436 49478 29438 49530
rect 29276 49476 29300 49478
rect 29356 49476 29380 49478
rect 29436 49476 29460 49478
rect 29220 49456 29516 49476
rect 29220 48444 29516 48464
rect 29276 48442 29300 48444
rect 29356 48442 29380 48444
rect 29436 48442 29460 48444
rect 29298 48390 29300 48442
rect 29362 48390 29374 48442
rect 29436 48390 29438 48442
rect 29276 48388 29300 48390
rect 29356 48388 29380 48390
rect 29436 48388 29460 48390
rect 29220 48368 29516 48388
rect 29220 47356 29516 47376
rect 29276 47354 29300 47356
rect 29356 47354 29380 47356
rect 29436 47354 29460 47356
rect 29298 47302 29300 47354
rect 29362 47302 29374 47354
rect 29436 47302 29438 47354
rect 29276 47300 29300 47302
rect 29356 47300 29380 47302
rect 29436 47300 29460 47302
rect 29220 47280 29516 47300
rect 29220 46268 29516 46288
rect 29276 46266 29300 46268
rect 29356 46266 29380 46268
rect 29436 46266 29460 46268
rect 29298 46214 29300 46266
rect 29362 46214 29374 46266
rect 29436 46214 29438 46266
rect 29276 46212 29300 46214
rect 29356 46212 29380 46214
rect 29436 46212 29460 46214
rect 29220 46192 29516 46212
rect 29220 45180 29516 45200
rect 29276 45178 29300 45180
rect 29356 45178 29380 45180
rect 29436 45178 29460 45180
rect 29298 45126 29300 45178
rect 29362 45126 29374 45178
rect 29436 45126 29438 45178
rect 29276 45124 29300 45126
rect 29356 45124 29380 45126
rect 29436 45124 29460 45126
rect 29220 45104 29516 45124
rect 29220 44092 29516 44112
rect 29276 44090 29300 44092
rect 29356 44090 29380 44092
rect 29436 44090 29460 44092
rect 29298 44038 29300 44090
rect 29362 44038 29374 44090
rect 29436 44038 29438 44090
rect 29276 44036 29300 44038
rect 29356 44036 29380 44038
rect 29436 44036 29460 44038
rect 29220 44016 29516 44036
rect 29220 43004 29516 43024
rect 29276 43002 29300 43004
rect 29356 43002 29380 43004
rect 29436 43002 29460 43004
rect 29298 42950 29300 43002
rect 29362 42950 29374 43002
rect 29436 42950 29438 43002
rect 29276 42948 29300 42950
rect 29356 42948 29380 42950
rect 29436 42948 29460 42950
rect 29220 42928 29516 42948
rect 29220 41916 29516 41936
rect 29276 41914 29300 41916
rect 29356 41914 29380 41916
rect 29436 41914 29460 41916
rect 29298 41862 29300 41914
rect 29362 41862 29374 41914
rect 29436 41862 29438 41914
rect 29276 41860 29300 41862
rect 29356 41860 29380 41862
rect 29436 41860 29460 41862
rect 29220 41840 29516 41860
rect 28264 41540 28316 41546
rect 28264 41482 28316 41488
rect 28448 41540 28500 41546
rect 28448 41482 28500 41488
rect 27896 26852 27948 26858
rect 27896 26794 27948 26800
rect 27908 26518 27936 26794
rect 28172 26580 28224 26586
rect 28172 26522 28224 26528
rect 27896 26512 27948 26518
rect 27896 26454 27948 26460
rect 28184 26450 28212 26522
rect 28460 26450 28488 41482
rect 29220 40828 29516 40848
rect 29276 40826 29300 40828
rect 29356 40826 29380 40828
rect 29436 40826 29460 40828
rect 29298 40774 29300 40826
rect 29362 40774 29374 40826
rect 29436 40774 29438 40826
rect 29276 40772 29300 40774
rect 29356 40772 29380 40774
rect 29436 40772 29460 40774
rect 29220 40752 29516 40772
rect 29220 39740 29516 39760
rect 29276 39738 29300 39740
rect 29356 39738 29380 39740
rect 29436 39738 29460 39740
rect 29298 39686 29300 39738
rect 29362 39686 29374 39738
rect 29436 39686 29438 39738
rect 29276 39684 29300 39686
rect 29356 39684 29380 39686
rect 29436 39684 29460 39686
rect 29220 39664 29516 39684
rect 29000 39296 29052 39302
rect 29000 39238 29052 39244
rect 29012 37942 29040 39238
rect 29220 38652 29516 38672
rect 29276 38650 29300 38652
rect 29356 38650 29380 38652
rect 29436 38650 29460 38652
rect 29298 38598 29300 38650
rect 29362 38598 29374 38650
rect 29436 38598 29438 38650
rect 29276 38596 29300 38598
rect 29356 38596 29380 38598
rect 29436 38596 29460 38598
rect 29220 38576 29516 38596
rect 29000 37936 29052 37942
rect 29000 37878 29052 37884
rect 29220 37564 29516 37584
rect 29276 37562 29300 37564
rect 29356 37562 29380 37564
rect 29436 37562 29460 37564
rect 29298 37510 29300 37562
rect 29362 37510 29374 37562
rect 29436 37510 29438 37562
rect 29276 37508 29300 37510
rect 29356 37508 29380 37510
rect 29436 37508 29460 37510
rect 29220 37488 29516 37508
rect 29220 36476 29516 36496
rect 29276 36474 29300 36476
rect 29356 36474 29380 36476
rect 29436 36474 29460 36476
rect 29298 36422 29300 36474
rect 29362 36422 29374 36474
rect 29436 36422 29438 36474
rect 29276 36420 29300 36422
rect 29356 36420 29380 36422
rect 29436 36420 29460 36422
rect 29220 36400 29516 36420
rect 29220 35388 29516 35408
rect 29276 35386 29300 35388
rect 29356 35386 29380 35388
rect 29436 35386 29460 35388
rect 29298 35334 29300 35386
rect 29362 35334 29374 35386
rect 29436 35334 29438 35386
rect 29276 35332 29300 35334
rect 29356 35332 29380 35334
rect 29436 35332 29460 35334
rect 29220 35312 29516 35332
rect 29220 34300 29516 34320
rect 29276 34298 29300 34300
rect 29356 34298 29380 34300
rect 29436 34298 29460 34300
rect 29298 34246 29300 34298
rect 29362 34246 29374 34298
rect 29436 34246 29438 34298
rect 29276 34244 29300 34246
rect 29356 34244 29380 34246
rect 29436 34244 29460 34246
rect 29220 34224 29516 34244
rect 29220 33212 29516 33232
rect 29276 33210 29300 33212
rect 29356 33210 29380 33212
rect 29436 33210 29460 33212
rect 29298 33158 29300 33210
rect 29362 33158 29374 33210
rect 29436 33158 29438 33210
rect 29276 33156 29300 33158
rect 29356 33156 29380 33158
rect 29436 33156 29460 33158
rect 29220 33136 29516 33156
rect 29220 32124 29516 32144
rect 29276 32122 29300 32124
rect 29356 32122 29380 32124
rect 29436 32122 29460 32124
rect 29298 32070 29300 32122
rect 29362 32070 29374 32122
rect 29436 32070 29438 32122
rect 29276 32068 29300 32070
rect 29356 32068 29380 32070
rect 29436 32068 29460 32070
rect 29220 32048 29516 32068
rect 29220 31036 29516 31056
rect 29276 31034 29300 31036
rect 29356 31034 29380 31036
rect 29436 31034 29460 31036
rect 29298 30982 29300 31034
rect 29362 30982 29374 31034
rect 29436 30982 29438 31034
rect 29276 30980 29300 30982
rect 29356 30980 29380 30982
rect 29436 30980 29460 30982
rect 29220 30960 29516 30980
rect 29220 29948 29516 29968
rect 29276 29946 29300 29948
rect 29356 29946 29380 29948
rect 29436 29946 29460 29948
rect 29298 29894 29300 29946
rect 29362 29894 29374 29946
rect 29436 29894 29438 29946
rect 29276 29892 29300 29894
rect 29356 29892 29380 29894
rect 29436 29892 29460 29894
rect 29220 29872 29516 29892
rect 28540 29844 28592 29850
rect 28540 29786 28592 29792
rect 28552 29646 28580 29786
rect 29564 29782 29592 53518
rect 30300 45014 30328 56238
rect 30288 45008 30340 45014
rect 30288 44950 30340 44956
rect 30484 32434 30512 66438
rect 32404 63232 32456 63238
rect 32404 63174 32456 63180
rect 31300 55888 31352 55894
rect 31300 55830 31352 55836
rect 31312 55350 31340 55830
rect 31300 55344 31352 55350
rect 31300 55286 31352 55292
rect 31312 55214 31340 55286
rect 31312 55186 31432 55214
rect 31300 51808 31352 51814
rect 31300 51750 31352 51756
rect 31312 51406 31340 51750
rect 31300 51400 31352 51406
rect 31300 51342 31352 51348
rect 30932 50380 30984 50386
rect 30932 50322 30984 50328
rect 30944 49910 30972 50322
rect 30932 49904 30984 49910
rect 30932 49846 30984 49852
rect 30564 43852 30616 43858
rect 30564 43794 30616 43800
rect 30576 34950 30604 43794
rect 30748 43648 30800 43654
rect 30748 43590 30800 43596
rect 30760 41750 30788 43590
rect 30748 41744 30800 41750
rect 30748 41686 30800 41692
rect 30564 34944 30616 34950
rect 30564 34886 30616 34892
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30576 30938 30604 34886
rect 30564 30932 30616 30938
rect 30564 30874 30616 30880
rect 29552 29776 29604 29782
rect 29552 29718 29604 29724
rect 28540 29640 28592 29646
rect 28540 29582 28592 29588
rect 29220 28860 29516 28880
rect 29276 28858 29300 28860
rect 29356 28858 29380 28860
rect 29436 28858 29460 28860
rect 29298 28806 29300 28858
rect 29362 28806 29374 28858
rect 29436 28806 29438 28858
rect 29276 28804 29300 28806
rect 29356 28804 29380 28806
rect 29436 28804 29460 28806
rect 29220 28784 29516 28804
rect 30944 28082 30972 49846
rect 31404 41750 31432 55186
rect 32036 51808 32088 51814
rect 32036 51750 32088 51756
rect 31668 47184 31720 47190
rect 31852 47184 31904 47190
rect 31720 47132 31852 47138
rect 31668 47126 31904 47132
rect 31680 47110 31892 47126
rect 31392 41744 31444 41750
rect 31392 41686 31444 41692
rect 32048 34678 32076 51750
rect 32036 34672 32088 34678
rect 32036 34614 32088 34620
rect 32048 34474 32076 34614
rect 31760 34468 31812 34474
rect 31760 34410 31812 34416
rect 32036 34468 32088 34474
rect 32036 34410 32088 34416
rect 31772 31482 31800 34410
rect 31760 31476 31812 31482
rect 31760 31418 31812 31424
rect 31772 28914 31800 31418
rect 32416 30054 32444 63174
rect 32496 62280 32548 62286
rect 32496 62222 32548 62228
rect 32508 34202 32536 62222
rect 33140 62212 33192 62218
rect 33140 62154 33192 62160
rect 33152 58954 33180 62154
rect 33140 58948 33192 58954
rect 33140 58890 33192 58896
rect 32864 53576 32916 53582
rect 32864 53518 32916 53524
rect 33140 53576 33192 53582
rect 33140 53518 33192 53524
rect 32876 52970 32904 53518
rect 32864 52964 32916 52970
rect 32864 52906 32916 52912
rect 32588 46980 32640 46986
rect 32588 46922 32640 46928
rect 32496 34196 32548 34202
rect 32496 34138 32548 34144
rect 32404 30048 32456 30054
rect 32404 29990 32456 29996
rect 31588 28886 31800 28914
rect 31484 28756 31536 28762
rect 31484 28698 31536 28704
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 31392 28076 31444 28082
rect 31392 28018 31444 28024
rect 29220 27772 29516 27792
rect 29276 27770 29300 27772
rect 29356 27770 29380 27772
rect 29436 27770 29460 27772
rect 29298 27718 29300 27770
rect 29362 27718 29374 27770
rect 29436 27718 29438 27770
rect 29276 27716 29300 27718
rect 29356 27716 29380 27718
rect 29436 27716 29460 27718
rect 29220 27696 29516 27716
rect 30196 27668 30248 27674
rect 30196 27610 30248 27616
rect 29220 26684 29516 26704
rect 29276 26682 29300 26684
rect 29356 26682 29380 26684
rect 29436 26682 29460 26684
rect 29298 26630 29300 26682
rect 29362 26630 29374 26682
rect 29436 26630 29438 26682
rect 29276 26628 29300 26630
rect 29356 26628 29380 26630
rect 29436 26628 29460 26630
rect 29220 26608 29516 26628
rect 30208 26586 30236 27610
rect 31116 27328 31168 27334
rect 31116 27270 31168 27276
rect 30196 26580 30248 26586
rect 30196 26522 30248 26528
rect 30208 26450 30236 26522
rect 28172 26444 28224 26450
rect 28172 26386 28224 26392
rect 28448 26444 28500 26450
rect 28448 26386 28500 26392
rect 30196 26444 30248 26450
rect 30196 26386 30248 26392
rect 28460 26042 28488 26386
rect 28448 26036 28500 26042
rect 28448 25978 28500 25984
rect 29220 25596 29516 25616
rect 29276 25594 29300 25596
rect 29356 25594 29380 25596
rect 29436 25594 29460 25596
rect 29298 25542 29300 25594
rect 29362 25542 29374 25594
rect 29436 25542 29438 25594
rect 29276 25540 29300 25542
rect 29356 25540 29380 25542
rect 29436 25540 29460 25542
rect 29220 25520 29516 25540
rect 29220 24508 29516 24528
rect 29276 24506 29300 24508
rect 29356 24506 29380 24508
rect 29436 24506 29460 24508
rect 29298 24454 29300 24506
rect 29362 24454 29374 24506
rect 29436 24454 29438 24506
rect 29276 24452 29300 24454
rect 29356 24452 29380 24454
rect 29436 24452 29460 24454
rect 29220 24432 29516 24452
rect 29092 24064 29144 24070
rect 29092 24006 29144 24012
rect 29104 23798 29132 24006
rect 29092 23792 29144 23798
rect 29092 23734 29144 23740
rect 29220 23420 29516 23440
rect 29276 23418 29300 23420
rect 29356 23418 29380 23420
rect 29436 23418 29460 23420
rect 29298 23366 29300 23418
rect 29362 23366 29374 23418
rect 29436 23366 29438 23418
rect 29276 23364 29300 23366
rect 29356 23364 29380 23366
rect 29436 23364 29460 23366
rect 29220 23344 29516 23364
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 29920 22976 29972 22982
rect 29920 22918 29972 22924
rect 29932 22710 29960 22918
rect 29920 22704 29972 22710
rect 29920 22646 29972 22652
rect 29932 22438 29960 22646
rect 30116 22506 30144 23054
rect 30104 22500 30156 22506
rect 30104 22442 30156 22448
rect 29920 22432 29972 22438
rect 29920 22374 29972 22380
rect 29220 22332 29516 22352
rect 29276 22330 29300 22332
rect 29356 22330 29380 22332
rect 29436 22330 29460 22332
rect 29298 22278 29300 22330
rect 29362 22278 29374 22330
rect 29436 22278 29438 22330
rect 29276 22276 29300 22278
rect 29356 22276 29380 22278
rect 29436 22276 29460 22278
rect 29220 22256 29516 22276
rect 30116 22234 30144 22442
rect 30104 22228 30156 22234
rect 30104 22170 30156 22176
rect 30208 22094 30236 26386
rect 30116 22066 30236 22094
rect 29220 21244 29516 21264
rect 29276 21242 29300 21244
rect 29356 21242 29380 21244
rect 29436 21242 29460 21244
rect 29298 21190 29300 21242
rect 29362 21190 29374 21242
rect 29436 21190 29438 21242
rect 29276 21188 29300 21190
rect 29356 21188 29380 21190
rect 29436 21188 29460 21190
rect 29220 21168 29516 21188
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27816 19854 27844 20538
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 28276 19514 28304 19654
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 29012 17678 29040 20334
rect 29220 20156 29516 20176
rect 29276 20154 29300 20156
rect 29356 20154 29380 20156
rect 29436 20154 29460 20156
rect 29298 20102 29300 20154
rect 29362 20102 29374 20154
rect 29436 20102 29438 20154
rect 29276 20100 29300 20102
rect 29356 20100 29380 20102
rect 29436 20100 29460 20102
rect 29220 20080 29516 20100
rect 30116 20058 30144 22066
rect 31128 20602 31156 27270
rect 31404 26450 31432 28018
rect 31496 28014 31524 28698
rect 31484 28008 31536 28014
rect 31484 27950 31536 27956
rect 31588 27946 31616 28886
rect 31760 28416 31812 28422
rect 31760 28358 31812 28364
rect 31772 28218 31800 28358
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31668 28144 31720 28150
rect 32036 28144 32088 28150
rect 31864 28104 32036 28132
rect 31864 28098 31892 28104
rect 31720 28092 31892 28098
rect 31668 28086 31892 28092
rect 32036 28086 32088 28092
rect 31680 28070 31892 28086
rect 32036 28008 32088 28014
rect 32088 27968 32260 27996
rect 32036 27950 32088 27956
rect 31576 27940 31628 27946
rect 31576 27882 31628 27888
rect 31588 27334 31616 27882
rect 32232 27878 32260 27968
rect 32220 27872 32272 27878
rect 32220 27814 32272 27820
rect 31576 27328 31628 27334
rect 31576 27270 31628 27276
rect 31392 26444 31444 26450
rect 31392 26386 31444 26392
rect 31668 26444 31720 26450
rect 31668 26386 31720 26392
rect 31576 22772 31628 22778
rect 31576 22714 31628 22720
rect 31588 22506 31616 22714
rect 31576 22500 31628 22506
rect 31576 22442 31628 22448
rect 31116 20596 31168 20602
rect 31116 20538 31168 20544
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 31128 19786 31156 20538
rect 31116 19780 31168 19786
rect 31116 19722 31168 19728
rect 31680 19718 31708 26386
rect 32416 22094 32444 29990
rect 32600 26994 32628 46922
rect 32770 34640 32826 34649
rect 32770 34575 32772 34584
rect 32824 34575 32826 34584
rect 32772 34546 32824 34552
rect 32876 30122 32904 52906
rect 33152 52902 33180 53518
rect 33140 52896 33192 52902
rect 33140 52838 33192 52844
rect 33152 44198 33180 52838
rect 33244 47666 33272 66982
rect 34164 66842 34192 67050
rect 36544 67040 36596 67046
rect 36544 66982 36596 66988
rect 34152 66836 34204 66842
rect 34152 66778 34204 66784
rect 34220 66396 34516 66416
rect 34276 66394 34300 66396
rect 34356 66394 34380 66396
rect 34436 66394 34460 66396
rect 34298 66342 34300 66394
rect 34362 66342 34374 66394
rect 34436 66342 34438 66394
rect 34276 66340 34300 66342
rect 34356 66340 34380 66342
rect 34436 66340 34460 66342
rect 34220 66320 34516 66340
rect 36176 66088 36228 66094
rect 36176 66030 36228 66036
rect 36452 66088 36504 66094
rect 36452 66030 36504 66036
rect 36188 65958 36216 66030
rect 34888 65952 34940 65958
rect 34888 65894 34940 65900
rect 36176 65952 36228 65958
rect 36176 65894 36228 65900
rect 34220 65308 34516 65328
rect 34276 65306 34300 65308
rect 34356 65306 34380 65308
rect 34436 65306 34460 65308
rect 34298 65254 34300 65306
rect 34362 65254 34374 65306
rect 34436 65254 34438 65306
rect 34276 65252 34300 65254
rect 34356 65252 34380 65254
rect 34436 65252 34460 65254
rect 34220 65232 34516 65252
rect 34220 64220 34516 64240
rect 34276 64218 34300 64220
rect 34356 64218 34380 64220
rect 34436 64218 34460 64220
rect 34298 64166 34300 64218
rect 34362 64166 34374 64218
rect 34436 64166 34438 64218
rect 34276 64164 34300 64166
rect 34356 64164 34380 64166
rect 34436 64164 34460 64166
rect 34220 64144 34516 64164
rect 34220 63132 34516 63152
rect 34276 63130 34300 63132
rect 34356 63130 34380 63132
rect 34436 63130 34460 63132
rect 34298 63078 34300 63130
rect 34362 63078 34374 63130
rect 34436 63078 34438 63130
rect 34276 63076 34300 63078
rect 34356 63076 34380 63078
rect 34436 63076 34460 63078
rect 34220 63056 34516 63076
rect 34220 62044 34516 62064
rect 34276 62042 34300 62044
rect 34356 62042 34380 62044
rect 34436 62042 34460 62044
rect 34298 61990 34300 62042
rect 34362 61990 34374 62042
rect 34436 61990 34438 62042
rect 34276 61988 34300 61990
rect 34356 61988 34380 61990
rect 34436 61988 34460 61990
rect 34220 61968 34516 61988
rect 34220 60956 34516 60976
rect 34276 60954 34300 60956
rect 34356 60954 34380 60956
rect 34436 60954 34460 60956
rect 34298 60902 34300 60954
rect 34362 60902 34374 60954
rect 34436 60902 34438 60954
rect 34276 60900 34300 60902
rect 34356 60900 34380 60902
rect 34436 60900 34460 60902
rect 34220 60880 34516 60900
rect 34220 59868 34516 59888
rect 34276 59866 34300 59868
rect 34356 59866 34380 59868
rect 34436 59866 34460 59868
rect 34298 59814 34300 59866
rect 34362 59814 34374 59866
rect 34436 59814 34438 59866
rect 34276 59812 34300 59814
rect 34356 59812 34380 59814
rect 34436 59812 34460 59814
rect 34220 59792 34516 59812
rect 33508 59492 33560 59498
rect 33508 59434 33560 59440
rect 33416 58948 33468 58954
rect 33416 58890 33468 58896
rect 33232 47660 33284 47666
rect 33232 47602 33284 47608
rect 33140 44192 33192 44198
rect 33140 44134 33192 44140
rect 33152 43110 33180 44134
rect 33140 43104 33192 43110
rect 33140 43046 33192 43052
rect 33152 39030 33180 43046
rect 33428 39302 33456 58890
rect 33416 39296 33468 39302
rect 33416 39238 33468 39244
rect 33140 39024 33192 39030
rect 33140 38966 33192 38972
rect 33520 38654 33548 59434
rect 34220 58780 34516 58800
rect 34276 58778 34300 58780
rect 34356 58778 34380 58780
rect 34436 58778 34460 58780
rect 34298 58726 34300 58778
rect 34362 58726 34374 58778
rect 34436 58726 34438 58778
rect 34276 58724 34300 58726
rect 34356 58724 34380 58726
rect 34436 58724 34460 58726
rect 34220 58704 34516 58724
rect 34520 58472 34572 58478
rect 34520 58414 34572 58420
rect 34532 58138 34560 58414
rect 34520 58132 34572 58138
rect 34520 58074 34572 58080
rect 34220 57692 34516 57712
rect 34276 57690 34300 57692
rect 34356 57690 34380 57692
rect 34436 57690 34460 57692
rect 34298 57638 34300 57690
rect 34362 57638 34374 57690
rect 34436 57638 34438 57690
rect 34276 57636 34300 57638
rect 34356 57636 34380 57638
rect 34436 57636 34460 57638
rect 34220 57616 34516 57636
rect 34220 56604 34516 56624
rect 34276 56602 34300 56604
rect 34356 56602 34380 56604
rect 34436 56602 34460 56604
rect 34298 56550 34300 56602
rect 34362 56550 34374 56602
rect 34436 56550 34438 56602
rect 34276 56548 34300 56550
rect 34356 56548 34380 56550
rect 34436 56548 34460 56550
rect 34220 56528 34516 56548
rect 34220 55516 34516 55536
rect 34276 55514 34300 55516
rect 34356 55514 34380 55516
rect 34436 55514 34460 55516
rect 34298 55462 34300 55514
rect 34362 55462 34374 55514
rect 34436 55462 34438 55514
rect 34276 55460 34300 55462
rect 34356 55460 34380 55462
rect 34436 55460 34460 55462
rect 34220 55440 34516 55460
rect 33876 54528 33928 54534
rect 33876 54470 33928 54476
rect 33888 49842 33916 54470
rect 34220 54428 34516 54448
rect 34276 54426 34300 54428
rect 34356 54426 34380 54428
rect 34436 54426 34460 54428
rect 34298 54374 34300 54426
rect 34362 54374 34374 54426
rect 34436 54374 34438 54426
rect 34276 54372 34300 54374
rect 34356 54372 34380 54374
rect 34436 54372 34460 54374
rect 34220 54352 34516 54372
rect 34220 53340 34516 53360
rect 34276 53338 34300 53340
rect 34356 53338 34380 53340
rect 34436 53338 34460 53340
rect 34298 53286 34300 53338
rect 34362 53286 34374 53338
rect 34436 53286 34438 53338
rect 34276 53284 34300 53286
rect 34356 53284 34380 53286
rect 34436 53284 34460 53286
rect 34220 53264 34516 53284
rect 34220 52252 34516 52272
rect 34276 52250 34300 52252
rect 34356 52250 34380 52252
rect 34436 52250 34460 52252
rect 34298 52198 34300 52250
rect 34362 52198 34374 52250
rect 34436 52198 34438 52250
rect 34276 52196 34300 52198
rect 34356 52196 34380 52198
rect 34436 52196 34460 52198
rect 34220 52176 34516 52196
rect 34220 51164 34516 51184
rect 34276 51162 34300 51164
rect 34356 51162 34380 51164
rect 34436 51162 34460 51164
rect 34298 51110 34300 51162
rect 34362 51110 34374 51162
rect 34436 51110 34438 51162
rect 34276 51108 34300 51110
rect 34356 51108 34380 51110
rect 34436 51108 34460 51110
rect 34220 51088 34516 51108
rect 34152 50244 34204 50250
rect 34152 50186 34204 50192
rect 33876 49836 33928 49842
rect 33876 49778 33928 49784
rect 33692 39296 33744 39302
rect 33692 39238 33744 39244
rect 33600 39024 33652 39030
rect 33600 38966 33652 38972
rect 33152 38626 33548 38654
rect 32956 35148 33008 35154
rect 32956 35090 33008 35096
rect 32968 34542 32996 35090
rect 33152 34610 33180 38626
rect 33612 38214 33640 38966
rect 33704 38962 33732 39238
rect 33692 38956 33744 38962
rect 33692 38898 33744 38904
rect 33600 38208 33652 38214
rect 33600 38150 33652 38156
rect 33232 34672 33284 34678
rect 33232 34614 33284 34620
rect 33140 34604 33192 34610
rect 33140 34546 33192 34552
rect 32956 34536 33008 34542
rect 32956 34478 33008 34484
rect 33140 34400 33192 34406
rect 33140 34342 33192 34348
rect 32864 30116 32916 30122
rect 32864 30058 32916 30064
rect 33152 28218 33180 34342
rect 33244 34134 33272 34614
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 33336 34202 33364 34478
rect 33324 34196 33376 34202
rect 33324 34138 33376 34144
rect 33232 34128 33284 34134
rect 33232 34070 33284 34076
rect 33140 28212 33192 28218
rect 33140 28154 33192 28160
rect 33152 27674 33180 28154
rect 33232 27872 33284 27878
rect 33232 27814 33284 27820
rect 33140 27668 33192 27674
rect 33140 27610 33192 27616
rect 32588 26988 32640 26994
rect 32588 26930 32640 26936
rect 32956 26988 33008 26994
rect 32956 26930 33008 26936
rect 32968 26518 32996 26930
rect 32956 26512 33008 26518
rect 32956 26454 33008 26460
rect 31864 22066 32444 22094
rect 31864 19922 31892 22066
rect 32404 19984 32456 19990
rect 32404 19926 32456 19932
rect 31852 19916 31904 19922
rect 31852 19858 31904 19864
rect 31668 19712 31720 19718
rect 31668 19654 31720 19660
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 27620 16584 27672 16590
rect 32416 16574 32444 19926
rect 33244 18970 33272 27814
rect 33612 26586 33640 38150
rect 33704 30598 33732 38898
rect 33888 38654 33916 49778
rect 33968 49700 34020 49706
rect 33968 49642 34020 49648
rect 33980 49094 34008 49642
rect 33968 49088 34020 49094
rect 33968 49030 34020 49036
rect 33980 46986 34008 49030
rect 33968 46980 34020 46986
rect 33968 46922 34020 46928
rect 34164 44946 34192 50186
rect 34220 50076 34516 50096
rect 34276 50074 34300 50076
rect 34356 50074 34380 50076
rect 34436 50074 34460 50076
rect 34298 50022 34300 50074
rect 34362 50022 34374 50074
rect 34436 50022 34438 50074
rect 34276 50020 34300 50022
rect 34356 50020 34380 50022
rect 34436 50020 34460 50022
rect 34220 50000 34516 50020
rect 34704 49768 34756 49774
rect 34704 49710 34756 49716
rect 34220 48988 34516 49008
rect 34276 48986 34300 48988
rect 34356 48986 34380 48988
rect 34436 48986 34460 48988
rect 34298 48934 34300 48986
rect 34362 48934 34374 48986
rect 34436 48934 34438 48986
rect 34276 48932 34300 48934
rect 34356 48932 34380 48934
rect 34436 48932 34460 48934
rect 34220 48912 34516 48932
rect 34220 47900 34516 47920
rect 34276 47898 34300 47900
rect 34356 47898 34380 47900
rect 34436 47898 34460 47900
rect 34298 47846 34300 47898
rect 34362 47846 34374 47898
rect 34436 47846 34438 47898
rect 34276 47844 34300 47846
rect 34356 47844 34380 47846
rect 34436 47844 34460 47846
rect 34220 47824 34516 47844
rect 34220 46812 34516 46832
rect 34276 46810 34300 46812
rect 34356 46810 34380 46812
rect 34436 46810 34460 46812
rect 34298 46758 34300 46810
rect 34362 46758 34374 46810
rect 34436 46758 34438 46810
rect 34276 46756 34300 46758
rect 34356 46756 34380 46758
rect 34436 46756 34460 46758
rect 34220 46736 34516 46756
rect 34220 45724 34516 45744
rect 34276 45722 34300 45724
rect 34356 45722 34380 45724
rect 34436 45722 34460 45724
rect 34298 45670 34300 45722
rect 34362 45670 34374 45722
rect 34436 45670 34438 45722
rect 34276 45668 34300 45670
rect 34356 45668 34380 45670
rect 34436 45668 34460 45670
rect 34220 45648 34516 45668
rect 34152 44940 34204 44946
rect 34152 44882 34204 44888
rect 34220 44636 34516 44656
rect 34276 44634 34300 44636
rect 34356 44634 34380 44636
rect 34436 44634 34460 44636
rect 34298 44582 34300 44634
rect 34362 44582 34374 44634
rect 34436 44582 34438 44634
rect 34276 44580 34300 44582
rect 34356 44580 34380 44582
rect 34436 44580 34460 44582
rect 34220 44560 34516 44580
rect 34220 43548 34516 43568
rect 34276 43546 34300 43548
rect 34356 43546 34380 43548
rect 34436 43546 34460 43548
rect 34298 43494 34300 43546
rect 34362 43494 34374 43546
rect 34436 43494 34438 43546
rect 34276 43492 34300 43494
rect 34356 43492 34380 43494
rect 34436 43492 34460 43494
rect 34220 43472 34516 43492
rect 34220 42460 34516 42480
rect 34276 42458 34300 42460
rect 34356 42458 34380 42460
rect 34436 42458 34460 42460
rect 34298 42406 34300 42458
rect 34362 42406 34374 42458
rect 34436 42406 34438 42458
rect 34276 42404 34300 42406
rect 34356 42404 34380 42406
rect 34436 42404 34460 42406
rect 34220 42384 34516 42404
rect 34220 41372 34516 41392
rect 34276 41370 34300 41372
rect 34356 41370 34380 41372
rect 34436 41370 34460 41372
rect 34298 41318 34300 41370
rect 34362 41318 34374 41370
rect 34436 41318 34438 41370
rect 34276 41316 34300 41318
rect 34356 41316 34380 41318
rect 34436 41316 34460 41318
rect 34220 41296 34516 41316
rect 34220 40284 34516 40304
rect 34276 40282 34300 40284
rect 34356 40282 34380 40284
rect 34436 40282 34460 40284
rect 34298 40230 34300 40282
rect 34362 40230 34374 40282
rect 34436 40230 34438 40282
rect 34276 40228 34300 40230
rect 34356 40228 34380 40230
rect 34436 40228 34460 40230
rect 34220 40208 34516 40228
rect 34220 39196 34516 39216
rect 34276 39194 34300 39196
rect 34356 39194 34380 39196
rect 34436 39194 34460 39196
rect 34298 39142 34300 39194
rect 34362 39142 34374 39194
rect 34436 39142 34438 39194
rect 34276 39140 34300 39142
rect 34356 39140 34380 39142
rect 34436 39140 34460 39142
rect 34220 39120 34516 39140
rect 34716 38826 34744 49710
rect 34704 38820 34756 38826
rect 34704 38762 34756 38768
rect 33796 38626 33916 38654
rect 33796 34134 33824 38626
rect 34220 38108 34516 38128
rect 34276 38106 34300 38108
rect 34356 38106 34380 38108
rect 34436 38106 34460 38108
rect 34298 38054 34300 38106
rect 34362 38054 34374 38106
rect 34436 38054 34438 38106
rect 34276 38052 34300 38054
rect 34356 38052 34380 38054
rect 34436 38052 34460 38054
rect 34220 38032 34516 38052
rect 34220 37020 34516 37040
rect 34276 37018 34300 37020
rect 34356 37018 34380 37020
rect 34436 37018 34460 37020
rect 34298 36966 34300 37018
rect 34362 36966 34374 37018
rect 34436 36966 34438 37018
rect 34276 36964 34300 36966
rect 34356 36964 34380 36966
rect 34436 36964 34460 36966
rect 34220 36944 34516 36964
rect 34220 35932 34516 35952
rect 34276 35930 34300 35932
rect 34356 35930 34380 35932
rect 34436 35930 34460 35932
rect 34298 35878 34300 35930
rect 34362 35878 34374 35930
rect 34436 35878 34438 35930
rect 34276 35876 34300 35878
rect 34356 35876 34380 35878
rect 34436 35876 34460 35878
rect 34220 35856 34516 35876
rect 34220 34844 34516 34864
rect 34276 34842 34300 34844
rect 34356 34842 34380 34844
rect 34436 34842 34460 34844
rect 34298 34790 34300 34842
rect 34362 34790 34374 34842
rect 34436 34790 34438 34842
rect 34276 34788 34300 34790
rect 34356 34788 34380 34790
rect 34436 34788 34460 34790
rect 34220 34768 34516 34788
rect 33874 34640 33930 34649
rect 33874 34575 33876 34584
rect 33928 34575 33930 34584
rect 33876 34546 33928 34552
rect 33784 34128 33836 34134
rect 33784 34070 33836 34076
rect 33796 31958 33824 34070
rect 34220 33756 34516 33776
rect 34276 33754 34300 33756
rect 34356 33754 34380 33756
rect 34436 33754 34460 33756
rect 34298 33702 34300 33754
rect 34362 33702 34374 33754
rect 34436 33702 34438 33754
rect 34276 33700 34300 33702
rect 34356 33700 34380 33702
rect 34436 33700 34460 33702
rect 34220 33680 34516 33700
rect 34220 32668 34516 32688
rect 34276 32666 34300 32668
rect 34356 32666 34380 32668
rect 34436 32666 34460 32668
rect 34298 32614 34300 32666
rect 34362 32614 34374 32666
rect 34436 32614 34438 32666
rect 34276 32612 34300 32614
rect 34356 32612 34380 32614
rect 34436 32612 34460 32614
rect 34220 32592 34516 32612
rect 33784 31952 33836 31958
rect 33784 31894 33836 31900
rect 34220 31580 34516 31600
rect 34276 31578 34300 31580
rect 34356 31578 34380 31580
rect 34436 31578 34460 31580
rect 34298 31526 34300 31578
rect 34362 31526 34374 31578
rect 34436 31526 34438 31578
rect 34276 31524 34300 31526
rect 34356 31524 34380 31526
rect 34436 31524 34460 31526
rect 34220 31504 34516 31524
rect 33692 30592 33744 30598
rect 33692 30534 33744 30540
rect 33600 26580 33652 26586
rect 33600 26522 33652 26528
rect 33612 22982 33640 26522
rect 33704 23118 33732 30534
rect 34220 30492 34516 30512
rect 34276 30490 34300 30492
rect 34356 30490 34380 30492
rect 34436 30490 34460 30492
rect 34298 30438 34300 30490
rect 34362 30438 34374 30490
rect 34436 30438 34438 30490
rect 34276 30436 34300 30438
rect 34356 30436 34380 30438
rect 34436 30436 34460 30438
rect 34220 30416 34516 30436
rect 34220 29404 34516 29424
rect 34276 29402 34300 29404
rect 34356 29402 34380 29404
rect 34436 29402 34460 29404
rect 34298 29350 34300 29402
rect 34362 29350 34374 29402
rect 34436 29350 34438 29402
rect 34276 29348 34300 29350
rect 34356 29348 34380 29350
rect 34436 29348 34460 29350
rect 34220 29328 34516 29348
rect 34220 28316 34516 28336
rect 34276 28314 34300 28316
rect 34356 28314 34380 28316
rect 34436 28314 34460 28316
rect 34298 28262 34300 28314
rect 34362 28262 34374 28314
rect 34436 28262 34438 28314
rect 34276 28260 34300 28262
rect 34356 28260 34380 28262
rect 34436 28260 34460 28262
rect 34220 28240 34516 28260
rect 34220 27228 34516 27248
rect 34276 27226 34300 27228
rect 34356 27226 34380 27228
rect 34436 27226 34460 27228
rect 34298 27174 34300 27226
rect 34362 27174 34374 27226
rect 34436 27174 34438 27226
rect 34276 27172 34300 27174
rect 34356 27172 34380 27174
rect 34436 27172 34460 27174
rect 34220 27152 34516 27172
rect 34220 26140 34516 26160
rect 34276 26138 34300 26140
rect 34356 26138 34380 26140
rect 34436 26138 34460 26140
rect 34298 26086 34300 26138
rect 34362 26086 34374 26138
rect 34436 26086 34438 26138
rect 34276 26084 34300 26086
rect 34356 26084 34380 26086
rect 34436 26084 34460 26086
rect 34220 26064 34516 26084
rect 34220 25052 34516 25072
rect 34276 25050 34300 25052
rect 34356 25050 34380 25052
rect 34436 25050 34460 25052
rect 34298 24998 34300 25050
rect 34362 24998 34374 25050
rect 34436 24998 34438 25050
rect 34276 24996 34300 24998
rect 34356 24996 34380 24998
rect 34436 24996 34460 24998
rect 34220 24976 34516 24996
rect 34220 23964 34516 23984
rect 34276 23962 34300 23964
rect 34356 23962 34380 23964
rect 34436 23962 34460 23964
rect 34298 23910 34300 23962
rect 34362 23910 34374 23962
rect 34436 23910 34438 23962
rect 34276 23908 34300 23910
rect 34356 23908 34380 23910
rect 34436 23908 34460 23910
rect 34220 23888 34516 23908
rect 33692 23112 33744 23118
rect 33692 23054 33744 23060
rect 33600 22976 33652 22982
rect 33600 22918 33652 22924
rect 34220 22876 34516 22896
rect 34276 22874 34300 22876
rect 34356 22874 34380 22876
rect 34436 22874 34460 22876
rect 34298 22822 34300 22874
rect 34362 22822 34374 22874
rect 34436 22822 34438 22874
rect 34276 22820 34300 22822
rect 34356 22820 34380 22822
rect 34436 22820 34460 22822
rect 34220 22800 34516 22820
rect 34716 22094 34744 38762
rect 34796 34944 34848 34950
rect 34796 34886 34848 34892
rect 34808 34406 34836 34886
rect 34796 34400 34848 34406
rect 34796 34342 34848 34348
rect 34900 29238 34928 65894
rect 36464 62966 36492 66030
rect 36452 62960 36504 62966
rect 36452 62902 36504 62908
rect 36176 57792 36228 57798
rect 36176 57734 36228 57740
rect 36188 57526 36216 57734
rect 36176 57520 36228 57526
rect 36176 57462 36228 57468
rect 34980 49904 35032 49910
rect 34980 49846 35032 49852
rect 34888 29232 34940 29238
rect 34888 29174 34940 29180
rect 34992 22778 35020 49846
rect 35716 43648 35768 43654
rect 35716 43590 35768 43596
rect 35072 35012 35124 35018
rect 35072 34954 35124 34960
rect 35084 34678 35112 34954
rect 35072 34672 35124 34678
rect 35072 34614 35124 34620
rect 35084 34542 35112 34614
rect 35072 34536 35124 34542
rect 35072 34478 35124 34484
rect 34980 22772 35032 22778
rect 34980 22714 35032 22720
rect 34624 22066 34744 22094
rect 34220 21788 34516 21808
rect 34276 21786 34300 21788
rect 34356 21786 34380 21788
rect 34436 21786 34460 21788
rect 34298 21734 34300 21786
rect 34362 21734 34374 21786
rect 34436 21734 34438 21786
rect 34276 21732 34300 21734
rect 34356 21732 34380 21734
rect 34436 21732 34460 21734
rect 34220 21712 34516 21732
rect 34220 20700 34516 20720
rect 34276 20698 34300 20700
rect 34356 20698 34380 20700
rect 34436 20698 34460 20700
rect 34298 20646 34300 20698
rect 34362 20646 34374 20698
rect 34436 20646 34438 20698
rect 34276 20644 34300 20646
rect 34356 20644 34380 20646
rect 34436 20644 34460 20646
rect 34220 20624 34516 20644
rect 33968 19712 34020 19718
rect 33968 19654 34020 19660
rect 33232 18964 33284 18970
rect 33232 18906 33284 18912
rect 33980 18902 34008 19654
rect 34220 19612 34516 19632
rect 34276 19610 34300 19612
rect 34356 19610 34380 19612
rect 34436 19610 34460 19612
rect 34298 19558 34300 19610
rect 34362 19558 34374 19610
rect 34436 19558 34438 19610
rect 34276 19556 34300 19558
rect 34356 19556 34380 19558
rect 34436 19556 34460 19558
rect 34220 19536 34516 19556
rect 33968 18896 34020 18902
rect 33968 18838 34020 18844
rect 34624 18154 34652 22066
rect 34612 18148 34664 18154
rect 34612 18090 34664 18096
rect 32416 16546 32812 16574
rect 27620 16526 27672 16532
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32600 13124 32628 15846
rect 23940 12436 23992 12442
rect 32784 12434 32812 16546
rect 35728 14346 35756 43590
rect 36452 35148 36504 35154
rect 36452 35090 36504 35096
rect 36464 34678 36492 35090
rect 36452 34672 36504 34678
rect 36452 34614 36504 34620
rect 36452 30728 36504 30734
rect 36452 30670 36504 30676
rect 36464 30394 36492 30670
rect 36452 30388 36504 30394
rect 36452 30330 36504 30336
rect 36556 24274 36584 66982
rect 39220 66940 39516 66960
rect 39276 66938 39300 66940
rect 39356 66938 39380 66940
rect 39436 66938 39460 66940
rect 39298 66886 39300 66938
rect 39362 66886 39374 66938
rect 39436 66886 39438 66938
rect 39276 66884 39300 66886
rect 39356 66884 39380 66886
rect 39436 66884 39460 66886
rect 39220 66864 39516 66884
rect 41524 66502 41552 67050
rect 47780 66842 47808 67050
rect 50804 67040 50856 67046
rect 50804 66982 50856 66988
rect 54760 67040 54812 67046
rect 54760 66982 54812 66988
rect 49220 66940 49516 66960
rect 49276 66938 49300 66940
rect 49356 66938 49380 66940
rect 49436 66938 49460 66940
rect 49298 66886 49300 66938
rect 49362 66886 49374 66938
rect 49436 66886 49438 66938
rect 49276 66884 49300 66886
rect 49356 66884 49380 66886
rect 49436 66884 49460 66886
rect 49220 66864 49516 66884
rect 47768 66836 47820 66842
rect 47768 66778 47820 66784
rect 41512 66496 41564 66502
rect 41512 66438 41564 66444
rect 36912 65952 36964 65958
rect 36912 65894 36964 65900
rect 36924 52970 36952 65894
rect 39220 65852 39516 65872
rect 39276 65850 39300 65852
rect 39356 65850 39380 65852
rect 39436 65850 39460 65852
rect 39298 65798 39300 65850
rect 39362 65798 39374 65850
rect 39436 65798 39438 65850
rect 39276 65796 39300 65798
rect 39356 65796 39380 65798
rect 39436 65796 39460 65798
rect 39220 65776 39516 65796
rect 37924 65748 37976 65754
rect 37924 65690 37976 65696
rect 37464 55140 37516 55146
rect 37464 55082 37516 55088
rect 37476 53786 37504 55082
rect 37464 53780 37516 53786
rect 37464 53722 37516 53728
rect 37188 53440 37240 53446
rect 37188 53382 37240 53388
rect 36912 52964 36964 52970
rect 36912 52906 36964 52912
rect 37200 42634 37228 53382
rect 37188 42628 37240 42634
rect 37188 42570 37240 42576
rect 37200 41478 37228 42570
rect 37832 41812 37884 41818
rect 37832 41754 37884 41760
rect 36728 41472 36780 41478
rect 36728 41414 36780 41420
rect 37188 41472 37240 41478
rect 37188 41414 37240 41420
rect 36636 31952 36688 31958
rect 36636 31894 36688 31900
rect 36544 24268 36596 24274
rect 36544 24210 36596 24216
rect 36648 23594 36676 31894
rect 36740 25906 36768 41414
rect 37004 31884 37056 31890
rect 37004 31826 37056 31832
rect 36728 25900 36780 25906
rect 36728 25842 36780 25848
rect 36912 24744 36964 24750
rect 36912 24686 36964 24692
rect 36636 23588 36688 23594
rect 36636 23530 36688 23536
rect 36648 19854 36676 23530
rect 36924 21622 36952 24686
rect 36912 21616 36964 21622
rect 36912 21558 36964 21564
rect 36636 19848 36688 19854
rect 36636 19790 36688 19796
rect 37016 17542 37044 31826
rect 37648 31748 37700 31754
rect 37648 31690 37700 31696
rect 37660 31482 37688 31690
rect 37648 31476 37700 31482
rect 37648 31418 37700 31424
rect 37096 30864 37148 30870
rect 37096 30806 37148 30812
rect 37108 30326 37136 30806
rect 37648 30796 37700 30802
rect 37648 30738 37700 30744
rect 37660 30598 37688 30738
rect 37556 30592 37608 30598
rect 37556 30534 37608 30540
rect 37648 30592 37700 30598
rect 37648 30534 37700 30540
rect 37096 30320 37148 30326
rect 37096 30262 37148 30268
rect 37568 23254 37596 30534
rect 37556 23248 37608 23254
rect 37556 23190 37608 23196
rect 37660 22438 37688 30534
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 37648 22432 37700 22438
rect 37648 22374 37700 22380
rect 37752 22094 37780 23666
rect 37844 22438 37872 41754
rect 37936 26450 37964 65690
rect 39220 64764 39516 64784
rect 39276 64762 39300 64764
rect 39356 64762 39380 64764
rect 39436 64762 39460 64764
rect 39298 64710 39300 64762
rect 39362 64710 39374 64762
rect 39436 64710 39438 64762
rect 39276 64708 39300 64710
rect 39356 64708 39380 64710
rect 39436 64708 39460 64710
rect 39220 64688 39516 64708
rect 38108 64116 38160 64122
rect 38108 64058 38160 64064
rect 38016 55616 38068 55622
rect 38016 55558 38068 55564
rect 38028 55214 38056 55558
rect 38016 55208 38068 55214
rect 38016 55150 38068 55156
rect 37924 26444 37976 26450
rect 37924 26386 37976 26392
rect 37924 22976 37976 22982
rect 37924 22918 37976 22924
rect 37936 22506 37964 22918
rect 37924 22500 37976 22506
rect 37924 22442 37976 22448
rect 37832 22432 37884 22438
rect 37832 22374 37884 22380
rect 37844 22234 37872 22374
rect 37832 22228 37884 22234
rect 37832 22170 37884 22176
rect 37752 22066 37964 22094
rect 37004 17536 37056 17542
rect 37004 17478 37056 17484
rect 35716 14340 35768 14346
rect 35716 14282 35768 14288
rect 37936 13870 37964 22066
rect 37648 13864 37700 13870
rect 37648 13806 37700 13812
rect 37924 13864 37976 13870
rect 37924 13806 37976 13812
rect 37464 13320 37516 13326
rect 37464 13262 37516 13268
rect 37188 12708 37240 12714
rect 37188 12650 37240 12656
rect 32784 12406 32904 12434
rect 23940 12378 23992 12384
rect 32680 10124 32732 10130
rect 32680 10066 32732 10072
rect 32588 9920 32640 9926
rect 32588 9862 32640 9868
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18786 6352 18842 6361
rect 18786 6287 18842 6296
rect 18800 4690 18828 6287
rect 18878 5808 18934 5817
rect 18878 5743 18934 5752
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18892 4570 18920 5743
rect 18800 4542 18920 4570
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18616 3862 18736 3890
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18236 1420 18288 1426
rect 18340 1414 18460 1442
rect 18236 1362 18288 1368
rect 18248 800 18276 1362
rect 18432 800 18460 1414
rect 18524 800 18552 2994
rect 18616 2514 18644 2994
rect 18708 2854 18736 3862
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18800 2666 18828 4542
rect 18984 4434 19012 6598
rect 18892 4406 19012 4434
rect 18892 2961 18920 4406
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18878 2952 18934 2961
rect 18878 2887 18934 2896
rect 18878 2816 18934 2825
rect 18878 2751 18934 2760
rect 18892 2689 18920 2751
rect 18708 2638 18828 2666
rect 18878 2680 18934 2689
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18708 800 18736 2638
rect 18878 2615 18934 2624
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18800 800 18828 2518
rect 18984 800 19012 3878
rect 19076 3466 19104 6802
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 19168 3398 19196 6258
rect 19352 6254 19380 8842
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 3874 19380 5646
rect 19340 3868 19392 3874
rect 19340 3810 19392 3816
rect 19444 3806 19472 7142
rect 19432 3800 19484 3806
rect 19432 3742 19484 3748
rect 19156 3392 19208 3398
rect 19062 3360 19118 3369
rect 19156 3334 19208 3340
rect 19062 3295 19118 3304
rect 19076 3262 19104 3295
rect 19064 3256 19116 3262
rect 19064 3198 19116 3204
rect 19154 2952 19210 2961
rect 19154 2887 19210 2896
rect 19064 1896 19116 1902
rect 19064 1838 19116 1844
rect 19076 800 19104 1838
rect 19168 1426 19196 2887
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19248 1760 19300 1766
rect 19248 1702 19300 1708
rect 19156 1420 19208 1426
rect 19156 1362 19208 1368
rect 19260 800 19288 1702
rect 19444 800 19472 2246
rect 19536 800 19564 7346
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19628 3942 19656 5578
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 19720 800 19748 3606
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19812 800 19840 2790
rect 19904 1426 19932 6190
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 19892 1420 19944 1426
rect 19892 1362 19944 1368
rect 19996 800 20024 4150
rect 20088 800 20116 5714
rect 20364 2922 20392 5850
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20272 800 20300 2858
rect 20456 2774 20484 6394
rect 20720 5296 20772 5302
rect 20720 5238 20772 5244
rect 20732 3992 20760 5238
rect 20732 3964 20852 3992
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20364 2746 20484 2774
rect 20364 800 20392 2746
rect 20536 1420 20588 1426
rect 20536 1362 20588 1368
rect 20548 800 20576 1362
rect 20640 800 20668 3538
rect 20824 800 20852 3964
rect 20916 3534 20944 6666
rect 21008 3738 21036 7822
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20916 800 20944 3334
rect 21100 3126 21128 8298
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21178 5672 21234 5681
rect 21178 5607 21234 5616
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 21192 2854 21220 5607
rect 21456 4548 21508 4554
rect 21456 4490 21508 4496
rect 21272 3936 21324 3942
rect 21272 3878 21324 3884
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21088 2032 21140 2038
rect 21088 1974 21140 1980
rect 21100 800 21128 1974
rect 21284 800 21312 3878
rect 21364 3868 21416 3874
rect 21364 3810 21416 3816
rect 21376 800 21404 3810
rect 21468 3398 21496 4490
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21560 800 21588 3946
rect 21744 3942 21772 7210
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21732 3936 21784 3942
rect 21638 3904 21694 3913
rect 21732 3878 21784 3884
rect 21638 3839 21694 3848
rect 21652 3670 21680 3839
rect 21640 3664 21692 3670
rect 21640 3606 21692 3612
rect 21640 3256 21692 3262
rect 21640 3198 21692 3204
rect 21652 800 21680 3198
rect 21836 800 21864 5170
rect 22572 3874 22600 6326
rect 22664 4010 22692 6734
rect 23308 4282 23336 7958
rect 23388 6180 23440 6186
rect 23388 6122 23440 6128
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 22652 4004 22704 4010
rect 22652 3946 22704 3952
rect 22560 3868 22612 3874
rect 22560 3810 22612 3816
rect 22650 3768 22706 3777
rect 22650 3703 22706 3712
rect 22664 3602 22692 3703
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22652 3460 22704 3466
rect 22652 3402 22704 3408
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 21916 1964 21968 1970
rect 21916 1906 21968 1912
rect 22100 1964 22152 1970
rect 22100 1906 22152 1912
rect 21928 800 21956 1906
rect 22112 800 22140 1906
rect 22192 1760 22244 1766
rect 22192 1702 22244 1708
rect 22204 800 22232 1702
rect 22572 1578 22600 2926
rect 22664 1766 22692 3402
rect 22744 2712 22796 2718
rect 22744 2654 22796 2660
rect 23112 2712 23164 2718
rect 23112 2654 23164 2660
rect 22652 1760 22704 1766
rect 22652 1702 22704 1708
rect 22756 1578 22784 2654
rect 22928 2168 22980 2174
rect 22928 2110 22980 2116
rect 22836 2032 22888 2038
rect 22836 1974 22888 1980
rect 22388 1550 22600 1578
rect 22664 1550 22784 1578
rect 22388 800 22416 1550
rect 22468 1488 22520 1494
rect 22468 1430 22520 1436
rect 22480 800 22508 1430
rect 22664 800 22692 1550
rect 22848 800 22876 1974
rect 22940 800 22968 2110
rect 23124 800 23152 2654
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 23216 800 23244 2042
rect 23308 2038 23336 4082
rect 23400 4026 23428 6122
rect 23478 5944 23534 5953
rect 23478 5879 23534 5888
rect 23492 5114 23520 5879
rect 23584 5302 23612 8774
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23492 5086 23612 5114
rect 23400 3998 23520 4026
rect 23492 3806 23520 3998
rect 23388 3800 23440 3806
rect 23388 3742 23440 3748
rect 23480 3800 23532 3806
rect 23480 3742 23532 3748
rect 23400 2854 23428 3742
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23388 2712 23440 2718
rect 23388 2654 23440 2660
rect 23296 2032 23348 2038
rect 23296 1974 23348 1980
rect 23400 800 23428 2654
rect 23492 800 23520 3470
rect 23584 2922 23612 5086
rect 23676 3466 23704 7754
rect 23768 4690 23796 7890
rect 23860 4962 23888 9386
rect 23952 6225 23980 9522
rect 32600 9180 32628 9862
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 23938 6216 23994 6225
rect 23938 6151 23994 6160
rect 23938 6080 23994 6089
rect 23938 6015 23994 6024
rect 23848 4956 23900 4962
rect 23848 4898 23900 4904
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23756 3800 23808 3806
rect 23756 3742 23808 3748
rect 23664 3460 23716 3466
rect 23664 3402 23716 3408
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23676 800 23704 3130
rect 23768 800 23796 3742
rect 23860 2122 23888 3946
rect 23952 3806 23980 6015
rect 24504 5574 24532 8434
rect 24964 5574 24992 8978
rect 32312 8900 32364 8906
rect 32312 8842 32364 8848
rect 31944 8492 31996 8498
rect 31944 8434 31996 8440
rect 31760 6996 31812 7002
rect 31760 6938 31812 6944
rect 31772 5574 31800 6938
rect 31956 5642 31984 8434
rect 32036 7948 32088 7954
rect 32036 7890 32088 7896
rect 31944 5636 31996 5642
rect 31944 5578 31996 5584
rect 32048 5574 32076 7890
rect 32324 5574 32352 8842
rect 32496 7200 32548 7206
rect 32496 7142 32548 7148
rect 32508 5574 32536 7142
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 31760 5568 31812 5574
rect 31760 5510 31812 5516
rect 32036 5568 32088 5574
rect 32036 5510 32088 5516
rect 32312 5568 32364 5574
rect 32312 5510 32364 5516
rect 32496 5568 32548 5574
rect 32496 5510 32548 5516
rect 23940 3800 23992 3806
rect 23940 3742 23992 3748
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 23952 2258 23980 3334
rect 24044 2650 24072 5236
rect 24492 4888 24544 4894
rect 24122 4856 24178 4865
rect 24492 4830 24544 4836
rect 31760 4888 31812 4894
rect 31760 4830 31812 4836
rect 32036 4888 32088 4894
rect 32036 4830 32088 4836
rect 24122 4791 24178 4800
rect 24136 2854 24164 4791
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24308 3868 24360 3874
rect 24308 3810 24360 3816
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 23952 2230 24072 2258
rect 23860 2094 23980 2122
rect 23952 800 23980 2094
rect 24044 800 24072 2230
rect 24228 800 24256 3538
rect 24320 800 24348 3810
rect 24412 3126 24440 4626
rect 24504 3194 24532 4830
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24964 4026 24992 4082
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 24492 1692 24544 1698
rect 24492 1634 24544 1640
rect 24504 800 24532 1634
rect 24688 800 24716 4014
rect 24964 3998 25084 4026
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24780 800 24808 3878
rect 24952 3052 25004 3058
rect 24952 2994 25004 3000
rect 24964 1494 24992 2994
rect 24952 1488 25004 1494
rect 24952 1430 25004 1436
rect 24952 1352 25004 1358
rect 24952 1294 25004 1300
rect 24964 800 24992 1294
rect 25056 800 25084 3998
rect 31668 3664 31720 3670
rect 31668 3606 31720 3612
rect 31680 2922 31708 3606
rect 31668 2916 31720 2922
rect 31668 2858 31720 2864
rect 31668 2508 31720 2514
rect 31668 2450 31720 2456
rect 26332 1964 26384 1970
rect 26332 1906 26384 1912
rect 26516 1964 26568 1970
rect 26516 1906 26568 1912
rect 26608 1964 26660 1970
rect 26608 1906 26660 1912
rect 26884 1964 26936 1970
rect 26884 1906 26936 1912
rect 27160 1964 27212 1970
rect 27160 1906 27212 1912
rect 27436 1964 27488 1970
rect 27436 1906 27488 1912
rect 27620 1964 27672 1970
rect 27620 1906 27672 1912
rect 27896 1964 27948 1970
rect 27896 1906 27948 1912
rect 28724 1964 28776 1970
rect 28724 1906 28776 1912
rect 29000 1964 29052 1970
rect 29000 1906 29052 1912
rect 29184 1964 29236 1970
rect 29184 1906 29236 1912
rect 29276 1964 29328 1970
rect 29276 1906 29328 1912
rect 25320 1896 25372 1902
rect 25320 1838 25372 1844
rect 25596 1896 25648 1902
rect 25596 1838 25648 1844
rect 25780 1896 25832 1902
rect 25780 1838 25832 1844
rect 25872 1896 25924 1902
rect 25872 1838 25924 1844
rect 26056 1896 26108 1902
rect 26056 1838 26108 1844
rect 26148 1896 26200 1902
rect 26148 1838 26200 1844
rect 25228 1488 25280 1494
rect 25228 1430 25280 1436
rect 25240 800 25268 1430
rect 25332 800 25360 1838
rect 25504 1828 25556 1834
rect 25504 1770 25556 1776
rect 25516 800 25544 1770
rect 25608 800 25636 1838
rect 25688 1760 25740 1766
rect 25688 1702 25740 1708
rect 25700 1426 25728 1702
rect 25688 1420 25740 1426
rect 25688 1362 25740 1368
rect 25792 800 25820 1838
rect 25884 800 25912 1838
rect 26068 800 26096 1838
rect 26160 800 26188 1838
rect 26344 800 26372 1906
rect 26528 800 26556 1906
rect 26620 800 26648 1906
rect 26792 1896 26844 1902
rect 26792 1838 26844 1844
rect 26804 800 26832 1838
rect 26896 800 26924 1906
rect 27068 1488 27120 1494
rect 27068 1430 27120 1436
rect 27080 800 27108 1430
rect 27172 800 27200 1906
rect 27344 1896 27396 1902
rect 27344 1838 27396 1844
rect 27356 800 27384 1838
rect 27448 800 27476 1906
rect 27632 800 27660 1906
rect 27710 1864 27766 1873
rect 27710 1799 27766 1808
rect 27724 800 27752 1799
rect 27908 800 27936 1906
rect 28448 1896 28500 1902
rect 28078 1864 28134 1873
rect 28448 1838 28500 1844
rect 28078 1799 28134 1808
rect 28092 800 28120 1799
rect 28170 1728 28226 1737
rect 28170 1663 28226 1672
rect 28184 800 28212 1663
rect 28356 1624 28408 1630
rect 28356 1566 28408 1572
rect 28368 800 28396 1566
rect 28460 800 28488 1838
rect 28632 1760 28684 1766
rect 28632 1702 28684 1708
rect 28644 800 28672 1702
rect 28736 800 28764 1906
rect 28906 1728 28962 1737
rect 28906 1663 28962 1672
rect 28920 800 28948 1663
rect 29012 800 29040 1906
rect 29196 800 29224 1906
rect 29288 800 29316 1906
rect 29918 1864 29974 1873
rect 29918 1799 29974 1808
rect 30194 1864 30250 1873
rect 30194 1799 30250 1808
rect 31022 1864 31078 1873
rect 31022 1799 31078 1808
rect 29552 1760 29604 1766
rect 29552 1702 29604 1708
rect 29460 1556 29512 1562
rect 29460 1498 29512 1504
rect 29472 800 29500 1498
rect 29564 800 29592 1702
rect 29736 1420 29788 1426
rect 29736 1362 29788 1368
rect 29748 800 29776 1362
rect 29932 800 29960 1799
rect 30012 1760 30064 1766
rect 30012 1702 30064 1708
rect 30024 800 30052 1702
rect 30208 800 30236 1799
rect 30288 1556 30340 1562
rect 30288 1498 30340 1504
rect 30564 1556 30616 1562
rect 30564 1498 30616 1504
rect 30840 1556 30892 1562
rect 30840 1498 30892 1504
rect 30300 800 30328 1498
rect 30472 1352 30524 1358
rect 30472 1294 30524 1300
rect 30484 800 30512 1294
rect 30576 800 30604 1498
rect 30748 1352 30800 1358
rect 30748 1294 30800 1300
rect 30760 800 30788 1294
rect 30852 800 30880 1498
rect 31036 800 31064 1799
rect 31116 1692 31168 1698
rect 31116 1634 31168 1640
rect 31300 1692 31352 1698
rect 31300 1634 31352 1640
rect 31576 1692 31628 1698
rect 31576 1634 31628 1640
rect 31128 800 31156 1634
rect 31312 800 31340 1634
rect 31392 1556 31444 1562
rect 31392 1498 31444 1504
rect 31404 800 31432 1498
rect 31588 800 31616 1634
rect 31680 1426 31708 2450
rect 31772 1970 31800 4830
rect 31944 4684 31996 4690
rect 31944 4626 31996 4632
rect 31850 3496 31906 3505
rect 31850 3431 31906 3440
rect 31864 2990 31892 3431
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 31852 2712 31904 2718
rect 31852 2654 31904 2660
rect 31760 1964 31812 1970
rect 31760 1906 31812 1912
rect 31864 1442 31892 2654
rect 31956 1902 31984 4626
rect 32048 2786 32076 4830
rect 32036 2780 32088 2786
rect 32036 2722 32088 2728
rect 32036 2576 32088 2582
rect 32036 2518 32088 2524
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 31944 1896 31996 1902
rect 31944 1838 31996 1844
rect 31668 1420 31720 1426
rect 31668 1362 31720 1368
rect 31772 1414 31892 1442
rect 31772 800 31800 1414
rect 31850 1184 31906 1193
rect 31850 1119 31906 1128
rect 31864 800 31892 1119
rect 32048 800 32076 2518
rect 32140 800 32168 2518
rect 32232 2106 32260 5236
rect 32312 4888 32364 4894
rect 32312 4830 32364 4836
rect 32496 4888 32548 4894
rect 32496 4830 32548 4836
rect 32220 2100 32272 2106
rect 32220 2042 32272 2048
rect 32324 800 32352 4830
rect 32402 3904 32458 3913
rect 32402 3839 32458 3848
rect 32416 3806 32444 3839
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32508 2774 32536 4830
rect 32588 4140 32640 4146
rect 32588 4082 32640 4088
rect 32600 2922 32628 4082
rect 32588 2916 32640 2922
rect 32588 2858 32640 2864
rect 32508 2746 32628 2774
rect 32600 1442 32628 2746
rect 32416 1414 32628 1442
rect 32416 800 32444 1414
rect 32588 1352 32640 1358
rect 32588 1294 32640 1300
rect 32600 800 32628 1294
rect 32692 800 32720 10066
rect 32772 9036 32824 9042
rect 32772 8978 32824 8984
rect 32784 3641 32812 8978
rect 32770 3632 32826 3641
rect 32770 3567 32826 3576
rect 32772 3528 32824 3534
rect 32772 3470 32824 3476
rect 32784 2854 32812 3470
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 32772 2644 32824 2650
rect 32772 2586 32824 2592
rect 32784 1426 32812 2586
rect 32876 2446 32904 12406
rect 37200 10062 37228 12650
rect 37372 10600 37424 10606
rect 37372 10542 37424 10548
rect 36084 10056 36136 10062
rect 36084 9998 36136 10004
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 34888 8968 34940 8974
rect 34888 8910 34940 8916
rect 32956 8356 33008 8362
rect 32956 8298 33008 8304
rect 32968 2990 32996 8298
rect 33048 7268 33100 7274
rect 33048 7210 33100 7216
rect 33060 5234 33088 7210
rect 33138 5808 33194 5817
rect 33138 5743 33194 5752
rect 33968 5772 34020 5778
rect 33048 5228 33100 5234
rect 33048 5170 33100 5176
rect 33046 5128 33102 5137
rect 33046 5063 33102 5072
rect 33060 4962 33088 5063
rect 33048 4956 33100 4962
rect 33048 4898 33100 4904
rect 33048 4412 33100 4418
rect 33048 4354 33100 4360
rect 33060 4060 33088 4354
rect 33152 4214 33180 5743
rect 33968 5714 34020 5720
rect 33140 4208 33192 4214
rect 33140 4150 33192 4156
rect 33980 4078 34008 5714
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 33968 4072 34020 4078
rect 33060 4032 33180 4060
rect 33048 3732 33100 3738
rect 33048 3674 33100 3680
rect 33060 3641 33088 3674
rect 33046 3632 33102 3641
rect 33046 3567 33102 3576
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32968 1578 32996 2790
rect 32876 1550 32996 1578
rect 32772 1420 32824 1426
rect 32772 1362 32824 1368
rect 32876 800 32904 1550
rect 32956 1352 33008 1358
rect 32956 1294 33008 1300
rect 32968 800 32996 1294
rect 33152 800 33180 4032
rect 33968 4014 34020 4020
rect 33966 3768 34022 3777
rect 33966 3703 33968 3712
rect 34020 3703 34022 3712
rect 33968 3674 34020 3680
rect 33874 3360 33930 3369
rect 33874 3295 33930 3304
rect 33888 3262 33916 3295
rect 33876 3256 33928 3262
rect 33876 3198 33928 3204
rect 33324 2712 33376 2718
rect 33324 2654 33376 2660
rect 33336 800 33364 2654
rect 33416 2576 33468 2582
rect 33416 2518 33468 2524
rect 33692 2576 33744 2582
rect 33692 2518 33744 2524
rect 33428 800 33456 2518
rect 33600 2372 33652 2378
rect 33600 2314 33652 2320
rect 33612 800 33640 2314
rect 33704 800 33732 2518
rect 34152 1964 34204 1970
rect 34152 1906 34204 1912
rect 34428 1964 34480 1970
rect 34428 1906 34480 1912
rect 33876 1284 33928 1290
rect 33876 1226 33928 1232
rect 33888 800 33916 1226
rect 33968 1012 34020 1018
rect 33968 954 34020 960
rect 33980 800 34008 954
rect 34164 800 34192 1906
rect 34244 1692 34296 1698
rect 34244 1634 34296 1640
rect 34256 800 34284 1634
rect 34440 800 34468 1906
rect 34624 1442 34652 4558
rect 34702 3224 34758 3233
rect 34702 3159 34704 3168
rect 34756 3159 34758 3168
rect 34704 3130 34756 3136
rect 34702 2816 34758 2825
rect 34900 2774 34928 8910
rect 34980 8016 35032 8022
rect 34980 7958 35032 7964
rect 34702 2751 34758 2760
rect 34532 1414 34652 1442
rect 34532 800 34560 1414
rect 34716 800 34744 2751
rect 34808 2746 34928 2774
rect 34808 800 34836 2746
rect 34992 800 35020 7958
rect 35256 7540 35308 7546
rect 35256 7482 35308 7488
rect 35162 6896 35218 6905
rect 35162 6831 35218 6840
rect 35072 4548 35124 4554
rect 35072 4490 35124 4496
rect 35084 3602 35112 4490
rect 35176 4418 35204 6831
rect 35164 4412 35216 4418
rect 35164 4354 35216 4360
rect 35072 3596 35124 3602
rect 35072 3538 35124 3544
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 35072 3120 35124 3126
rect 35072 3062 35124 3068
rect 35084 2825 35112 3062
rect 35070 2816 35126 2825
rect 35070 2751 35126 2760
rect 35176 800 35204 3538
rect 35268 800 35296 7482
rect 35624 7472 35676 7478
rect 35624 7414 35676 7420
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 35348 6180 35400 6186
rect 35348 6122 35400 6128
rect 35360 3262 35388 6122
rect 35440 6112 35492 6118
rect 35440 6054 35492 6060
rect 35452 3806 35480 6054
rect 35440 3800 35492 3806
rect 35440 3742 35492 3748
rect 35544 3738 35572 6258
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 35636 3652 35664 7414
rect 35992 5908 36044 5914
rect 35992 5850 36044 5856
rect 36004 4060 36032 5850
rect 35820 4032 36032 4060
rect 35636 3624 35756 3652
rect 35532 3324 35584 3330
rect 35532 3266 35584 3272
rect 35348 3256 35400 3262
rect 35348 3198 35400 3204
rect 35440 3256 35492 3262
rect 35440 3198 35492 3204
rect 35452 800 35480 3198
rect 35544 800 35572 3266
rect 35728 800 35756 3624
rect 35820 800 35848 4032
rect 35990 3768 36046 3777
rect 35990 3703 36046 3712
rect 36004 3097 36032 3703
rect 35990 3088 36046 3097
rect 35990 3023 36046 3032
rect 36096 1154 36124 9998
rect 37280 9512 37332 9518
rect 37280 9454 37332 9460
rect 37096 8424 37148 8430
rect 37096 8366 37148 8372
rect 36912 8084 36964 8090
rect 36912 8026 36964 8032
rect 36268 7404 36320 7410
rect 36268 7346 36320 7352
rect 36176 5364 36228 5370
rect 36176 5306 36228 5312
rect 36084 1148 36136 1154
rect 36084 1090 36136 1096
rect 36188 1034 36216 5306
rect 36004 1006 36216 1034
rect 36004 800 36032 1006
rect 36084 944 36136 950
rect 36084 886 36136 892
rect 36096 800 36124 886
rect 36280 800 36308 7346
rect 36726 6488 36782 6497
rect 36726 6423 36782 6432
rect 36544 6384 36596 6390
rect 36544 6326 36596 6332
rect 36360 3664 36412 3670
rect 36360 3606 36412 3612
rect 36372 800 36400 3606
rect 36556 800 36584 6326
rect 36740 2718 36768 6423
rect 36820 5636 36872 5642
rect 36820 5578 36872 5584
rect 36728 2712 36780 2718
rect 36728 2654 36780 2660
rect 36634 2408 36690 2417
rect 36634 2343 36690 2352
rect 36648 800 36676 2343
rect 36832 800 36860 5578
rect 36924 2774 36952 8026
rect 37004 6724 37056 6730
rect 37004 6666 37056 6672
rect 37016 3074 37044 6666
rect 37108 3262 37136 8366
rect 37292 5506 37320 9454
rect 37280 5500 37332 5506
rect 37280 5442 37332 5448
rect 37188 5024 37240 5030
rect 37188 4966 37240 4972
rect 37200 3602 37228 4966
rect 37280 3732 37332 3738
rect 37280 3674 37332 3680
rect 37188 3596 37240 3602
rect 37188 3538 37240 3544
rect 37096 3256 37148 3262
rect 37096 3198 37148 3204
rect 37016 3046 37136 3074
rect 36924 2746 37044 2774
rect 37016 800 37044 2746
rect 37108 800 37136 3046
rect 37292 800 37320 3674
rect 37384 800 37412 10542
rect 37476 2990 37504 13262
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37568 4690 37596 12786
rect 37556 4684 37608 4690
rect 37556 4626 37608 4632
rect 37660 3670 37688 13806
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 37752 10606 37780 13126
rect 37832 12640 37884 12646
rect 37832 12582 37884 12588
rect 37740 10600 37792 10606
rect 37740 10542 37792 10548
rect 37844 10130 37872 12582
rect 37922 12200 37978 12209
rect 37922 12135 37978 12144
rect 37936 11218 37964 12135
rect 38028 11898 38056 55150
rect 38120 16574 38148 64058
rect 39220 63676 39516 63696
rect 39276 63674 39300 63676
rect 39356 63674 39380 63676
rect 39436 63674 39460 63676
rect 39298 63622 39300 63674
rect 39362 63622 39374 63674
rect 39436 63622 39438 63674
rect 39276 63620 39300 63622
rect 39356 63620 39380 63622
rect 39436 63620 39460 63622
rect 39220 63600 39516 63620
rect 39220 62588 39516 62608
rect 39276 62586 39300 62588
rect 39356 62586 39380 62588
rect 39436 62586 39460 62588
rect 39298 62534 39300 62586
rect 39362 62534 39374 62586
rect 39436 62534 39438 62586
rect 39276 62532 39300 62534
rect 39356 62532 39380 62534
rect 39436 62532 39460 62534
rect 39220 62512 39516 62532
rect 39220 61500 39516 61520
rect 39276 61498 39300 61500
rect 39356 61498 39380 61500
rect 39436 61498 39460 61500
rect 39298 61446 39300 61498
rect 39362 61446 39374 61498
rect 39436 61446 39438 61498
rect 39276 61444 39300 61446
rect 39356 61444 39380 61446
rect 39436 61444 39460 61446
rect 39220 61424 39516 61444
rect 39220 60412 39516 60432
rect 39276 60410 39300 60412
rect 39356 60410 39380 60412
rect 39436 60410 39460 60412
rect 39298 60358 39300 60410
rect 39362 60358 39374 60410
rect 39436 60358 39438 60410
rect 39276 60356 39300 60358
rect 39356 60356 39380 60358
rect 39436 60356 39460 60358
rect 39220 60336 39516 60356
rect 39220 59324 39516 59344
rect 39276 59322 39300 59324
rect 39356 59322 39380 59324
rect 39436 59322 39460 59324
rect 39298 59270 39300 59322
rect 39362 59270 39374 59322
rect 39436 59270 39438 59322
rect 39276 59268 39300 59270
rect 39356 59268 39380 59270
rect 39436 59268 39460 59270
rect 39220 59248 39516 59268
rect 39220 58236 39516 58256
rect 39276 58234 39300 58236
rect 39356 58234 39380 58236
rect 39436 58234 39460 58236
rect 39298 58182 39300 58234
rect 39362 58182 39374 58234
rect 39436 58182 39438 58234
rect 39276 58180 39300 58182
rect 39356 58180 39380 58182
rect 39436 58180 39460 58182
rect 39220 58160 39516 58180
rect 39220 57148 39516 57168
rect 39276 57146 39300 57148
rect 39356 57146 39380 57148
rect 39436 57146 39460 57148
rect 39298 57094 39300 57146
rect 39362 57094 39374 57146
rect 39436 57094 39438 57146
rect 39276 57092 39300 57094
rect 39356 57092 39380 57094
rect 39436 57092 39460 57094
rect 39220 57072 39516 57092
rect 39220 56060 39516 56080
rect 39276 56058 39300 56060
rect 39356 56058 39380 56060
rect 39436 56058 39460 56060
rect 39298 56006 39300 56058
rect 39362 56006 39374 56058
rect 39436 56006 39438 56058
rect 39276 56004 39300 56006
rect 39356 56004 39380 56006
rect 39436 56004 39460 56006
rect 39220 55984 39516 56004
rect 39948 55344 40000 55350
rect 39948 55286 40000 55292
rect 38752 55208 38804 55214
rect 38752 55150 38804 55156
rect 38384 55072 38436 55078
rect 38384 55014 38436 55020
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38212 28422 38240 35974
rect 38200 28416 38252 28422
rect 38200 28358 38252 28364
rect 38396 26790 38424 55014
rect 38764 54534 38792 55150
rect 39220 54972 39516 54992
rect 39276 54970 39300 54972
rect 39356 54970 39380 54972
rect 39436 54970 39460 54972
rect 39298 54918 39300 54970
rect 39362 54918 39374 54970
rect 39436 54918 39438 54970
rect 39276 54916 39300 54918
rect 39356 54916 39380 54918
rect 39436 54916 39460 54918
rect 39220 54896 39516 54916
rect 38752 54528 38804 54534
rect 38752 54470 38804 54476
rect 39220 53884 39516 53904
rect 39276 53882 39300 53884
rect 39356 53882 39380 53884
rect 39436 53882 39460 53884
rect 39298 53830 39300 53882
rect 39362 53830 39374 53882
rect 39436 53830 39438 53882
rect 39276 53828 39300 53830
rect 39356 53828 39380 53830
rect 39436 53828 39460 53830
rect 39220 53808 39516 53828
rect 39220 52796 39516 52816
rect 39276 52794 39300 52796
rect 39356 52794 39380 52796
rect 39436 52794 39460 52796
rect 39298 52742 39300 52794
rect 39362 52742 39374 52794
rect 39436 52742 39438 52794
rect 39276 52740 39300 52742
rect 39356 52740 39380 52742
rect 39436 52740 39460 52742
rect 39220 52720 39516 52740
rect 39960 52698 39988 55286
rect 39948 52692 40000 52698
rect 39948 52634 40000 52640
rect 39220 51708 39516 51728
rect 39276 51706 39300 51708
rect 39356 51706 39380 51708
rect 39436 51706 39460 51708
rect 39298 51654 39300 51706
rect 39362 51654 39374 51706
rect 39436 51654 39438 51706
rect 39276 51652 39300 51654
rect 39356 51652 39380 51654
rect 39436 51652 39460 51654
rect 39220 51632 39516 51652
rect 39960 51474 39988 52634
rect 39948 51468 40000 51474
rect 39948 51410 40000 51416
rect 39220 50620 39516 50640
rect 39276 50618 39300 50620
rect 39356 50618 39380 50620
rect 39436 50618 39460 50620
rect 39298 50566 39300 50618
rect 39362 50566 39374 50618
rect 39436 50566 39438 50618
rect 39276 50564 39300 50566
rect 39356 50564 39380 50566
rect 39436 50564 39460 50566
rect 39220 50544 39516 50564
rect 40132 49700 40184 49706
rect 40132 49642 40184 49648
rect 39220 49532 39516 49552
rect 39276 49530 39300 49532
rect 39356 49530 39380 49532
rect 39436 49530 39460 49532
rect 39298 49478 39300 49530
rect 39362 49478 39374 49530
rect 39436 49478 39438 49530
rect 39276 49476 39300 49478
rect 39356 49476 39380 49478
rect 39436 49476 39460 49478
rect 39220 49456 39516 49476
rect 40144 49094 40172 49642
rect 40132 49088 40184 49094
rect 40132 49030 40184 49036
rect 39220 48444 39516 48464
rect 39276 48442 39300 48444
rect 39356 48442 39380 48444
rect 39436 48442 39460 48444
rect 39298 48390 39300 48442
rect 39362 48390 39374 48442
rect 39436 48390 39438 48442
rect 39276 48388 39300 48390
rect 39356 48388 39380 48390
rect 39436 48388 39460 48390
rect 39220 48368 39516 48388
rect 39220 47356 39516 47376
rect 39276 47354 39300 47356
rect 39356 47354 39380 47356
rect 39436 47354 39460 47356
rect 39298 47302 39300 47354
rect 39362 47302 39374 47354
rect 39436 47302 39438 47354
rect 39276 47300 39300 47302
rect 39356 47300 39380 47302
rect 39436 47300 39460 47302
rect 39220 47280 39516 47300
rect 39220 46268 39516 46288
rect 39276 46266 39300 46268
rect 39356 46266 39380 46268
rect 39436 46266 39460 46268
rect 39298 46214 39300 46266
rect 39362 46214 39374 46266
rect 39436 46214 39438 46266
rect 39276 46212 39300 46214
rect 39356 46212 39380 46214
rect 39436 46212 39460 46214
rect 39220 46192 39516 46212
rect 39120 45824 39172 45830
rect 39120 45766 39172 45772
rect 39132 45354 39160 45766
rect 39948 45552 40000 45558
rect 39948 45494 40000 45500
rect 39120 45348 39172 45354
rect 39120 45290 39172 45296
rect 39132 42090 39160 45290
rect 39856 45280 39908 45286
rect 39856 45222 39908 45228
rect 39220 45180 39516 45200
rect 39276 45178 39300 45180
rect 39356 45178 39380 45180
rect 39436 45178 39460 45180
rect 39298 45126 39300 45178
rect 39362 45126 39374 45178
rect 39436 45126 39438 45178
rect 39276 45124 39300 45126
rect 39356 45124 39380 45126
rect 39436 45124 39460 45126
rect 39220 45104 39516 45124
rect 39220 44092 39516 44112
rect 39276 44090 39300 44092
rect 39356 44090 39380 44092
rect 39436 44090 39460 44092
rect 39298 44038 39300 44090
rect 39362 44038 39374 44090
rect 39436 44038 39438 44090
rect 39276 44036 39300 44038
rect 39356 44036 39380 44038
rect 39436 44036 39460 44038
rect 39220 44016 39516 44036
rect 39220 43004 39516 43024
rect 39276 43002 39300 43004
rect 39356 43002 39380 43004
rect 39436 43002 39460 43004
rect 39298 42950 39300 43002
rect 39362 42950 39374 43002
rect 39436 42950 39438 43002
rect 39276 42948 39300 42950
rect 39356 42948 39380 42950
rect 39436 42948 39460 42950
rect 39220 42928 39516 42948
rect 39120 42084 39172 42090
rect 39120 42026 39172 42032
rect 39220 41916 39516 41936
rect 39276 41914 39300 41916
rect 39356 41914 39380 41916
rect 39436 41914 39460 41916
rect 39298 41862 39300 41914
rect 39362 41862 39374 41914
rect 39436 41862 39438 41914
rect 39276 41860 39300 41862
rect 39356 41860 39380 41862
rect 39436 41860 39460 41862
rect 39220 41840 39516 41860
rect 39120 40928 39172 40934
rect 39120 40870 39172 40876
rect 39132 40526 39160 40870
rect 39220 40828 39516 40848
rect 39276 40826 39300 40828
rect 39356 40826 39380 40828
rect 39436 40826 39460 40828
rect 39298 40774 39300 40826
rect 39362 40774 39374 40826
rect 39436 40774 39438 40826
rect 39276 40772 39300 40774
rect 39356 40772 39380 40774
rect 39436 40772 39460 40774
rect 39220 40752 39516 40772
rect 39868 40526 39896 45222
rect 39120 40520 39172 40526
rect 39120 40462 39172 40468
rect 39856 40520 39908 40526
rect 39856 40462 39908 40468
rect 39132 30802 39160 40462
rect 39220 39740 39516 39760
rect 39276 39738 39300 39740
rect 39356 39738 39380 39740
rect 39436 39738 39460 39740
rect 39298 39686 39300 39738
rect 39362 39686 39374 39738
rect 39436 39686 39438 39738
rect 39276 39684 39300 39686
rect 39356 39684 39380 39686
rect 39436 39684 39460 39686
rect 39220 39664 39516 39684
rect 39220 38652 39516 38672
rect 39276 38650 39300 38652
rect 39356 38650 39380 38652
rect 39436 38650 39460 38652
rect 39298 38598 39300 38650
rect 39362 38598 39374 38650
rect 39436 38598 39438 38650
rect 39276 38596 39300 38598
rect 39356 38596 39380 38598
rect 39436 38596 39460 38598
rect 39220 38576 39516 38596
rect 39220 37564 39516 37584
rect 39276 37562 39300 37564
rect 39356 37562 39380 37564
rect 39436 37562 39460 37564
rect 39298 37510 39300 37562
rect 39362 37510 39374 37562
rect 39436 37510 39438 37562
rect 39276 37508 39300 37510
rect 39356 37508 39380 37510
rect 39436 37508 39460 37510
rect 39220 37488 39516 37508
rect 39220 36476 39516 36496
rect 39276 36474 39300 36476
rect 39356 36474 39380 36476
rect 39436 36474 39460 36476
rect 39298 36422 39300 36474
rect 39362 36422 39374 36474
rect 39436 36422 39438 36474
rect 39276 36420 39300 36422
rect 39356 36420 39380 36422
rect 39436 36420 39460 36422
rect 39220 36400 39516 36420
rect 39220 35388 39516 35408
rect 39276 35386 39300 35388
rect 39356 35386 39380 35388
rect 39436 35386 39460 35388
rect 39298 35334 39300 35386
rect 39362 35334 39374 35386
rect 39436 35334 39438 35386
rect 39276 35332 39300 35334
rect 39356 35332 39380 35334
rect 39436 35332 39460 35334
rect 39220 35312 39516 35332
rect 39960 35086 39988 45494
rect 40144 45422 40172 49030
rect 40408 47660 40460 47666
rect 40408 47602 40460 47608
rect 40316 47592 40368 47598
rect 40316 47534 40368 47540
rect 40328 45422 40356 47534
rect 40132 45416 40184 45422
rect 40132 45358 40184 45364
rect 40316 45416 40368 45422
rect 40316 45358 40368 45364
rect 40328 44742 40356 45358
rect 40316 44736 40368 44742
rect 40316 44678 40368 44684
rect 39948 35080 40000 35086
rect 39948 35022 40000 35028
rect 39220 34300 39516 34320
rect 39276 34298 39300 34300
rect 39356 34298 39380 34300
rect 39436 34298 39460 34300
rect 39298 34246 39300 34298
rect 39362 34246 39374 34298
rect 39436 34246 39438 34298
rect 39276 34244 39300 34246
rect 39356 34244 39380 34246
rect 39436 34244 39460 34246
rect 39220 34224 39516 34244
rect 39220 33212 39516 33232
rect 39276 33210 39300 33212
rect 39356 33210 39380 33212
rect 39436 33210 39460 33212
rect 39298 33158 39300 33210
rect 39362 33158 39374 33210
rect 39436 33158 39438 33210
rect 39276 33156 39300 33158
rect 39356 33156 39380 33158
rect 39436 33156 39460 33158
rect 39220 33136 39516 33156
rect 39220 32124 39516 32144
rect 39276 32122 39300 32124
rect 39356 32122 39380 32124
rect 39436 32122 39460 32124
rect 39298 32070 39300 32122
rect 39362 32070 39374 32122
rect 39436 32070 39438 32122
rect 39276 32068 39300 32070
rect 39356 32068 39380 32070
rect 39436 32068 39460 32070
rect 39220 32048 39516 32068
rect 39580 32020 39632 32026
rect 39580 31962 39632 31968
rect 39220 31036 39516 31056
rect 39276 31034 39300 31036
rect 39356 31034 39380 31036
rect 39436 31034 39460 31036
rect 39298 30982 39300 31034
rect 39362 30982 39374 31034
rect 39436 30982 39438 31034
rect 39276 30980 39300 30982
rect 39356 30980 39380 30982
rect 39436 30980 39460 30982
rect 39220 30960 39516 30980
rect 38660 30796 38712 30802
rect 38660 30738 38712 30744
rect 39120 30796 39172 30802
rect 39120 30738 39172 30744
rect 38384 26784 38436 26790
rect 38384 26726 38436 26732
rect 38672 22982 38700 30738
rect 38936 30184 38988 30190
rect 38936 30126 38988 30132
rect 38200 22976 38252 22982
rect 38200 22918 38252 22924
rect 38660 22976 38712 22982
rect 38660 22918 38712 22924
rect 38212 22574 38240 22918
rect 38568 22772 38620 22778
rect 38568 22714 38620 22720
rect 38200 22568 38252 22574
rect 38200 22510 38252 22516
rect 38580 22438 38608 22714
rect 38568 22432 38620 22438
rect 38568 22374 38620 22380
rect 38752 21616 38804 21622
rect 38752 21558 38804 21564
rect 38120 16546 38240 16574
rect 38108 14544 38160 14550
rect 38108 14486 38160 14492
rect 38120 14006 38148 14486
rect 38212 14278 38240 16546
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 38384 14272 38436 14278
rect 38384 14214 38436 14220
rect 38108 14000 38160 14006
rect 38108 13942 38160 13948
rect 38292 12980 38344 12986
rect 38292 12922 38344 12928
rect 38108 12096 38160 12102
rect 38108 12038 38160 12044
rect 38200 12096 38252 12102
rect 38304 12073 38332 12922
rect 38200 12038 38252 12044
rect 38290 12064 38346 12073
rect 38016 11892 38068 11898
rect 38016 11834 38068 11840
rect 38120 11830 38148 12038
rect 38108 11824 38160 11830
rect 38108 11766 38160 11772
rect 37924 11212 37976 11218
rect 37924 11154 37976 11160
rect 38108 11076 38160 11082
rect 38108 11018 38160 11024
rect 38016 10600 38068 10606
rect 38016 10542 38068 10548
rect 37924 10464 37976 10470
rect 37924 10406 37976 10412
rect 37832 10124 37884 10130
rect 37832 10066 37884 10072
rect 37740 9648 37792 9654
rect 37740 9590 37792 9596
rect 37752 8906 37780 9590
rect 37740 8900 37792 8906
rect 37740 8842 37792 8848
rect 37752 5574 37780 8842
rect 37936 7954 37964 10406
rect 38028 9654 38056 10542
rect 38016 9648 38068 9654
rect 38016 9590 38068 9596
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 37924 7948 37976 7954
rect 37924 7890 37976 7896
rect 37832 6656 37884 6662
rect 37832 6598 37884 6604
rect 37740 5568 37792 5574
rect 37740 5510 37792 5516
rect 37740 5160 37792 5166
rect 37740 5102 37792 5108
rect 37556 3664 37608 3670
rect 37556 3606 37608 3612
rect 37648 3664 37700 3670
rect 37648 3606 37700 3612
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37568 800 37596 3606
rect 37752 2774 37780 5102
rect 37660 2746 37780 2774
rect 37660 800 37688 2746
rect 37844 800 37872 6598
rect 37922 6352 37978 6361
rect 37922 6287 37924 6296
rect 37976 6287 37978 6296
rect 37924 6258 37976 6264
rect 37924 5704 37976 5710
rect 37924 5646 37976 5652
rect 37936 800 37964 5646
rect 38028 4026 38056 9318
rect 38120 7342 38148 11018
rect 38212 9042 38240 12038
rect 38290 11999 38346 12008
rect 38304 11694 38332 11999
rect 38292 11688 38344 11694
rect 38292 11630 38344 11636
rect 38292 9988 38344 9994
rect 38292 9930 38344 9936
rect 38200 9036 38252 9042
rect 38200 8978 38252 8984
rect 38108 7336 38160 7342
rect 38108 7278 38160 7284
rect 38120 4146 38148 7278
rect 38304 5250 38332 9930
rect 38396 5846 38424 14214
rect 38568 14000 38620 14006
rect 38568 13942 38620 13948
rect 38476 11552 38528 11558
rect 38476 11494 38528 11500
rect 38488 8430 38516 11494
rect 38580 10606 38608 13942
rect 38764 12986 38792 21558
rect 38844 20800 38896 20806
rect 38844 20742 38896 20748
rect 38752 12980 38804 12986
rect 38752 12922 38804 12928
rect 38660 11688 38712 11694
rect 38660 11630 38712 11636
rect 38568 10600 38620 10606
rect 38568 10542 38620 10548
rect 38568 10464 38620 10470
rect 38568 10406 38620 10412
rect 38476 8424 38528 8430
rect 38476 8366 38528 8372
rect 38476 6928 38528 6934
rect 38476 6870 38528 6876
rect 38384 5840 38436 5846
rect 38384 5782 38436 5788
rect 38304 5222 38424 5250
rect 38396 5098 38424 5222
rect 38384 5092 38436 5098
rect 38384 5034 38436 5040
rect 38488 4978 38516 6870
rect 38580 6866 38608 10406
rect 38672 8362 38700 11630
rect 38752 11076 38804 11082
rect 38752 11018 38804 11024
rect 38660 8356 38712 8362
rect 38660 8298 38712 8304
rect 38764 8106 38792 11018
rect 38672 8078 38792 8106
rect 38672 8022 38700 8078
rect 38660 8016 38712 8022
rect 38660 7958 38712 7964
rect 38660 7812 38712 7818
rect 38660 7754 38712 7760
rect 38568 6860 38620 6866
rect 38568 6802 38620 6808
rect 38580 5953 38608 6802
rect 38672 6089 38700 7754
rect 38750 7440 38806 7449
rect 38750 7375 38806 7384
rect 38764 7342 38792 7375
rect 38752 7336 38804 7342
rect 38752 7278 38804 7284
rect 38764 7206 38792 7278
rect 38752 7200 38804 7206
rect 38752 7142 38804 7148
rect 38752 6860 38804 6866
rect 38752 6802 38804 6808
rect 38658 6080 38714 6089
rect 38658 6015 38714 6024
rect 38566 5944 38622 5953
rect 38566 5879 38622 5888
rect 38568 5568 38620 5574
rect 38568 5510 38620 5516
rect 38396 4950 38516 4978
rect 38108 4140 38160 4146
rect 38108 4082 38160 4088
rect 38292 4140 38344 4146
rect 38292 4082 38344 4088
rect 38028 3998 38240 4026
rect 38108 1420 38160 1426
rect 38108 1362 38160 1368
rect 38120 800 38148 1362
rect 38212 800 38240 3998
rect 38304 3738 38332 4082
rect 38292 3732 38344 3738
rect 38292 3674 38344 3680
rect 38396 800 38424 4950
rect 38580 4876 38608 5510
rect 38488 4848 38608 4876
rect 38488 4010 38516 4848
rect 38568 4208 38620 4214
rect 38568 4150 38620 4156
rect 38658 4176 38714 4185
rect 38580 4010 38608 4150
rect 38658 4111 38714 4120
rect 38672 4078 38700 4111
rect 38660 4072 38712 4078
rect 38660 4014 38712 4020
rect 38476 4004 38528 4010
rect 38476 3946 38528 3952
rect 38568 4004 38620 4010
rect 38568 3946 38620 3952
rect 38764 3942 38792 6802
rect 38856 5166 38884 20742
rect 38948 18834 38976 30126
rect 39220 29948 39516 29968
rect 39276 29946 39300 29948
rect 39356 29946 39380 29948
rect 39436 29946 39460 29948
rect 39298 29894 39300 29946
rect 39362 29894 39374 29946
rect 39436 29894 39438 29946
rect 39276 29892 39300 29894
rect 39356 29892 39380 29894
rect 39436 29892 39460 29894
rect 39220 29872 39516 29892
rect 39220 28860 39516 28880
rect 39276 28858 39300 28860
rect 39356 28858 39380 28860
rect 39436 28858 39460 28860
rect 39298 28806 39300 28858
rect 39362 28806 39374 28858
rect 39436 28806 39438 28858
rect 39276 28804 39300 28806
rect 39356 28804 39380 28806
rect 39436 28804 39460 28806
rect 39220 28784 39516 28804
rect 39220 27772 39516 27792
rect 39276 27770 39300 27772
rect 39356 27770 39380 27772
rect 39436 27770 39460 27772
rect 39298 27718 39300 27770
rect 39362 27718 39374 27770
rect 39436 27718 39438 27770
rect 39276 27716 39300 27718
rect 39356 27716 39380 27718
rect 39436 27716 39460 27718
rect 39220 27696 39516 27716
rect 39220 26684 39516 26704
rect 39276 26682 39300 26684
rect 39356 26682 39380 26684
rect 39436 26682 39460 26684
rect 39298 26630 39300 26682
rect 39362 26630 39374 26682
rect 39436 26630 39438 26682
rect 39276 26628 39300 26630
rect 39356 26628 39380 26630
rect 39436 26628 39460 26630
rect 39220 26608 39516 26628
rect 39220 25596 39516 25616
rect 39276 25594 39300 25596
rect 39356 25594 39380 25596
rect 39436 25594 39460 25596
rect 39298 25542 39300 25594
rect 39362 25542 39374 25594
rect 39436 25542 39438 25594
rect 39276 25540 39300 25542
rect 39356 25540 39380 25542
rect 39436 25540 39460 25542
rect 39220 25520 39516 25540
rect 39220 24508 39516 24528
rect 39276 24506 39300 24508
rect 39356 24506 39380 24508
rect 39436 24506 39460 24508
rect 39298 24454 39300 24506
rect 39362 24454 39374 24506
rect 39436 24454 39438 24506
rect 39276 24452 39300 24454
rect 39356 24452 39380 24454
rect 39436 24452 39460 24454
rect 39220 24432 39516 24452
rect 39220 23420 39516 23440
rect 39276 23418 39300 23420
rect 39356 23418 39380 23420
rect 39436 23418 39460 23420
rect 39298 23366 39300 23418
rect 39362 23366 39374 23418
rect 39436 23366 39438 23418
rect 39276 23364 39300 23366
rect 39356 23364 39380 23366
rect 39436 23364 39460 23366
rect 39220 23344 39516 23364
rect 39220 22332 39516 22352
rect 39276 22330 39300 22332
rect 39356 22330 39380 22332
rect 39436 22330 39460 22332
rect 39298 22278 39300 22330
rect 39362 22278 39374 22330
rect 39436 22278 39438 22330
rect 39276 22276 39300 22278
rect 39356 22276 39380 22278
rect 39436 22276 39460 22278
rect 39220 22256 39516 22276
rect 39220 21244 39516 21264
rect 39276 21242 39300 21244
rect 39356 21242 39380 21244
rect 39436 21242 39460 21244
rect 39298 21190 39300 21242
rect 39362 21190 39374 21242
rect 39436 21190 39438 21242
rect 39276 21188 39300 21190
rect 39356 21188 39380 21190
rect 39436 21188 39460 21190
rect 39220 21168 39516 21188
rect 39220 20156 39516 20176
rect 39276 20154 39300 20156
rect 39356 20154 39380 20156
rect 39436 20154 39460 20156
rect 39298 20102 39300 20154
rect 39362 20102 39374 20154
rect 39436 20102 39438 20154
rect 39276 20100 39300 20102
rect 39356 20100 39380 20102
rect 39436 20100 39460 20102
rect 39220 20080 39516 20100
rect 39220 19068 39516 19088
rect 39276 19066 39300 19068
rect 39356 19066 39380 19068
rect 39436 19066 39460 19068
rect 39298 19014 39300 19066
rect 39362 19014 39374 19066
rect 39436 19014 39438 19066
rect 39276 19012 39300 19014
rect 39356 19012 39380 19014
rect 39436 19012 39460 19014
rect 39220 18992 39516 19012
rect 38936 18828 38988 18834
rect 38936 18770 38988 18776
rect 39220 17980 39516 18000
rect 39276 17978 39300 17980
rect 39356 17978 39380 17980
rect 39436 17978 39460 17980
rect 39298 17926 39300 17978
rect 39362 17926 39374 17978
rect 39436 17926 39438 17978
rect 39276 17924 39300 17926
rect 39356 17924 39380 17926
rect 39436 17924 39460 17926
rect 39220 17904 39516 17924
rect 39220 16892 39516 16912
rect 39276 16890 39300 16892
rect 39356 16890 39380 16892
rect 39436 16890 39460 16892
rect 39298 16838 39300 16890
rect 39362 16838 39374 16890
rect 39436 16838 39438 16890
rect 39276 16836 39300 16838
rect 39356 16836 39380 16838
rect 39436 16836 39460 16838
rect 39220 16816 39516 16836
rect 39220 15804 39516 15824
rect 39276 15802 39300 15804
rect 39356 15802 39380 15804
rect 39436 15802 39460 15804
rect 39298 15750 39300 15802
rect 39362 15750 39374 15802
rect 39436 15750 39438 15802
rect 39276 15748 39300 15750
rect 39356 15748 39380 15750
rect 39436 15748 39460 15750
rect 39220 15728 39516 15748
rect 39220 14716 39516 14736
rect 39276 14714 39300 14716
rect 39356 14714 39380 14716
rect 39436 14714 39460 14716
rect 39298 14662 39300 14714
rect 39362 14662 39374 14714
rect 39436 14662 39438 14714
rect 39276 14660 39300 14662
rect 39356 14660 39380 14662
rect 39436 14660 39460 14662
rect 39220 14640 39516 14660
rect 39220 13628 39516 13648
rect 39276 13626 39300 13628
rect 39356 13626 39380 13628
rect 39436 13626 39460 13628
rect 39298 13574 39300 13626
rect 39362 13574 39374 13626
rect 39436 13574 39438 13626
rect 39276 13572 39300 13574
rect 39356 13572 39380 13574
rect 39436 13572 39460 13574
rect 39220 13552 39516 13572
rect 39212 13184 39264 13190
rect 39210 13152 39212 13161
rect 39264 13152 39266 13161
rect 39210 13087 39266 13096
rect 39592 12646 39620 31962
rect 39948 31952 40000 31958
rect 39948 31894 40000 31900
rect 39960 26450 39988 31894
rect 40328 30870 40356 44678
rect 40316 30864 40368 30870
rect 40316 30806 40368 30812
rect 39948 26444 40000 26450
rect 39948 26386 40000 26392
rect 39672 23180 39724 23186
rect 39672 23122 39724 23128
rect 39684 22778 39712 23122
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 39764 21480 39816 21486
rect 39764 21422 39816 21428
rect 39776 16574 39804 21422
rect 39856 21412 39908 21418
rect 39856 21354 39908 21360
rect 39684 16546 39804 16574
rect 39684 13190 39712 16546
rect 39764 14000 39816 14006
rect 39764 13942 39816 13948
rect 39776 13870 39804 13942
rect 39764 13864 39816 13870
rect 39764 13806 39816 13812
rect 39672 13184 39724 13190
rect 39672 13126 39724 13132
rect 39120 12640 39172 12646
rect 39120 12582 39172 12588
rect 39580 12640 39632 12646
rect 39580 12582 39632 12588
rect 39132 12434 39160 12582
rect 39220 12540 39516 12560
rect 39276 12538 39300 12540
rect 39356 12538 39380 12540
rect 39436 12538 39460 12540
rect 39298 12486 39300 12538
rect 39362 12486 39374 12538
rect 39436 12486 39438 12538
rect 39276 12484 39300 12486
rect 39356 12484 39380 12486
rect 39436 12484 39460 12486
rect 39220 12464 39516 12484
rect 39684 12458 39712 13126
rect 39776 12481 39804 13806
rect 38948 12406 39160 12434
rect 39592 12430 39712 12458
rect 39762 12472 39818 12481
rect 38844 5160 38896 5166
rect 38844 5102 38896 5108
rect 38844 4548 38896 4554
rect 38844 4490 38896 4496
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 38568 3732 38620 3738
rect 38568 3674 38620 3680
rect 38580 2774 38608 3674
rect 38658 3632 38714 3641
rect 38658 3567 38714 3576
rect 38672 3369 38700 3567
rect 38764 3398 38792 3878
rect 38752 3392 38804 3398
rect 38658 3360 38714 3369
rect 38752 3334 38804 3340
rect 38658 3295 38714 3304
rect 38488 2746 38608 2774
rect 38488 1426 38516 2746
rect 38750 2544 38806 2553
rect 38750 2479 38806 2488
rect 38568 2032 38620 2038
rect 38568 1974 38620 1980
rect 38658 2000 38714 2009
rect 38476 1420 38528 1426
rect 38476 1362 38528 1368
rect 38580 800 38608 1974
rect 38658 1935 38714 1944
rect 38672 800 38700 1935
rect 38764 1306 38792 2479
rect 38856 1442 38884 4490
rect 38948 2582 38976 12406
rect 39120 12096 39172 12102
rect 39120 12038 39172 12044
rect 39028 10464 39080 10470
rect 39028 10406 39080 10412
rect 39040 9194 39068 10406
rect 39132 9518 39160 12038
rect 39220 11452 39516 11472
rect 39276 11450 39300 11452
rect 39356 11450 39380 11452
rect 39436 11450 39460 11452
rect 39298 11398 39300 11450
rect 39362 11398 39374 11450
rect 39436 11398 39438 11450
rect 39276 11396 39300 11398
rect 39356 11396 39380 11398
rect 39436 11396 39460 11398
rect 39220 11376 39516 11396
rect 39220 10364 39516 10384
rect 39276 10362 39300 10364
rect 39356 10362 39380 10364
rect 39436 10362 39460 10364
rect 39298 10310 39300 10362
rect 39362 10310 39374 10362
rect 39436 10310 39438 10362
rect 39276 10308 39300 10310
rect 39356 10308 39380 10310
rect 39436 10308 39460 10310
rect 39220 10288 39516 10308
rect 39396 10192 39448 10198
rect 39396 10134 39448 10140
rect 39408 9518 39436 10134
rect 39488 9920 39540 9926
rect 39488 9862 39540 9868
rect 39120 9512 39172 9518
rect 39120 9454 39172 9460
rect 39396 9512 39448 9518
rect 39500 9489 39528 9862
rect 39396 9454 39448 9460
rect 39486 9480 39542 9489
rect 39486 9415 39542 9424
rect 39220 9276 39516 9296
rect 39276 9274 39300 9276
rect 39356 9274 39380 9276
rect 39436 9274 39460 9276
rect 39298 9222 39300 9274
rect 39362 9222 39374 9274
rect 39436 9222 39438 9274
rect 39276 9220 39300 9222
rect 39356 9220 39380 9222
rect 39436 9220 39460 9222
rect 39220 9200 39516 9220
rect 39040 9166 39160 9194
rect 39026 9072 39082 9081
rect 39026 9007 39028 9016
rect 39080 9007 39082 9016
rect 39028 8978 39080 8984
rect 39028 8016 39080 8022
rect 39028 7958 39080 7964
rect 39040 4729 39068 7958
rect 39132 7274 39160 9166
rect 39394 8528 39450 8537
rect 39394 8463 39450 8472
rect 39408 8430 39436 8463
rect 39396 8424 39448 8430
rect 39396 8366 39448 8372
rect 39220 8188 39516 8208
rect 39276 8186 39300 8188
rect 39356 8186 39380 8188
rect 39436 8186 39460 8188
rect 39298 8134 39300 8186
rect 39362 8134 39374 8186
rect 39436 8134 39438 8186
rect 39276 8132 39300 8134
rect 39356 8132 39380 8134
rect 39436 8132 39460 8134
rect 39220 8112 39516 8132
rect 39120 7268 39172 7274
rect 39120 7210 39172 7216
rect 39220 7100 39516 7120
rect 39276 7098 39300 7100
rect 39356 7098 39380 7100
rect 39436 7098 39460 7100
rect 39298 7046 39300 7098
rect 39362 7046 39374 7098
rect 39436 7046 39438 7098
rect 39276 7044 39300 7046
rect 39356 7044 39380 7046
rect 39436 7044 39460 7046
rect 39220 7024 39516 7044
rect 39220 6012 39516 6032
rect 39276 6010 39300 6012
rect 39356 6010 39380 6012
rect 39436 6010 39460 6012
rect 39298 5958 39300 6010
rect 39362 5958 39374 6010
rect 39436 5958 39438 6010
rect 39276 5956 39300 5958
rect 39356 5956 39380 5958
rect 39436 5956 39460 5958
rect 39220 5936 39516 5956
rect 39210 5672 39266 5681
rect 39210 5607 39212 5616
rect 39264 5607 39266 5616
rect 39212 5578 39264 5584
rect 39220 4924 39516 4944
rect 39276 4922 39300 4924
rect 39356 4922 39380 4924
rect 39436 4922 39460 4924
rect 39298 4870 39300 4922
rect 39362 4870 39374 4922
rect 39436 4870 39438 4922
rect 39276 4868 39300 4870
rect 39356 4868 39380 4870
rect 39436 4868 39460 4870
rect 39220 4848 39516 4868
rect 39026 4720 39082 4729
rect 39592 4706 39620 12430
rect 39762 12407 39818 12416
rect 39764 12232 39816 12238
rect 39762 12200 39764 12209
rect 39816 12200 39818 12209
rect 39868 12170 39896 21354
rect 40040 13456 40092 13462
rect 40040 13398 40092 13404
rect 40052 13326 40080 13398
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 40132 13320 40184 13326
rect 40132 13262 40184 13268
rect 39946 13016 40002 13025
rect 39946 12951 39948 12960
rect 40000 12951 40002 12960
rect 39948 12922 40000 12928
rect 39762 12135 39818 12144
rect 39856 12164 39908 12170
rect 39856 12106 39908 12112
rect 39764 12096 39816 12102
rect 39764 12038 39816 12044
rect 39670 11384 39726 11393
rect 39670 11319 39726 11328
rect 39684 11121 39712 11319
rect 39776 11218 39804 12038
rect 39764 11212 39816 11218
rect 39764 11154 39816 11160
rect 39670 11112 39726 11121
rect 39670 11047 39726 11056
rect 39764 11076 39816 11082
rect 39764 11018 39816 11024
rect 39672 11008 39724 11014
rect 39672 10950 39724 10956
rect 39684 10198 39712 10950
rect 39672 10192 39724 10198
rect 39672 10134 39724 10140
rect 39776 9874 39804 11018
rect 39684 9846 39804 9874
rect 39684 7954 39712 9846
rect 39764 9716 39816 9722
rect 39764 9658 39816 9664
rect 39672 7948 39724 7954
rect 39672 7890 39724 7896
rect 39672 7744 39724 7750
rect 39672 7686 39724 7692
rect 39684 7546 39712 7686
rect 39672 7540 39724 7546
rect 39672 7482 39724 7488
rect 39670 7032 39726 7041
rect 39670 6967 39726 6976
rect 39026 4655 39082 4664
rect 39224 4678 39620 4706
rect 39684 4690 39712 6967
rect 39776 6458 39804 9658
rect 39868 8945 39896 12106
rect 39854 8936 39910 8945
rect 39854 8871 39910 8880
rect 39856 8832 39908 8838
rect 39856 8774 39908 8780
rect 39868 6798 39896 8774
rect 39856 6792 39908 6798
rect 39856 6734 39908 6740
rect 39854 6624 39910 6633
rect 39854 6559 39910 6568
rect 39868 6458 39896 6559
rect 39764 6452 39816 6458
rect 39764 6394 39816 6400
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 39856 6316 39908 6322
rect 39856 6258 39908 6264
rect 39868 5574 39896 6258
rect 39856 5568 39908 5574
rect 39856 5510 39908 5516
rect 39764 5160 39816 5166
rect 39764 5102 39816 5108
rect 39672 4684 39724 4690
rect 39120 4208 39172 4214
rect 39120 4150 39172 4156
rect 39026 3768 39082 3777
rect 39026 3703 39082 3712
rect 39040 3602 39068 3703
rect 39028 3596 39080 3602
rect 39028 3538 39080 3544
rect 39132 3466 39160 4150
rect 39224 4078 39252 4678
rect 39672 4626 39724 4632
rect 39670 4584 39726 4593
rect 39670 4519 39726 4528
rect 39394 4176 39450 4185
rect 39394 4111 39450 4120
rect 39408 4078 39436 4111
rect 39212 4072 39264 4078
rect 39212 4014 39264 4020
rect 39396 4072 39448 4078
rect 39396 4014 39448 4020
rect 39684 4010 39712 4519
rect 39672 4004 39724 4010
rect 39672 3946 39724 3952
rect 39220 3836 39516 3856
rect 39276 3834 39300 3836
rect 39356 3834 39380 3836
rect 39436 3834 39460 3836
rect 39298 3782 39300 3834
rect 39362 3782 39374 3834
rect 39436 3782 39438 3834
rect 39276 3780 39300 3782
rect 39356 3780 39380 3782
rect 39436 3780 39460 3782
rect 39220 3760 39516 3780
rect 39776 3652 39804 5102
rect 39854 4720 39910 4729
rect 39854 4655 39856 4664
rect 39908 4655 39910 4664
rect 39856 4626 39908 4632
rect 39592 3624 39804 3652
rect 39212 3596 39264 3602
rect 39212 3538 39264 3544
rect 39224 3466 39252 3538
rect 39120 3460 39172 3466
rect 39120 3402 39172 3408
rect 39212 3460 39264 3466
rect 39212 3402 39264 3408
rect 39488 3460 39540 3466
rect 39488 3402 39540 3408
rect 39500 3369 39528 3402
rect 39210 3360 39266 3369
rect 39210 3295 39266 3304
rect 39486 3360 39542 3369
rect 39486 3295 39542 3304
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 38936 2576 38988 2582
rect 38936 2518 38988 2524
rect 38856 1414 38976 1442
rect 38764 1278 38884 1306
rect 38856 800 38884 1278
rect 38948 800 38976 1414
rect 39132 800 39160 2994
rect 39224 2990 39252 3295
rect 39212 2984 39264 2990
rect 39212 2926 39264 2932
rect 39220 2748 39516 2768
rect 39276 2746 39300 2748
rect 39356 2746 39380 2748
rect 39436 2746 39460 2748
rect 39298 2694 39300 2746
rect 39362 2694 39374 2746
rect 39436 2694 39438 2746
rect 39276 2692 39300 2694
rect 39356 2692 39380 2694
rect 39436 2692 39460 2694
rect 39220 2672 39516 2692
rect 39592 2530 39620 3624
rect 39868 3584 39896 4626
rect 39408 2502 39620 2530
rect 39684 3556 39896 3584
rect 39210 2272 39266 2281
rect 39210 2207 39266 2216
rect 39224 800 39252 2207
rect 39408 800 39436 2502
rect 39684 2106 39712 3556
rect 39762 3496 39818 3505
rect 39762 3431 39818 3440
rect 39776 3126 39804 3431
rect 39856 3392 39908 3398
rect 39856 3334 39908 3340
rect 39764 3120 39816 3126
rect 39764 3062 39816 3068
rect 39868 2666 39896 3334
rect 39960 2990 39988 12922
rect 40144 12434 40172 13262
rect 40316 13184 40368 13190
rect 40316 13126 40368 13132
rect 40328 12850 40356 13126
rect 40316 12844 40368 12850
rect 40316 12786 40368 12792
rect 40144 12406 40264 12434
rect 40132 11552 40184 11558
rect 40132 11494 40184 11500
rect 40040 11076 40092 11082
rect 40040 11018 40092 11024
rect 40052 8430 40080 11018
rect 40144 10577 40172 11494
rect 40130 10568 40186 10577
rect 40130 10503 40186 10512
rect 40132 10464 40184 10470
rect 40132 10406 40184 10412
rect 40040 8424 40092 8430
rect 40040 8366 40092 8372
rect 40052 5545 40080 8366
rect 40144 7410 40172 10406
rect 40132 7404 40184 7410
rect 40132 7346 40184 7352
rect 40132 7268 40184 7274
rect 40132 7210 40184 7216
rect 40144 6934 40172 7210
rect 40132 6928 40184 6934
rect 40132 6870 40184 6876
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 40038 5536 40094 5545
rect 40038 5471 40094 5480
rect 40144 4282 40172 6734
rect 40236 5370 40264 12406
rect 40316 12096 40368 12102
rect 40316 12038 40368 12044
rect 40328 9518 40356 12038
rect 40316 9512 40368 9518
rect 40316 9454 40368 9460
rect 40316 9376 40368 9382
rect 40316 9318 40368 9324
rect 40328 8430 40356 9318
rect 40316 8424 40368 8430
rect 40316 8366 40368 8372
rect 40316 8084 40368 8090
rect 40316 8026 40368 8032
rect 40328 7478 40356 8026
rect 40316 7472 40368 7478
rect 40316 7414 40368 7420
rect 40316 7336 40368 7342
rect 40316 7278 40368 7284
rect 40328 7002 40356 7278
rect 40316 6996 40368 7002
rect 40316 6938 40368 6944
rect 40316 6656 40368 6662
rect 40420 6633 40448 47602
rect 40776 47184 40828 47190
rect 40776 47126 40828 47132
rect 40788 38554 40816 47126
rect 40776 38548 40828 38554
rect 40776 38490 40828 38496
rect 40960 38208 41012 38214
rect 40960 38150 41012 38156
rect 40972 38010 41000 38150
rect 40960 38004 41012 38010
rect 40960 37946 41012 37952
rect 40684 37800 40736 37806
rect 40684 37742 40736 37748
rect 40696 13462 40724 37742
rect 41236 32428 41288 32434
rect 41236 32370 41288 32376
rect 40684 13456 40736 13462
rect 40684 13398 40736 13404
rect 41144 13456 41196 13462
rect 41144 13398 41196 13404
rect 41156 13190 41184 13398
rect 41144 13184 41196 13190
rect 41144 13126 41196 13132
rect 40960 12912 41012 12918
rect 40960 12854 41012 12860
rect 40592 12776 40644 12782
rect 40592 12718 40644 12724
rect 40500 11552 40552 11558
rect 40500 11494 40552 11500
rect 40512 9382 40540 11494
rect 40500 9376 40552 9382
rect 40500 9318 40552 9324
rect 40498 9208 40554 9217
rect 40498 9143 40554 9152
rect 40512 9042 40540 9143
rect 40500 9036 40552 9042
rect 40500 8978 40552 8984
rect 40500 8560 40552 8566
rect 40500 8502 40552 8508
rect 40316 6598 40368 6604
rect 40406 6624 40462 6633
rect 40328 5778 40356 6598
rect 40406 6559 40462 6568
rect 40512 6202 40540 8502
rect 40420 6174 40540 6202
rect 40316 5772 40368 5778
rect 40316 5714 40368 5720
rect 40316 5636 40368 5642
rect 40316 5578 40368 5584
rect 40224 5364 40276 5370
rect 40224 5306 40276 5312
rect 40236 5098 40264 5306
rect 40224 5092 40276 5098
rect 40224 5034 40276 5040
rect 40224 4548 40276 4554
rect 40224 4490 40276 4496
rect 40132 4276 40184 4282
rect 40132 4218 40184 4224
rect 40132 4072 40184 4078
rect 40132 4014 40184 4020
rect 40040 4004 40092 4010
rect 40040 3946 40092 3952
rect 40052 3194 40080 3946
rect 40040 3188 40092 3194
rect 40040 3130 40092 3136
rect 40144 3058 40172 4014
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 40132 2848 40184 2854
rect 40130 2816 40132 2825
rect 40184 2816 40186 2825
rect 40130 2751 40186 2760
rect 39868 2638 39988 2666
rect 39856 2576 39908 2582
rect 39856 2518 39908 2524
rect 39672 2100 39724 2106
rect 39672 2042 39724 2048
rect 39486 1320 39542 1329
rect 39486 1255 39542 1264
rect 39500 800 39528 1255
rect 39868 1170 39896 2518
rect 39960 2106 39988 2638
rect 39948 2100 40000 2106
rect 39948 2042 40000 2048
rect 39948 1828 40000 1834
rect 39948 1770 40000 1776
rect 39684 1142 39896 1170
rect 39684 800 39712 1142
rect 39764 1080 39816 1086
rect 39764 1022 39816 1028
rect 39776 800 39804 1022
rect 39960 800 39988 1770
rect 40040 1420 40092 1426
rect 40040 1362 40092 1368
rect 40052 800 40080 1362
rect 40236 800 40264 4490
rect 40328 4078 40356 5578
rect 40316 4072 40368 4078
rect 40316 4014 40368 4020
rect 40316 3188 40368 3194
rect 40316 3130 40368 3136
rect 40328 2582 40356 3130
rect 40316 2576 40368 2582
rect 40316 2518 40368 2524
rect 40420 800 40448 6174
rect 40498 6080 40554 6089
rect 40498 6015 40554 6024
rect 40512 3924 40540 6015
rect 40604 4078 40632 12718
rect 40684 12708 40736 12714
rect 40684 12650 40736 12656
rect 40592 4072 40644 4078
rect 40592 4014 40644 4020
rect 40512 3896 40632 3924
rect 40498 3088 40554 3097
rect 40498 3023 40500 3032
rect 40552 3023 40554 3032
rect 40500 2994 40552 3000
rect 40500 2916 40552 2922
rect 40500 2858 40552 2864
rect 40512 800 40540 2858
rect 40604 1290 40632 3896
rect 40696 3670 40724 12650
rect 40868 12640 40920 12646
rect 40866 12608 40868 12617
rect 40920 12608 40922 12617
rect 40866 12543 40922 12552
rect 40972 12102 41000 12854
rect 40960 12096 41012 12102
rect 40960 12038 41012 12044
rect 40868 11076 40920 11082
rect 40868 11018 40920 11024
rect 40776 10464 40828 10470
rect 40776 10406 40828 10412
rect 40788 7342 40816 10406
rect 40880 10033 40908 11018
rect 40866 10024 40922 10033
rect 40866 9959 40922 9968
rect 40868 9920 40920 9926
rect 40868 9862 40920 9868
rect 40776 7336 40828 7342
rect 40776 7278 40828 7284
rect 40776 7200 40828 7206
rect 40776 7142 40828 7148
rect 40788 5642 40816 7142
rect 40880 6254 40908 9862
rect 40868 6248 40920 6254
rect 40868 6190 40920 6196
rect 40776 5636 40828 5642
rect 40776 5578 40828 5584
rect 40684 3664 40736 3670
rect 40684 3606 40736 3612
rect 40868 3596 40920 3602
rect 40868 3538 40920 3544
rect 40682 3088 40738 3097
rect 40682 3023 40738 3032
rect 40776 3052 40828 3058
rect 40696 2990 40724 3023
rect 40776 2994 40828 3000
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40788 1442 40816 2994
rect 40696 1414 40816 1442
rect 40880 1442 40908 3538
rect 40972 2582 41000 12038
rect 41052 11552 41104 11558
rect 41052 11494 41104 11500
rect 41064 8974 41092 11494
rect 41248 9994 41276 32370
rect 41328 19168 41380 19174
rect 41328 19110 41380 19116
rect 41236 9988 41288 9994
rect 41236 9930 41288 9936
rect 41144 9920 41196 9926
rect 41144 9862 41196 9868
rect 41052 8968 41104 8974
rect 41052 8910 41104 8916
rect 41052 8628 41104 8634
rect 41052 8570 41104 8576
rect 41064 4690 41092 8570
rect 41156 6866 41184 9862
rect 41340 9722 41368 19110
rect 41524 14521 41552 66438
rect 44220 66396 44516 66416
rect 44276 66394 44300 66396
rect 44356 66394 44380 66396
rect 44436 66394 44460 66396
rect 44298 66342 44300 66394
rect 44362 66342 44374 66394
rect 44436 66342 44438 66394
rect 44276 66340 44300 66342
rect 44356 66340 44380 66342
rect 44436 66340 44460 66342
rect 44220 66320 44516 66340
rect 49220 65852 49516 65872
rect 49276 65850 49300 65852
rect 49356 65850 49380 65852
rect 49436 65850 49460 65852
rect 49298 65798 49300 65850
rect 49362 65798 49374 65850
rect 49436 65798 49438 65850
rect 49276 65796 49300 65798
rect 49356 65796 49380 65798
rect 49436 65796 49460 65798
rect 49220 65776 49516 65796
rect 44220 65308 44516 65328
rect 44276 65306 44300 65308
rect 44356 65306 44380 65308
rect 44436 65306 44460 65308
rect 44298 65254 44300 65306
rect 44362 65254 44374 65306
rect 44436 65254 44438 65306
rect 44276 65252 44300 65254
rect 44356 65252 44380 65254
rect 44436 65252 44460 65254
rect 44220 65232 44516 65252
rect 49220 64764 49516 64784
rect 49276 64762 49300 64764
rect 49356 64762 49380 64764
rect 49436 64762 49460 64764
rect 49298 64710 49300 64762
rect 49362 64710 49374 64762
rect 49436 64710 49438 64762
rect 49276 64708 49300 64710
rect 49356 64708 49380 64710
rect 49436 64708 49460 64710
rect 49220 64688 49516 64708
rect 44220 64220 44516 64240
rect 44276 64218 44300 64220
rect 44356 64218 44380 64220
rect 44436 64218 44460 64220
rect 44298 64166 44300 64218
rect 44362 64166 44374 64218
rect 44436 64166 44438 64218
rect 44276 64164 44300 64166
rect 44356 64164 44380 64166
rect 44436 64164 44460 64166
rect 44220 64144 44516 64164
rect 49220 63676 49516 63696
rect 49276 63674 49300 63676
rect 49356 63674 49380 63676
rect 49436 63674 49460 63676
rect 49298 63622 49300 63674
rect 49362 63622 49374 63674
rect 49436 63622 49438 63674
rect 49276 63620 49300 63622
rect 49356 63620 49380 63622
rect 49436 63620 49460 63622
rect 49220 63600 49516 63620
rect 50068 63232 50120 63238
rect 50068 63174 50120 63180
rect 44220 63132 44516 63152
rect 44276 63130 44300 63132
rect 44356 63130 44380 63132
rect 44436 63130 44460 63132
rect 44298 63078 44300 63130
rect 44362 63078 44374 63130
rect 44436 63078 44438 63130
rect 44276 63076 44300 63078
rect 44356 63076 44380 63078
rect 44436 63076 44460 63078
rect 44220 63056 44516 63076
rect 48964 62960 49016 62966
rect 48964 62902 49016 62908
rect 48976 62422 49004 62902
rect 49148 62824 49200 62830
rect 49148 62766 49200 62772
rect 48964 62416 49016 62422
rect 48964 62358 49016 62364
rect 44220 62044 44516 62064
rect 44276 62042 44300 62044
rect 44356 62042 44380 62044
rect 44436 62042 44460 62044
rect 44298 61990 44300 62042
rect 44362 61990 44374 62042
rect 44436 61990 44438 62042
rect 44276 61988 44300 61990
rect 44356 61988 44380 61990
rect 44436 61988 44460 61990
rect 44220 61968 44516 61988
rect 44220 60956 44516 60976
rect 44276 60954 44300 60956
rect 44356 60954 44380 60956
rect 44436 60954 44460 60956
rect 44298 60902 44300 60954
rect 44362 60902 44374 60954
rect 44436 60902 44438 60954
rect 44276 60900 44300 60902
rect 44356 60900 44380 60902
rect 44436 60900 44460 60902
rect 44220 60880 44516 60900
rect 44088 60104 44140 60110
rect 44088 60046 44140 60052
rect 43996 58948 44048 58954
rect 43996 58890 44048 58896
rect 42524 58676 42576 58682
rect 42524 58618 42576 58624
rect 42536 58342 42564 58618
rect 44008 58546 44036 58890
rect 44100 58546 44128 60046
rect 47400 59968 47452 59974
rect 47400 59910 47452 59916
rect 44220 59868 44516 59888
rect 44276 59866 44300 59868
rect 44356 59866 44380 59868
rect 44436 59866 44460 59868
rect 44298 59814 44300 59866
rect 44362 59814 44374 59866
rect 44436 59814 44438 59866
rect 44276 59812 44300 59814
rect 44356 59812 44380 59814
rect 44436 59812 44460 59814
rect 44220 59792 44516 59812
rect 44220 58780 44516 58800
rect 44276 58778 44300 58780
rect 44356 58778 44380 58780
rect 44436 58778 44460 58780
rect 44298 58726 44300 58778
rect 44362 58726 44374 58778
rect 44436 58726 44438 58778
rect 44276 58724 44300 58726
rect 44356 58724 44380 58726
rect 44436 58724 44460 58726
rect 44220 58704 44516 58724
rect 44180 58608 44232 58614
rect 44456 58608 44508 58614
rect 44232 58556 44456 58562
rect 44180 58550 44508 58556
rect 43996 58540 44048 58546
rect 43996 58482 44048 58488
rect 44088 58540 44140 58546
rect 44192 58534 44496 58550
rect 44088 58482 44140 58488
rect 43260 58472 43312 58478
rect 43260 58414 43312 58420
rect 43272 58342 43300 58414
rect 42524 58336 42576 58342
rect 42524 58278 42576 58284
rect 43260 58336 43312 58342
rect 43260 58278 43312 58284
rect 43812 58336 43864 58342
rect 43812 58278 43864 58284
rect 42340 55412 42392 55418
rect 42340 55354 42392 55360
rect 41696 55276 41748 55282
rect 41696 55218 41748 55224
rect 41604 41608 41656 41614
rect 41604 41550 41656 41556
rect 41616 36174 41644 41550
rect 41604 36168 41656 36174
rect 41604 36110 41656 36116
rect 41616 35494 41644 36110
rect 41604 35488 41656 35494
rect 41604 35430 41656 35436
rect 41510 14512 41566 14521
rect 41510 14447 41566 14456
rect 41420 11076 41472 11082
rect 41420 11018 41472 11024
rect 41328 9716 41380 9722
rect 41328 9658 41380 9664
rect 41236 9512 41288 9518
rect 41236 9454 41288 9460
rect 41248 7206 41276 9454
rect 41432 8430 41460 11018
rect 41512 10464 41564 10470
rect 41512 10406 41564 10412
rect 41420 8424 41472 8430
rect 41420 8366 41472 8372
rect 41328 8356 41380 8362
rect 41328 8298 41380 8304
rect 41340 8265 41368 8298
rect 41420 8288 41472 8294
rect 41326 8256 41382 8265
rect 41420 8230 41472 8236
rect 41326 8191 41382 8200
rect 41432 7954 41460 8230
rect 41420 7948 41472 7954
rect 41420 7890 41472 7896
rect 41236 7200 41288 7206
rect 41432 7188 41460 7890
rect 41524 7342 41552 10406
rect 41708 10062 41736 55218
rect 42064 36168 42116 36174
rect 42064 36110 42116 36116
rect 42076 36038 42104 36110
rect 42064 36032 42116 36038
rect 42064 35974 42116 35980
rect 41972 13184 42024 13190
rect 41972 13126 42024 13132
rect 41984 10849 42012 13126
rect 42156 11892 42208 11898
rect 42156 11834 42208 11840
rect 42168 11082 42196 11834
rect 42248 11620 42300 11626
rect 42248 11562 42300 11568
rect 42064 11076 42116 11082
rect 42064 11018 42116 11024
rect 42156 11076 42208 11082
rect 42156 11018 42208 11024
rect 41970 10840 42026 10849
rect 41970 10775 42026 10784
rect 41880 10464 41932 10470
rect 41880 10406 41932 10412
rect 41696 10056 41748 10062
rect 41696 9998 41748 10004
rect 41696 9920 41748 9926
rect 41696 9862 41748 9868
rect 41604 9376 41656 9382
rect 41604 9318 41656 9324
rect 41512 7336 41564 7342
rect 41512 7278 41564 7284
rect 41432 7160 41552 7188
rect 41236 7142 41288 7148
rect 41248 7002 41460 7018
rect 41248 6996 41472 7002
rect 41248 6990 41420 6996
rect 41144 6860 41196 6866
rect 41144 6802 41196 6808
rect 41144 6112 41196 6118
rect 41142 6080 41144 6089
rect 41196 6080 41198 6089
rect 41142 6015 41198 6024
rect 41052 4684 41104 4690
rect 41052 4626 41104 4632
rect 41142 4584 41198 4593
rect 41052 4548 41104 4554
rect 41142 4519 41198 4528
rect 41052 4490 41104 4496
rect 41064 2961 41092 4490
rect 41050 2952 41106 2961
rect 41050 2887 41106 2896
rect 40960 2576 41012 2582
rect 40960 2518 41012 2524
rect 41052 2100 41104 2106
rect 41052 2042 41104 2048
rect 40880 1414 41000 1442
rect 40592 1284 40644 1290
rect 40592 1226 40644 1232
rect 40696 800 40724 1414
rect 40776 1284 40828 1290
rect 40776 1226 40828 1232
rect 40788 800 40816 1226
rect 40972 800 41000 1414
rect 41064 800 41092 2042
rect 41156 1426 41184 4519
rect 41144 1420 41196 1426
rect 41144 1362 41196 1368
rect 41248 800 41276 6990
rect 41420 6938 41472 6944
rect 41420 6860 41472 6866
rect 41420 6802 41472 6808
rect 41328 5772 41380 5778
rect 41328 5714 41380 5720
rect 41340 4554 41368 5714
rect 41328 4548 41380 4554
rect 41328 4490 41380 4496
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 41340 800 41368 3334
rect 41432 3194 41460 6802
rect 41524 6100 41552 7160
rect 41616 6254 41644 9318
rect 41708 8294 41736 9862
rect 41788 8832 41840 8838
rect 41788 8774 41840 8780
rect 41696 8288 41748 8294
rect 41696 8230 41748 8236
rect 41696 7336 41748 7342
rect 41696 7278 41748 7284
rect 41708 6497 41736 7278
rect 41694 6488 41750 6497
rect 41694 6423 41750 6432
rect 41604 6248 41656 6254
rect 41604 6190 41656 6196
rect 41524 6072 41644 6100
rect 41512 3936 41564 3942
rect 41512 3878 41564 3884
rect 41420 3188 41472 3194
rect 41420 3130 41472 3136
rect 41418 3088 41474 3097
rect 41418 3023 41474 3032
rect 41432 2990 41460 3023
rect 41420 2984 41472 2990
rect 41420 2926 41472 2932
rect 41524 800 41552 3878
rect 41616 2553 41644 6072
rect 41800 5778 41828 8774
rect 41892 7954 41920 10406
rect 41880 7948 41932 7954
rect 41880 7890 41932 7896
rect 41892 7818 41920 7890
rect 41880 7812 41932 7818
rect 41880 7754 41932 7760
rect 41788 5772 41840 5778
rect 41788 5714 41840 5720
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41708 3369 41736 5510
rect 41800 5273 41828 5714
rect 41786 5264 41842 5273
rect 41786 5199 41842 5208
rect 41984 5166 42012 10775
rect 42076 9518 42104 11018
rect 42156 9920 42208 9926
rect 42156 9862 42208 9868
rect 42064 9512 42116 9518
rect 42064 9454 42116 9460
rect 42064 9376 42116 9382
rect 42064 9318 42116 9324
rect 42076 6254 42104 9318
rect 42168 6866 42196 9862
rect 42156 6860 42208 6866
rect 42156 6802 42208 6808
rect 42064 6248 42116 6254
rect 42064 6190 42116 6196
rect 42076 5914 42104 6190
rect 42064 5908 42116 5914
rect 42064 5850 42116 5856
rect 42156 5636 42208 5642
rect 42156 5578 42208 5584
rect 41972 5160 42024 5166
rect 41972 5102 42024 5108
rect 41788 4276 41840 4282
rect 41788 4218 41840 4224
rect 41694 3360 41750 3369
rect 41694 3295 41750 3304
rect 41800 3210 41828 4218
rect 42064 4140 42116 4146
rect 42064 4082 42116 4088
rect 42076 3602 42104 4082
rect 42168 3670 42196 5578
rect 42260 4010 42288 11562
rect 42352 11121 42380 55354
rect 42432 32020 42484 32026
rect 42432 31962 42484 31968
rect 42444 31754 42472 31962
rect 42432 31748 42484 31754
rect 42432 31690 42484 31696
rect 42432 30388 42484 30394
rect 42432 30330 42484 30336
rect 42444 11626 42472 30330
rect 42536 25770 42564 58278
rect 43272 53650 43300 58278
rect 43444 57792 43496 57798
rect 43444 57734 43496 57740
rect 43260 53644 43312 53650
rect 43260 53586 43312 53592
rect 43456 53446 43484 57734
rect 43444 53440 43496 53446
rect 43444 53382 43496 53388
rect 43720 38548 43772 38554
rect 43720 38490 43772 38496
rect 43168 36032 43220 36038
rect 43168 35974 43220 35980
rect 42616 26580 42668 26586
rect 42616 26522 42668 26528
rect 42628 26450 42656 26522
rect 42616 26444 42668 26450
rect 42616 26386 42668 26392
rect 42524 25764 42576 25770
rect 42524 25706 42576 25712
rect 42524 17060 42576 17066
rect 42524 17002 42576 17008
rect 42432 11620 42484 11626
rect 42432 11562 42484 11568
rect 42432 11144 42484 11150
rect 42338 11112 42394 11121
rect 42536 11132 42564 17002
rect 43180 13326 43208 35974
rect 43628 27668 43680 27674
rect 43628 27610 43680 27616
rect 43168 13320 43220 13326
rect 43168 13262 43220 13268
rect 42616 12912 42668 12918
rect 42616 12854 42668 12860
rect 42628 12714 42656 12854
rect 42616 12708 42668 12714
rect 42616 12650 42668 12656
rect 42708 12096 42760 12102
rect 42708 12038 42760 12044
rect 43260 12096 43312 12102
rect 43260 12038 43312 12044
rect 42720 11234 42748 12038
rect 42892 11552 42944 11558
rect 42892 11494 42944 11500
rect 42720 11206 42840 11234
rect 42484 11104 42564 11132
rect 42706 11112 42762 11121
rect 42432 11086 42484 11092
rect 42338 11047 42394 11056
rect 42340 11008 42392 11014
rect 42340 10950 42392 10956
rect 42352 8945 42380 10950
rect 42338 8936 42394 8945
rect 42338 8871 42394 8880
rect 42340 8832 42392 8838
rect 42340 8774 42392 8780
rect 42352 5953 42380 8774
rect 42338 5944 42394 5953
rect 42338 5879 42394 5888
rect 42352 5778 42380 5879
rect 42340 5772 42392 5778
rect 42340 5714 42392 5720
rect 42340 5296 42392 5302
rect 42340 5238 42392 5244
rect 42248 4004 42300 4010
rect 42248 3946 42300 3952
rect 42352 3720 42380 5238
rect 42444 4078 42472 11086
rect 42616 11076 42668 11082
rect 42706 11047 42708 11056
rect 42616 11018 42668 11024
rect 42760 11047 42762 11056
rect 42708 11018 42760 11024
rect 42524 10600 42576 10606
rect 42524 10542 42576 10548
rect 42536 10062 42564 10542
rect 42524 10056 42576 10062
rect 42524 9998 42576 10004
rect 42536 5098 42564 9998
rect 42628 8430 42656 11018
rect 42812 10962 42840 11206
rect 42720 10934 42840 10962
rect 42616 8424 42668 8430
rect 42616 8366 42668 8372
rect 42720 6066 42748 10934
rect 42800 9920 42852 9926
rect 42800 9862 42852 9868
rect 42812 7954 42840 9862
rect 42904 9081 42932 11494
rect 42984 10464 43036 10470
rect 42984 10406 43036 10412
rect 42890 9072 42946 9081
rect 42890 9007 42946 9016
rect 42892 8832 42944 8838
rect 42892 8774 42944 8780
rect 42800 7948 42852 7954
rect 42800 7890 42852 7896
rect 42904 6984 42932 8774
rect 42996 8090 43024 10406
rect 43168 9512 43220 9518
rect 43168 9454 43220 9460
rect 43076 9376 43128 9382
rect 43076 9318 43128 9324
rect 42984 8084 43036 8090
rect 42984 8026 43036 8032
rect 42996 7954 43024 8026
rect 42984 7948 43036 7954
rect 42984 7890 43036 7896
rect 43088 7342 43116 9318
rect 43076 7336 43128 7342
rect 43076 7278 43128 7284
rect 42812 6956 42932 6984
rect 42812 6390 42840 6956
rect 43180 6934 43208 9454
rect 43168 6928 43220 6934
rect 42890 6896 42946 6905
rect 43168 6870 43220 6876
rect 42890 6831 42892 6840
rect 42944 6831 42946 6840
rect 42892 6802 42944 6808
rect 42800 6384 42852 6390
rect 42800 6326 42852 6332
rect 42628 6038 42748 6066
rect 42628 5302 42656 6038
rect 42708 5908 42760 5914
rect 42708 5850 42760 5856
rect 42616 5296 42668 5302
rect 42616 5238 42668 5244
rect 42524 5092 42576 5098
rect 42524 5034 42576 5040
rect 42616 5092 42668 5098
rect 42616 5034 42668 5040
rect 42628 4978 42656 5034
rect 42536 4950 42656 4978
rect 42536 4282 42564 4950
rect 42614 4720 42670 4729
rect 42614 4655 42616 4664
rect 42668 4655 42670 4664
rect 42616 4626 42668 4632
rect 42524 4276 42576 4282
rect 42524 4218 42576 4224
rect 42616 4276 42668 4282
rect 42616 4218 42668 4224
rect 42524 4140 42576 4146
rect 42524 4082 42576 4088
rect 42432 4072 42484 4078
rect 42432 4014 42484 4020
rect 42352 3692 42472 3720
rect 42156 3664 42208 3670
rect 42156 3606 42208 3612
rect 42064 3596 42116 3602
rect 42064 3538 42116 3544
rect 42340 3596 42392 3602
rect 42340 3538 42392 3544
rect 42248 3528 42300 3534
rect 42248 3470 42300 3476
rect 42062 3360 42118 3369
rect 42062 3295 42118 3304
rect 41708 3182 41828 3210
rect 41880 3188 41932 3194
rect 41602 2544 41658 2553
rect 41602 2479 41658 2488
rect 41604 2304 41656 2310
rect 41604 2246 41656 2252
rect 41616 1970 41644 2246
rect 41604 1964 41656 1970
rect 41604 1906 41656 1912
rect 41708 1034 41736 3182
rect 41880 3130 41932 3136
rect 41788 2848 41840 2854
rect 41788 2790 41840 2796
rect 41616 1006 41736 1034
rect 41616 800 41644 1006
rect 41800 800 41828 2790
rect 41892 800 41920 3130
rect 41972 2984 42024 2990
rect 41972 2926 42024 2932
rect 41984 2825 42012 2926
rect 41970 2816 42026 2825
rect 41970 2751 42026 2760
rect 42076 800 42104 3295
rect 42260 800 42288 3470
rect 42352 2417 42380 3538
rect 42444 2922 42472 3692
rect 42432 2916 42484 2922
rect 42432 2858 42484 2864
rect 42430 2680 42486 2689
rect 42430 2615 42486 2624
rect 42444 2582 42472 2615
rect 42432 2576 42484 2582
rect 42432 2518 42484 2524
rect 42338 2408 42394 2417
rect 42338 2343 42394 2352
rect 42432 2372 42484 2378
rect 42432 2314 42484 2320
rect 42340 2304 42392 2310
rect 42340 2246 42392 2252
rect 42352 1902 42380 2246
rect 42340 1896 42392 1902
rect 42340 1838 42392 1844
rect 42444 1170 42472 2314
rect 42352 1142 42472 1170
rect 42352 800 42380 1142
rect 42536 800 42564 4082
rect 42628 800 42656 4218
rect 42720 3398 42748 5850
rect 42812 5778 42840 6326
rect 43076 6248 43128 6254
rect 43076 6190 43128 6196
rect 42984 6180 43036 6186
rect 42984 6122 43036 6128
rect 42800 5772 42852 5778
rect 42800 5714 42852 5720
rect 42800 5636 42852 5642
rect 42800 5578 42852 5584
rect 42812 3534 42840 5578
rect 42892 4684 42944 4690
rect 42892 4626 42944 4632
rect 42904 3738 42932 4626
rect 42892 3732 42944 3738
rect 42892 3674 42944 3680
rect 42800 3528 42852 3534
rect 42800 3470 42852 3476
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 42706 3088 42762 3097
rect 42706 3023 42762 3032
rect 42720 2514 42748 3023
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 42812 800 42840 3334
rect 42904 3233 42932 3674
rect 42890 3224 42946 3233
rect 42890 3159 42946 3168
rect 42892 3120 42944 3126
rect 42892 3062 42944 3068
rect 42904 800 42932 3062
rect 42996 2854 43024 6122
rect 43088 6089 43116 6190
rect 43074 6080 43130 6089
rect 43074 6015 43130 6024
rect 43076 4480 43128 4486
rect 43076 4422 43128 4428
rect 42984 2848 43036 2854
rect 42984 2790 43036 2796
rect 43088 800 43116 4422
rect 43180 2990 43208 6870
rect 43272 4049 43300 12038
rect 43536 10464 43588 10470
rect 43536 10406 43588 10412
rect 43352 9920 43404 9926
rect 43352 9862 43404 9868
rect 43364 7342 43392 9862
rect 43444 8832 43496 8838
rect 43444 8774 43496 8780
rect 43352 7336 43404 7342
rect 43352 7278 43404 7284
rect 43364 5409 43392 7278
rect 43456 6254 43484 8774
rect 43548 8566 43576 10406
rect 43640 9217 43668 27610
rect 43732 16574 43760 38490
rect 43824 31890 43852 58278
rect 44100 57798 44128 58482
rect 46848 58132 46900 58138
rect 46848 58074 46900 58080
rect 44088 57792 44140 57798
rect 44088 57734 44140 57740
rect 45284 57792 45336 57798
rect 45284 57734 45336 57740
rect 44220 57692 44516 57712
rect 44276 57690 44300 57692
rect 44356 57690 44380 57692
rect 44436 57690 44460 57692
rect 44298 57638 44300 57690
rect 44362 57638 44374 57690
rect 44436 57638 44438 57690
rect 44276 57636 44300 57638
rect 44356 57636 44380 57638
rect 44436 57636 44460 57638
rect 44220 57616 44516 57636
rect 45296 57594 45324 57734
rect 44916 57588 44968 57594
rect 44916 57530 44968 57536
rect 45284 57588 45336 57594
rect 45284 57530 45336 57536
rect 44220 56604 44516 56624
rect 44276 56602 44300 56604
rect 44356 56602 44380 56604
rect 44436 56602 44460 56604
rect 44298 56550 44300 56602
rect 44362 56550 44374 56602
rect 44436 56550 44438 56602
rect 44276 56548 44300 56550
rect 44356 56548 44380 56550
rect 44436 56548 44460 56550
rect 44220 56528 44516 56548
rect 44640 56296 44692 56302
rect 44640 56238 44692 56244
rect 44220 55516 44516 55536
rect 44276 55514 44300 55516
rect 44356 55514 44380 55516
rect 44436 55514 44460 55516
rect 44298 55462 44300 55514
rect 44362 55462 44374 55514
rect 44436 55462 44438 55514
rect 44276 55460 44300 55462
rect 44356 55460 44380 55462
rect 44436 55460 44460 55462
rect 44220 55440 44516 55460
rect 44220 54428 44516 54448
rect 44276 54426 44300 54428
rect 44356 54426 44380 54428
rect 44436 54426 44460 54428
rect 44298 54374 44300 54426
rect 44362 54374 44374 54426
rect 44436 54374 44438 54426
rect 44276 54372 44300 54374
rect 44356 54372 44380 54374
rect 44436 54372 44460 54374
rect 44220 54352 44516 54372
rect 44220 53340 44516 53360
rect 44276 53338 44300 53340
rect 44356 53338 44380 53340
rect 44436 53338 44460 53340
rect 44298 53286 44300 53338
rect 44362 53286 44374 53338
rect 44436 53286 44438 53338
rect 44276 53284 44300 53286
rect 44356 53284 44380 53286
rect 44436 53284 44460 53286
rect 44220 53264 44516 53284
rect 44220 52252 44516 52272
rect 44276 52250 44300 52252
rect 44356 52250 44380 52252
rect 44436 52250 44460 52252
rect 44298 52198 44300 52250
rect 44362 52198 44374 52250
rect 44436 52198 44438 52250
rect 44276 52196 44300 52198
rect 44356 52196 44380 52198
rect 44436 52196 44460 52198
rect 44220 52176 44516 52196
rect 44220 51164 44516 51184
rect 44276 51162 44300 51164
rect 44356 51162 44380 51164
rect 44436 51162 44460 51164
rect 44298 51110 44300 51162
rect 44362 51110 44374 51162
rect 44436 51110 44438 51162
rect 44276 51108 44300 51110
rect 44356 51108 44380 51110
rect 44436 51108 44460 51110
rect 44220 51088 44516 51108
rect 44220 50076 44516 50096
rect 44276 50074 44300 50076
rect 44356 50074 44380 50076
rect 44436 50074 44460 50076
rect 44298 50022 44300 50074
rect 44362 50022 44374 50074
rect 44436 50022 44438 50074
rect 44276 50020 44300 50022
rect 44356 50020 44380 50022
rect 44436 50020 44460 50022
rect 44220 50000 44516 50020
rect 44220 48988 44516 49008
rect 44276 48986 44300 48988
rect 44356 48986 44380 48988
rect 44436 48986 44460 48988
rect 44298 48934 44300 48986
rect 44362 48934 44374 48986
rect 44436 48934 44438 48986
rect 44276 48932 44300 48934
rect 44356 48932 44380 48934
rect 44436 48932 44460 48934
rect 44220 48912 44516 48932
rect 44220 47900 44516 47920
rect 44276 47898 44300 47900
rect 44356 47898 44380 47900
rect 44436 47898 44460 47900
rect 44298 47846 44300 47898
rect 44362 47846 44374 47898
rect 44436 47846 44438 47898
rect 44276 47844 44300 47846
rect 44356 47844 44380 47846
rect 44436 47844 44460 47846
rect 44220 47824 44516 47844
rect 44220 46812 44516 46832
rect 44276 46810 44300 46812
rect 44356 46810 44380 46812
rect 44436 46810 44460 46812
rect 44298 46758 44300 46810
rect 44362 46758 44374 46810
rect 44436 46758 44438 46810
rect 44276 46756 44300 46758
rect 44356 46756 44380 46758
rect 44436 46756 44460 46758
rect 44220 46736 44516 46756
rect 44220 45724 44516 45744
rect 44276 45722 44300 45724
rect 44356 45722 44380 45724
rect 44436 45722 44460 45724
rect 44298 45670 44300 45722
rect 44362 45670 44374 45722
rect 44436 45670 44438 45722
rect 44276 45668 44300 45670
rect 44356 45668 44380 45670
rect 44436 45668 44460 45670
rect 44220 45648 44516 45668
rect 44220 44636 44516 44656
rect 44276 44634 44300 44636
rect 44356 44634 44380 44636
rect 44436 44634 44460 44636
rect 44298 44582 44300 44634
rect 44362 44582 44374 44634
rect 44436 44582 44438 44634
rect 44276 44580 44300 44582
rect 44356 44580 44380 44582
rect 44436 44580 44460 44582
rect 44220 44560 44516 44580
rect 44220 43548 44516 43568
rect 44276 43546 44300 43548
rect 44356 43546 44380 43548
rect 44436 43546 44460 43548
rect 44298 43494 44300 43546
rect 44362 43494 44374 43546
rect 44436 43494 44438 43546
rect 44276 43492 44300 43494
rect 44356 43492 44380 43494
rect 44436 43492 44460 43494
rect 44220 43472 44516 43492
rect 44220 42460 44516 42480
rect 44276 42458 44300 42460
rect 44356 42458 44380 42460
rect 44436 42458 44460 42460
rect 44298 42406 44300 42458
rect 44362 42406 44374 42458
rect 44436 42406 44438 42458
rect 44276 42404 44300 42406
rect 44356 42404 44380 42406
rect 44436 42404 44460 42406
rect 44220 42384 44516 42404
rect 44220 41372 44516 41392
rect 44276 41370 44300 41372
rect 44356 41370 44380 41372
rect 44436 41370 44460 41372
rect 44298 41318 44300 41370
rect 44362 41318 44374 41370
rect 44436 41318 44438 41370
rect 44276 41316 44300 41318
rect 44356 41316 44380 41318
rect 44436 41316 44460 41318
rect 44220 41296 44516 41316
rect 44220 40284 44516 40304
rect 44276 40282 44300 40284
rect 44356 40282 44380 40284
rect 44436 40282 44460 40284
rect 44298 40230 44300 40282
rect 44362 40230 44374 40282
rect 44436 40230 44438 40282
rect 44276 40228 44300 40230
rect 44356 40228 44380 40230
rect 44436 40228 44460 40230
rect 44220 40208 44516 40228
rect 44220 39196 44516 39216
rect 44276 39194 44300 39196
rect 44356 39194 44380 39196
rect 44436 39194 44460 39196
rect 44298 39142 44300 39194
rect 44362 39142 44374 39194
rect 44436 39142 44438 39194
rect 44276 39140 44300 39142
rect 44356 39140 44380 39142
rect 44436 39140 44460 39142
rect 44220 39120 44516 39140
rect 44220 38108 44516 38128
rect 44276 38106 44300 38108
rect 44356 38106 44380 38108
rect 44436 38106 44460 38108
rect 44298 38054 44300 38106
rect 44362 38054 44374 38106
rect 44436 38054 44438 38106
rect 44276 38052 44300 38054
rect 44356 38052 44380 38054
rect 44436 38052 44460 38054
rect 44220 38032 44516 38052
rect 44220 37020 44516 37040
rect 44276 37018 44300 37020
rect 44356 37018 44380 37020
rect 44436 37018 44460 37020
rect 44298 36966 44300 37018
rect 44362 36966 44374 37018
rect 44436 36966 44438 37018
rect 44276 36964 44300 36966
rect 44356 36964 44380 36966
rect 44436 36964 44460 36966
rect 44220 36944 44516 36964
rect 44220 35932 44516 35952
rect 44276 35930 44300 35932
rect 44356 35930 44380 35932
rect 44436 35930 44460 35932
rect 44298 35878 44300 35930
rect 44362 35878 44374 35930
rect 44436 35878 44438 35930
rect 44276 35876 44300 35878
rect 44356 35876 44380 35878
rect 44436 35876 44460 35878
rect 44220 35856 44516 35876
rect 44088 35216 44140 35222
rect 44088 35158 44140 35164
rect 44100 34542 44128 35158
rect 44220 34844 44516 34864
rect 44276 34842 44300 34844
rect 44356 34842 44380 34844
rect 44436 34842 44460 34844
rect 44298 34790 44300 34842
rect 44362 34790 44374 34842
rect 44436 34790 44438 34842
rect 44276 34788 44300 34790
rect 44356 34788 44380 34790
rect 44436 34788 44460 34790
rect 44220 34768 44516 34788
rect 44088 34536 44140 34542
rect 44088 34478 44140 34484
rect 44220 33756 44516 33776
rect 44276 33754 44300 33756
rect 44356 33754 44380 33756
rect 44436 33754 44460 33756
rect 44298 33702 44300 33754
rect 44362 33702 44374 33754
rect 44436 33702 44438 33754
rect 44276 33700 44300 33702
rect 44356 33700 44380 33702
rect 44436 33700 44460 33702
rect 44220 33680 44516 33700
rect 44220 32668 44516 32688
rect 44276 32666 44300 32668
rect 44356 32666 44380 32668
rect 44436 32666 44460 32668
rect 44298 32614 44300 32666
rect 44362 32614 44374 32666
rect 44436 32614 44438 32666
rect 44276 32612 44300 32614
rect 44356 32612 44380 32614
rect 44436 32612 44460 32614
rect 44220 32592 44516 32612
rect 43812 31884 43864 31890
rect 43812 31826 43864 31832
rect 44220 31580 44516 31600
rect 44276 31578 44300 31580
rect 44356 31578 44380 31580
rect 44436 31578 44460 31580
rect 44298 31526 44300 31578
rect 44362 31526 44374 31578
rect 44436 31526 44438 31578
rect 44276 31524 44300 31526
rect 44356 31524 44380 31526
rect 44436 31524 44460 31526
rect 44220 31504 44516 31524
rect 44220 30492 44516 30512
rect 44276 30490 44300 30492
rect 44356 30490 44380 30492
rect 44436 30490 44460 30492
rect 44298 30438 44300 30490
rect 44362 30438 44374 30490
rect 44436 30438 44438 30490
rect 44276 30436 44300 30438
rect 44356 30436 44380 30438
rect 44436 30436 44460 30438
rect 44220 30416 44516 30436
rect 44220 29404 44516 29424
rect 44276 29402 44300 29404
rect 44356 29402 44380 29404
rect 44436 29402 44460 29404
rect 44298 29350 44300 29402
rect 44362 29350 44374 29402
rect 44436 29350 44438 29402
rect 44276 29348 44300 29350
rect 44356 29348 44380 29350
rect 44436 29348 44460 29350
rect 44220 29328 44516 29348
rect 44220 28316 44516 28336
rect 44276 28314 44300 28316
rect 44356 28314 44380 28316
rect 44436 28314 44460 28316
rect 44298 28262 44300 28314
rect 44362 28262 44374 28314
rect 44436 28262 44438 28314
rect 44276 28260 44300 28262
rect 44356 28260 44380 28262
rect 44436 28260 44460 28262
rect 44220 28240 44516 28260
rect 44220 27228 44516 27248
rect 44276 27226 44300 27228
rect 44356 27226 44380 27228
rect 44436 27226 44460 27228
rect 44298 27174 44300 27226
rect 44362 27174 44374 27226
rect 44436 27174 44438 27226
rect 44276 27172 44300 27174
rect 44356 27172 44380 27174
rect 44436 27172 44460 27174
rect 44220 27152 44516 27172
rect 44220 26140 44516 26160
rect 44276 26138 44300 26140
rect 44356 26138 44380 26140
rect 44436 26138 44460 26140
rect 44298 26086 44300 26138
rect 44362 26086 44374 26138
rect 44436 26086 44438 26138
rect 44276 26084 44300 26086
rect 44356 26084 44380 26086
rect 44436 26084 44460 26086
rect 44220 26064 44516 26084
rect 44220 25052 44516 25072
rect 44276 25050 44300 25052
rect 44356 25050 44380 25052
rect 44436 25050 44460 25052
rect 44298 24998 44300 25050
rect 44362 24998 44374 25050
rect 44436 24998 44438 25050
rect 44276 24996 44300 24998
rect 44356 24996 44380 24998
rect 44436 24996 44460 24998
rect 44220 24976 44516 24996
rect 44220 23964 44516 23984
rect 44276 23962 44300 23964
rect 44356 23962 44380 23964
rect 44436 23962 44460 23964
rect 44298 23910 44300 23962
rect 44362 23910 44374 23962
rect 44436 23910 44438 23962
rect 44276 23908 44300 23910
rect 44356 23908 44380 23910
rect 44436 23908 44460 23910
rect 44220 23888 44516 23908
rect 44220 22876 44516 22896
rect 44276 22874 44300 22876
rect 44356 22874 44380 22876
rect 44436 22874 44460 22876
rect 44298 22822 44300 22874
rect 44362 22822 44374 22874
rect 44436 22822 44438 22874
rect 44276 22820 44300 22822
rect 44356 22820 44380 22822
rect 44436 22820 44460 22822
rect 44220 22800 44516 22820
rect 44220 21788 44516 21808
rect 44276 21786 44300 21788
rect 44356 21786 44380 21788
rect 44436 21786 44460 21788
rect 44298 21734 44300 21786
rect 44362 21734 44374 21786
rect 44436 21734 44438 21786
rect 44276 21732 44300 21734
rect 44356 21732 44380 21734
rect 44436 21732 44460 21734
rect 44220 21712 44516 21732
rect 44220 20700 44516 20720
rect 44276 20698 44300 20700
rect 44356 20698 44380 20700
rect 44436 20698 44460 20700
rect 44298 20646 44300 20698
rect 44362 20646 44374 20698
rect 44436 20646 44438 20698
rect 44276 20644 44300 20646
rect 44356 20644 44380 20646
rect 44436 20644 44460 20646
rect 44220 20624 44516 20644
rect 44220 19612 44516 19632
rect 44276 19610 44300 19612
rect 44356 19610 44380 19612
rect 44436 19610 44460 19612
rect 44298 19558 44300 19610
rect 44362 19558 44374 19610
rect 44436 19558 44438 19610
rect 44276 19556 44300 19558
rect 44356 19556 44380 19558
rect 44436 19556 44460 19558
rect 44220 19536 44516 19556
rect 44220 18524 44516 18544
rect 44276 18522 44300 18524
rect 44356 18522 44380 18524
rect 44436 18522 44460 18524
rect 44298 18470 44300 18522
rect 44362 18470 44374 18522
rect 44436 18470 44438 18522
rect 44276 18468 44300 18470
rect 44356 18468 44380 18470
rect 44436 18468 44460 18470
rect 44220 18448 44516 18468
rect 44220 17436 44516 17456
rect 44276 17434 44300 17436
rect 44356 17434 44380 17436
rect 44436 17434 44460 17436
rect 44298 17382 44300 17434
rect 44362 17382 44374 17434
rect 44436 17382 44438 17434
rect 44276 17380 44300 17382
rect 44356 17380 44380 17382
rect 44436 17380 44460 17382
rect 44220 17360 44516 17380
rect 43732 16546 43944 16574
rect 43810 11384 43866 11393
rect 43810 11319 43866 11328
rect 43824 11082 43852 11319
rect 43812 11076 43864 11082
rect 43812 11018 43864 11024
rect 43626 9208 43682 9217
rect 43626 9143 43682 9152
rect 43824 8922 43852 11018
rect 43916 9586 43944 16546
rect 44220 16348 44516 16368
rect 44276 16346 44300 16348
rect 44356 16346 44380 16348
rect 44436 16346 44460 16348
rect 44298 16294 44300 16346
rect 44362 16294 44374 16346
rect 44436 16294 44438 16346
rect 44276 16292 44300 16294
rect 44356 16292 44380 16294
rect 44436 16292 44460 16294
rect 44220 16272 44516 16292
rect 44220 15260 44516 15280
rect 44276 15258 44300 15260
rect 44356 15258 44380 15260
rect 44436 15258 44460 15260
rect 44298 15206 44300 15258
rect 44362 15206 44374 15258
rect 44436 15206 44438 15258
rect 44276 15204 44300 15206
rect 44356 15204 44380 15206
rect 44436 15204 44460 15206
rect 44220 15184 44516 15204
rect 44220 14172 44516 14192
rect 44276 14170 44300 14172
rect 44356 14170 44380 14172
rect 44436 14170 44460 14172
rect 44298 14118 44300 14170
rect 44362 14118 44374 14170
rect 44436 14118 44438 14170
rect 44276 14116 44300 14118
rect 44356 14116 44380 14118
rect 44436 14116 44460 14118
rect 44220 14096 44516 14116
rect 44220 13084 44516 13104
rect 44276 13082 44300 13084
rect 44356 13082 44380 13084
rect 44436 13082 44460 13084
rect 44298 13030 44300 13082
rect 44362 13030 44374 13082
rect 44436 13030 44438 13082
rect 44276 13028 44300 13030
rect 44356 13028 44380 13030
rect 44436 13028 44460 13030
rect 44220 13008 44516 13028
rect 44220 11996 44516 12016
rect 44276 11994 44300 11996
rect 44356 11994 44380 11996
rect 44436 11994 44460 11996
rect 44298 11942 44300 11994
rect 44362 11942 44374 11994
rect 44436 11942 44438 11994
rect 44276 11940 44300 11942
rect 44356 11940 44380 11942
rect 44436 11940 44460 11942
rect 44220 11920 44516 11940
rect 44652 11558 44680 56238
rect 44824 54528 44876 54534
rect 44824 54470 44876 54476
rect 44836 54330 44864 54470
rect 44824 54324 44876 54330
rect 44824 54266 44876 54272
rect 44824 47048 44876 47054
rect 44824 46990 44876 46996
rect 44640 11552 44692 11558
rect 44640 11494 44692 11500
rect 44548 11076 44600 11082
rect 44548 11018 44600 11024
rect 44086 10976 44142 10985
rect 44086 10911 44142 10920
rect 43996 10668 44048 10674
rect 43996 10610 44048 10616
rect 43904 9580 43956 9586
rect 43904 9522 43956 9528
rect 44008 9489 44036 10610
rect 44100 10130 44128 10911
rect 44220 10908 44516 10928
rect 44276 10906 44300 10908
rect 44356 10906 44380 10908
rect 44436 10906 44460 10908
rect 44298 10854 44300 10906
rect 44362 10854 44374 10906
rect 44436 10854 44438 10906
rect 44276 10852 44300 10854
rect 44356 10852 44380 10854
rect 44436 10852 44460 10854
rect 44220 10832 44516 10852
rect 44180 10464 44232 10470
rect 44180 10406 44232 10412
rect 44088 10124 44140 10130
rect 44088 10066 44140 10072
rect 44192 9908 44220 10406
rect 44100 9880 44220 9908
rect 44100 9704 44128 9880
rect 44220 9820 44516 9840
rect 44276 9818 44300 9820
rect 44356 9818 44380 9820
rect 44436 9818 44460 9820
rect 44298 9766 44300 9818
rect 44362 9766 44374 9818
rect 44436 9766 44438 9818
rect 44276 9764 44300 9766
rect 44356 9764 44380 9766
rect 44436 9764 44460 9766
rect 44220 9744 44516 9764
rect 44560 9704 44588 11018
rect 44100 9676 44220 9704
rect 44088 9580 44140 9586
rect 44088 9522 44140 9528
rect 43994 9480 44050 9489
rect 43994 9415 44050 9424
rect 44100 9330 44128 9522
rect 43640 8894 43852 8922
rect 44008 9302 44128 9330
rect 43536 8560 43588 8566
rect 43536 8502 43588 8508
rect 43548 8430 43576 8502
rect 43536 8424 43588 8430
rect 43536 8366 43588 8372
rect 43640 8242 43668 8894
rect 43812 8832 43864 8838
rect 43812 8774 43864 8780
rect 43720 8560 43772 8566
rect 43720 8502 43772 8508
rect 43548 8214 43668 8242
rect 43444 6248 43496 6254
rect 43444 6190 43496 6196
rect 43350 5400 43406 5409
rect 43350 5335 43406 5344
rect 43352 5160 43404 5166
rect 43352 5102 43404 5108
rect 43364 4457 43392 5102
rect 43444 4548 43496 4554
rect 43444 4490 43496 4496
rect 43350 4448 43406 4457
rect 43350 4383 43406 4392
rect 43352 4072 43404 4078
rect 43258 4040 43314 4049
rect 43352 4014 43404 4020
rect 43258 3975 43314 3984
rect 43272 3602 43300 3975
rect 43260 3596 43312 3602
rect 43260 3538 43312 3544
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 43260 2848 43312 2854
rect 43166 2816 43222 2825
rect 43260 2790 43312 2796
rect 43166 2751 43222 2760
rect 43180 2582 43208 2751
rect 43168 2576 43220 2582
rect 43168 2518 43220 2524
rect 43272 1034 43300 2790
rect 43180 1006 43300 1034
rect 43180 800 43208 1006
rect 43364 800 43392 4014
rect 43456 800 43484 4490
rect 43548 2825 43576 8214
rect 43628 7880 43680 7886
rect 43628 7822 43680 7828
rect 43640 4729 43668 7822
rect 43626 4720 43682 4729
rect 43626 4655 43682 4664
rect 43628 4004 43680 4010
rect 43628 3946 43680 3952
rect 43534 2816 43590 2825
rect 43534 2751 43590 2760
rect 43536 2304 43588 2310
rect 43536 2246 43588 2252
rect 43548 1766 43576 2246
rect 43536 1760 43588 1766
rect 43536 1702 43588 1708
rect 43640 800 43668 3946
rect 43732 3942 43760 8502
rect 43824 6186 43852 8774
rect 44008 8566 44036 9302
rect 44192 8820 44220 9676
rect 44284 9676 44588 9704
rect 44284 8945 44312 9676
rect 44270 8936 44326 8945
rect 44270 8871 44326 8880
rect 44100 8792 44220 8820
rect 44548 8832 44600 8838
rect 43996 8560 44048 8566
rect 43996 8502 44048 8508
rect 43996 8288 44048 8294
rect 43996 8230 44048 8236
rect 43904 7948 43956 7954
rect 43904 7890 43956 7896
rect 43812 6180 43864 6186
rect 43812 6122 43864 6128
rect 43812 5840 43864 5846
rect 43812 5782 43864 5788
rect 43720 3936 43772 3942
rect 43720 3878 43772 3884
rect 43718 3768 43774 3777
rect 43718 3703 43774 3712
rect 43732 3602 43760 3703
rect 43720 3596 43772 3602
rect 43720 3538 43772 3544
rect 43718 3088 43774 3097
rect 43718 3023 43774 3032
rect 43732 2990 43760 3023
rect 43720 2984 43772 2990
rect 43720 2926 43772 2932
rect 43720 2304 43772 2310
rect 43720 2246 43772 2252
rect 43732 1698 43760 2246
rect 43720 1692 43772 1698
rect 43720 1634 43772 1640
rect 43824 800 43852 5782
rect 43916 4146 43944 7890
rect 44008 5778 44036 8230
rect 44100 7954 44128 8792
rect 44548 8774 44600 8780
rect 44220 8732 44516 8752
rect 44276 8730 44300 8732
rect 44356 8730 44380 8732
rect 44436 8730 44460 8732
rect 44298 8678 44300 8730
rect 44362 8678 44374 8730
rect 44436 8678 44438 8730
rect 44276 8676 44300 8678
rect 44356 8676 44380 8678
rect 44436 8676 44460 8678
rect 44220 8656 44516 8676
rect 44088 7948 44140 7954
rect 44088 7890 44140 7896
rect 44220 7644 44516 7664
rect 44276 7642 44300 7644
rect 44356 7642 44380 7644
rect 44436 7642 44460 7644
rect 44298 7590 44300 7642
rect 44362 7590 44374 7642
rect 44436 7590 44438 7642
rect 44276 7588 44300 7590
rect 44356 7588 44380 7590
rect 44436 7588 44460 7590
rect 44220 7568 44516 7588
rect 44088 7404 44140 7410
rect 44088 7346 44140 7352
rect 44100 5846 44128 7346
rect 44364 7268 44416 7274
rect 44364 7210 44416 7216
rect 44376 7002 44404 7210
rect 44364 6996 44416 7002
rect 44364 6938 44416 6944
rect 44560 6798 44588 8774
rect 44548 6792 44600 6798
rect 44548 6734 44600 6740
rect 44220 6556 44516 6576
rect 44276 6554 44300 6556
rect 44356 6554 44380 6556
rect 44436 6554 44460 6556
rect 44298 6502 44300 6554
rect 44362 6502 44374 6554
rect 44436 6502 44438 6554
rect 44276 6500 44300 6502
rect 44356 6500 44380 6502
rect 44436 6500 44460 6502
rect 44220 6480 44516 6500
rect 44180 6316 44232 6322
rect 44180 6258 44232 6264
rect 44088 5840 44140 5846
rect 44088 5782 44140 5788
rect 43996 5772 44048 5778
rect 43996 5714 44048 5720
rect 44192 5624 44220 6258
rect 44456 5908 44508 5914
rect 44456 5850 44508 5856
rect 44468 5642 44496 5850
rect 44008 5596 44220 5624
rect 44456 5636 44508 5642
rect 43904 4140 43956 4146
rect 43904 4082 43956 4088
rect 43904 3460 43956 3466
rect 43904 3402 43956 3408
rect 43916 800 43944 3402
rect 44008 1834 44036 5596
rect 44456 5578 44508 5584
rect 44548 5568 44600 5574
rect 44548 5510 44600 5516
rect 44220 5468 44516 5488
rect 44276 5466 44300 5468
rect 44356 5466 44380 5468
rect 44436 5466 44460 5468
rect 44298 5414 44300 5466
rect 44362 5414 44374 5466
rect 44436 5414 44438 5466
rect 44276 5412 44300 5414
rect 44356 5412 44380 5414
rect 44436 5412 44460 5414
rect 44220 5392 44516 5412
rect 44180 5296 44232 5302
rect 44180 5238 44232 5244
rect 44192 4593 44220 5238
rect 44560 5234 44588 5510
rect 44548 5228 44600 5234
rect 44548 5170 44600 5176
rect 44456 5160 44508 5166
rect 44508 5108 44588 5114
rect 44456 5102 44588 5108
rect 44468 5086 44588 5102
rect 44178 4584 44234 4593
rect 44178 4519 44234 4528
rect 44220 4380 44516 4400
rect 44276 4378 44300 4380
rect 44356 4378 44380 4380
rect 44436 4378 44460 4380
rect 44298 4326 44300 4378
rect 44362 4326 44374 4378
rect 44436 4326 44438 4378
rect 44276 4324 44300 4326
rect 44356 4324 44380 4326
rect 44436 4324 44460 4326
rect 44220 4304 44516 4324
rect 44560 3641 44588 5086
rect 44546 3632 44602 3641
rect 44546 3567 44602 3576
rect 44220 3292 44516 3312
rect 44276 3290 44300 3292
rect 44356 3290 44380 3292
rect 44436 3290 44460 3292
rect 44298 3238 44300 3290
rect 44362 3238 44374 3290
rect 44436 3238 44438 3290
rect 44276 3236 44300 3238
rect 44356 3236 44380 3238
rect 44436 3236 44460 3238
rect 44220 3216 44516 3236
rect 44088 3052 44140 3058
rect 44088 2994 44140 3000
rect 43996 1828 44048 1834
rect 43996 1770 44048 1776
rect 44100 800 44128 2994
rect 44652 2990 44680 11494
rect 44836 10538 44864 46990
rect 44824 10532 44876 10538
rect 44824 10474 44876 10480
rect 44928 10062 44956 57530
rect 45100 53032 45152 53038
rect 45100 52974 45152 52980
rect 45008 48000 45060 48006
rect 45008 47942 45060 47948
rect 45020 18766 45048 47942
rect 45008 18760 45060 18766
rect 45008 18702 45060 18708
rect 45112 11082 45140 52974
rect 46204 51400 46256 51406
rect 46204 51342 46256 51348
rect 46112 28144 46164 28150
rect 46112 28086 46164 28092
rect 46124 12434 46152 28086
rect 46216 14006 46244 51342
rect 46756 46980 46808 46986
rect 46756 46922 46808 46928
rect 46480 24880 46532 24886
rect 46480 24822 46532 24828
rect 46388 22568 46440 22574
rect 46388 22510 46440 22516
rect 46204 14000 46256 14006
rect 46204 13942 46256 13948
rect 46124 12406 46336 12434
rect 45652 11892 45704 11898
rect 45652 11834 45704 11840
rect 45560 11756 45612 11762
rect 45560 11698 45612 11704
rect 45572 11626 45600 11698
rect 45664 11626 45692 11834
rect 45560 11620 45612 11626
rect 45560 11562 45612 11568
rect 45652 11620 45704 11626
rect 45652 11562 45704 11568
rect 45374 11248 45430 11257
rect 45374 11183 45430 11192
rect 45100 11076 45152 11082
rect 45100 11018 45152 11024
rect 45008 10532 45060 10538
rect 45008 10474 45060 10480
rect 44916 10056 44968 10062
rect 44916 9998 44968 10004
rect 44916 9920 44968 9926
rect 44916 9862 44968 9868
rect 44824 9444 44876 9450
rect 44824 9386 44876 9392
rect 44732 9376 44784 9382
rect 44732 9318 44784 9324
rect 44744 7750 44772 9318
rect 44732 7744 44784 7750
rect 44732 7686 44784 7692
rect 44744 7342 44772 7686
rect 44732 7336 44784 7342
rect 44732 7278 44784 7284
rect 44732 6860 44784 6866
rect 44836 6848 44864 9386
rect 44928 7954 44956 9862
rect 44916 7948 44968 7954
rect 44916 7890 44968 7896
rect 44784 6820 44864 6848
rect 44732 6802 44784 6808
rect 44732 6248 44784 6254
rect 44732 6190 44784 6196
rect 44640 2984 44692 2990
rect 44640 2926 44692 2932
rect 44744 2836 44772 6190
rect 44824 3528 44876 3534
rect 44824 3470 44876 3476
rect 44546 2816 44602 2825
rect 44546 2751 44602 2760
rect 44652 2808 44772 2836
rect 44560 2582 44588 2751
rect 44548 2576 44600 2582
rect 44548 2518 44600 2524
rect 44220 2204 44516 2224
rect 44276 2202 44300 2204
rect 44356 2202 44380 2204
rect 44436 2202 44460 2204
rect 44298 2150 44300 2202
rect 44362 2150 44374 2202
rect 44436 2150 44438 2202
rect 44276 2148 44300 2150
rect 44356 2148 44380 2150
rect 44436 2148 44460 2150
rect 44220 2128 44516 2148
rect 44652 2088 44680 2808
rect 44836 2774 44864 3470
rect 44928 3126 44956 7890
rect 44916 3120 44968 3126
rect 44916 3062 44968 3068
rect 45020 2922 45048 10474
rect 45100 10464 45152 10470
rect 45100 10406 45152 10412
rect 45112 10198 45140 10406
rect 45100 10192 45152 10198
rect 45100 10134 45152 10140
rect 45112 8537 45140 10134
rect 45284 9988 45336 9994
rect 45284 9930 45336 9936
rect 45192 9376 45244 9382
rect 45192 9318 45244 9324
rect 45098 8528 45154 8537
rect 45098 8463 45154 8472
rect 45100 8424 45152 8430
rect 45100 8366 45152 8372
rect 45112 5302 45140 8366
rect 45204 6866 45232 9318
rect 45192 6860 45244 6866
rect 45192 6802 45244 6808
rect 45192 6724 45244 6730
rect 45192 6666 45244 6672
rect 45100 5296 45152 5302
rect 45100 5238 45152 5244
rect 45204 4146 45232 6666
rect 45192 4140 45244 4146
rect 45112 4100 45192 4128
rect 45112 3602 45140 4100
rect 45192 4082 45244 4088
rect 45296 4078 45324 9930
rect 45388 9518 45416 11183
rect 45468 11076 45520 11082
rect 45468 11018 45520 11024
rect 45376 9512 45428 9518
rect 45376 9454 45428 9460
rect 45376 8288 45428 8294
rect 45376 8230 45428 8236
rect 45388 5778 45416 8230
rect 45376 5772 45428 5778
rect 45376 5714 45428 5720
rect 45376 5636 45428 5642
rect 45376 5578 45428 5584
rect 45284 4072 45336 4078
rect 45284 4014 45336 4020
rect 45192 3732 45244 3738
rect 45192 3674 45244 3680
rect 45100 3596 45152 3602
rect 45100 3538 45152 3544
rect 45098 3496 45154 3505
rect 45098 3431 45154 3440
rect 45008 2916 45060 2922
rect 45008 2858 45060 2864
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44376 2060 44680 2088
rect 44744 2746 44864 2774
rect 44180 1896 44232 1902
rect 44180 1838 44232 1844
rect 44192 800 44220 1838
rect 44376 800 44404 2060
rect 44456 1420 44508 1426
rect 44456 1362 44508 1368
rect 44468 800 44496 1362
rect 44640 1216 44692 1222
rect 44640 1158 44692 1164
rect 44652 800 44680 1158
rect 44744 800 44772 2746
rect 44928 800 44956 2790
rect 45112 2774 45140 3431
rect 45020 2746 45140 2774
rect 45020 800 45048 2746
rect 45100 2304 45152 2310
rect 45100 2246 45152 2252
rect 45112 2038 45140 2246
rect 45100 2032 45152 2038
rect 45100 1974 45152 1980
rect 45204 800 45232 3674
rect 45284 3120 45336 3126
rect 45284 3062 45336 3068
rect 45296 800 45324 3062
rect 45388 1222 45416 5578
rect 45480 3670 45508 11018
rect 45572 7886 45600 11562
rect 46308 9926 46336 12406
rect 46296 9920 46348 9926
rect 46296 9862 46348 9868
rect 46020 9444 46072 9450
rect 46020 9386 46072 9392
rect 45836 9376 45888 9382
rect 45836 9318 45888 9324
rect 45652 8832 45704 8838
rect 45652 8774 45704 8780
rect 45560 7880 45612 7886
rect 45560 7822 45612 7828
rect 45560 7744 45612 7750
rect 45560 7686 45612 7692
rect 45572 6934 45600 7686
rect 45560 6928 45612 6934
rect 45560 6870 45612 6876
rect 45560 6792 45612 6798
rect 45560 6734 45612 6740
rect 45468 3664 45520 3670
rect 45468 3606 45520 3612
rect 45466 3360 45522 3369
rect 45466 3295 45522 3304
rect 45480 2922 45508 3295
rect 45468 2916 45520 2922
rect 45468 2858 45520 2864
rect 45572 2774 45600 6734
rect 45664 6458 45692 8774
rect 45744 8356 45796 8362
rect 45744 8298 45796 8304
rect 45652 6452 45704 6458
rect 45652 6394 45704 6400
rect 45664 6254 45692 6394
rect 45652 6248 45704 6254
rect 45652 6190 45704 6196
rect 45756 5386 45784 8298
rect 45848 6866 45876 9318
rect 45928 7200 45980 7206
rect 45928 7142 45980 7148
rect 45836 6860 45888 6866
rect 45836 6802 45888 6808
rect 45664 5358 45784 5386
rect 45664 5166 45692 5358
rect 45848 5250 45876 6802
rect 45756 5222 45876 5250
rect 45652 5160 45704 5166
rect 45652 5102 45704 5108
rect 45664 4486 45692 5102
rect 45652 4480 45704 4486
rect 45652 4422 45704 4428
rect 45652 4276 45704 4282
rect 45652 4218 45704 4224
rect 45664 3754 45692 4218
rect 45756 3942 45784 5222
rect 45836 5160 45888 5166
rect 45836 5102 45888 5108
rect 45848 4282 45876 5102
rect 45940 4690 45968 7142
rect 45928 4684 45980 4690
rect 45928 4626 45980 4632
rect 45836 4276 45888 4282
rect 45836 4218 45888 4224
rect 45836 4004 45888 4010
rect 45836 3946 45888 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45664 3726 45784 3754
rect 45652 3664 45704 3670
rect 45650 3632 45652 3641
rect 45704 3632 45706 3641
rect 45650 3567 45706 3576
rect 45756 3534 45784 3726
rect 45744 3528 45796 3534
rect 45744 3470 45796 3476
rect 45744 3392 45796 3398
rect 45744 3334 45796 3340
rect 45652 3188 45704 3194
rect 45652 3130 45704 3136
rect 45480 2746 45600 2774
rect 45376 1216 45428 1222
rect 45376 1158 45428 1164
rect 45480 800 45508 2746
rect 45664 800 45692 3130
rect 45756 800 45784 3334
rect 45848 1442 45876 3946
rect 45928 3936 45980 3942
rect 45928 3878 45980 3884
rect 45940 1578 45968 3878
rect 46032 2582 46060 9386
rect 46112 8832 46164 8838
rect 46112 8774 46164 8780
rect 46124 7274 46152 8774
rect 46204 8288 46256 8294
rect 46204 8230 46256 8236
rect 46216 8022 46244 8230
rect 46204 8016 46256 8022
rect 46204 7958 46256 7964
rect 46204 7744 46256 7750
rect 46204 7686 46256 7692
rect 46112 7268 46164 7274
rect 46112 7210 46164 7216
rect 46112 6724 46164 6730
rect 46112 6666 46164 6672
rect 46124 5914 46152 6666
rect 46112 5908 46164 5914
rect 46112 5850 46164 5856
rect 46216 5522 46244 7686
rect 46124 5494 46244 5522
rect 46124 4690 46152 5494
rect 46204 5364 46256 5370
rect 46204 5306 46256 5312
rect 46112 4684 46164 4690
rect 46112 4626 46164 4632
rect 46124 4554 46152 4626
rect 46216 4554 46244 5306
rect 46112 4548 46164 4554
rect 46112 4490 46164 4496
rect 46204 4548 46256 4554
rect 46204 4490 46256 4496
rect 46202 4448 46258 4457
rect 46202 4383 46258 4392
rect 46112 3052 46164 3058
rect 46112 2994 46164 3000
rect 46020 2576 46072 2582
rect 46020 2518 46072 2524
rect 45940 1550 46060 1578
rect 45848 1414 45968 1442
rect 45940 800 45968 1414
rect 46032 800 46060 1550
rect 46124 1068 46152 2994
rect 46216 1170 46244 4383
rect 46308 2582 46336 9862
rect 46400 9450 46428 22510
rect 46492 10470 46520 24822
rect 46480 10464 46532 10470
rect 46480 10406 46532 10412
rect 46388 9444 46440 9450
rect 46388 9386 46440 9392
rect 46388 8832 46440 8838
rect 46388 8774 46440 8780
rect 46400 7410 46428 8774
rect 46388 7404 46440 7410
rect 46388 7346 46440 7352
rect 46388 7200 46440 7206
rect 46388 7142 46440 7148
rect 46400 6662 46428 7142
rect 46388 6656 46440 6662
rect 46388 6598 46440 6604
rect 46388 5092 46440 5098
rect 46388 5034 46440 5040
rect 46400 4690 46428 5034
rect 46388 4684 46440 4690
rect 46388 4626 46440 4632
rect 46388 4480 46440 4486
rect 46388 4422 46440 4428
rect 46400 3738 46428 4422
rect 46388 3732 46440 3738
rect 46388 3674 46440 3680
rect 46388 3528 46440 3534
rect 46388 3470 46440 3476
rect 46400 2774 46428 3470
rect 46492 2990 46520 10406
rect 46768 9926 46796 46922
rect 46756 9920 46808 9926
rect 46756 9862 46808 9868
rect 46572 9376 46624 9382
rect 46572 9318 46624 9324
rect 46584 6798 46612 9318
rect 46664 8356 46716 8362
rect 46664 8298 46716 8304
rect 46572 6792 46624 6798
rect 46572 6734 46624 6740
rect 46572 6656 46624 6662
rect 46572 6598 46624 6604
rect 46584 4078 46612 6598
rect 46676 5817 46704 8298
rect 46662 5808 46718 5817
rect 46662 5743 46664 5752
rect 46716 5743 46718 5752
rect 46664 5714 46716 5720
rect 46768 5658 46796 9862
rect 46860 8974 46888 58074
rect 47032 41064 47084 41070
rect 47032 41006 47084 41012
rect 46938 12336 46994 12345
rect 46938 12271 46994 12280
rect 46848 8968 46900 8974
rect 46848 8910 46900 8916
rect 46860 7857 46888 8910
rect 46952 7954 46980 12271
rect 47044 10266 47072 41006
rect 47216 26852 47268 26858
rect 47216 26794 47268 26800
rect 47228 26314 47256 26794
rect 47216 26308 47268 26314
rect 47216 26250 47268 26256
rect 47412 13938 47440 59910
rect 48872 57996 48924 58002
rect 48872 57938 48924 57944
rect 47584 55684 47636 55690
rect 47584 55626 47636 55632
rect 47596 35894 47624 55626
rect 48780 54120 48832 54126
rect 48780 54062 48832 54068
rect 48228 52692 48280 52698
rect 48228 52634 48280 52640
rect 47504 35866 47624 35894
rect 47504 31890 47532 35866
rect 47492 31884 47544 31890
rect 47492 31826 47544 31832
rect 47504 26586 47532 31826
rect 48240 27606 48268 52634
rect 48688 46980 48740 46986
rect 48688 46922 48740 46928
rect 47584 27600 47636 27606
rect 47584 27542 47636 27548
rect 48228 27600 48280 27606
rect 48228 27542 48280 27548
rect 47492 26580 47544 26586
rect 47492 26522 47544 26528
rect 47596 26246 47624 27542
rect 48412 26444 48464 26450
rect 48412 26386 48464 26392
rect 47584 26240 47636 26246
rect 47584 26182 47636 26188
rect 47596 25702 47624 26182
rect 48424 25702 48452 26386
rect 48504 26376 48556 26382
rect 48504 26318 48556 26324
rect 47584 25696 47636 25702
rect 47584 25638 47636 25644
rect 48412 25696 48464 25702
rect 48412 25638 48464 25644
rect 47596 23662 47624 25638
rect 47584 23656 47636 23662
rect 47584 23598 47636 23604
rect 47596 15910 47624 23598
rect 47860 21344 47912 21350
rect 47860 21286 47912 21292
rect 47584 15904 47636 15910
rect 47584 15846 47636 15852
rect 47400 13932 47452 13938
rect 47400 13874 47452 13880
rect 47872 12434 47900 21286
rect 48424 18630 48452 25638
rect 48412 18624 48464 18630
rect 48412 18566 48464 18572
rect 48516 17610 48544 26318
rect 48504 17604 48556 17610
rect 48504 17546 48556 17552
rect 48596 14544 48648 14550
rect 48596 14486 48648 14492
rect 47780 12406 47900 12434
rect 47676 10464 47728 10470
rect 47676 10406 47728 10412
rect 47032 10260 47084 10266
rect 47032 10202 47084 10208
rect 47032 8832 47084 8838
rect 47032 8774 47084 8780
rect 47492 8832 47544 8838
rect 47492 8774 47544 8780
rect 46940 7948 46992 7954
rect 46940 7890 46992 7896
rect 46846 7848 46902 7857
rect 46846 7783 46902 7792
rect 46848 7744 46900 7750
rect 46848 7686 46900 7692
rect 46676 5630 46796 5658
rect 46572 4072 46624 4078
rect 46572 4014 46624 4020
rect 46570 3904 46626 3913
rect 46570 3839 46626 3848
rect 46584 3602 46612 3839
rect 46572 3596 46624 3602
rect 46572 3538 46624 3544
rect 46572 3460 46624 3466
rect 46572 3402 46624 3408
rect 46480 2984 46532 2990
rect 46480 2926 46532 2932
rect 46400 2746 46520 2774
rect 46296 2576 46348 2582
rect 46296 2518 46348 2524
rect 46216 1142 46336 1170
rect 46124 1040 46244 1068
rect 46216 800 46244 1040
rect 46308 800 46336 1142
rect 46492 800 46520 2746
rect 46584 800 46612 3402
rect 46676 2582 46704 5630
rect 46756 5160 46808 5166
rect 46860 5148 46888 7686
rect 47044 6254 47072 8774
rect 47124 8356 47176 8362
rect 47124 8298 47176 8304
rect 47136 6798 47164 8298
rect 47216 7744 47268 7750
rect 47216 7686 47268 7692
rect 47124 6792 47176 6798
rect 47124 6734 47176 6740
rect 47124 6656 47176 6662
rect 47124 6598 47176 6604
rect 47032 6248 47084 6254
rect 47032 6190 47084 6196
rect 46940 6112 46992 6118
rect 46940 6054 46992 6060
rect 46952 5846 46980 6054
rect 46940 5840 46992 5846
rect 46940 5782 46992 5788
rect 46808 5120 46888 5148
rect 46756 5102 46808 5108
rect 46768 4486 46796 5102
rect 46756 4480 46808 4486
rect 46756 4422 46808 4428
rect 46940 4276 46992 4282
rect 46940 4218 46992 4224
rect 46952 4162 46980 4218
rect 46768 4134 46980 4162
rect 46664 2576 46716 2582
rect 46664 2518 46716 2524
rect 46768 800 46796 4134
rect 47044 4060 47072 6190
rect 47136 4078 47164 6598
rect 47228 6390 47256 7686
rect 47400 7200 47452 7206
rect 47400 7142 47452 7148
rect 47308 6792 47360 6798
rect 47308 6734 47360 6740
rect 47216 6384 47268 6390
rect 47216 6326 47268 6332
rect 47320 5166 47348 6734
rect 47308 5160 47360 5166
rect 47308 5102 47360 5108
rect 46952 4032 47072 4060
rect 47124 4072 47176 4078
rect 46848 2372 46900 2378
rect 46848 2314 46900 2320
rect 46860 2106 46888 2314
rect 46848 2100 46900 2106
rect 46848 2042 46900 2048
rect 46848 1964 46900 1970
rect 46848 1906 46900 1912
rect 46860 800 46888 1906
rect 46952 1902 46980 4032
rect 47124 4014 47176 4020
rect 47136 3670 47164 4014
rect 47320 3942 47348 5102
rect 47412 4690 47440 7142
rect 47504 6866 47532 8774
rect 47584 7336 47636 7342
rect 47584 7278 47636 7284
rect 47492 6860 47544 6866
rect 47492 6802 47544 6808
rect 47400 4684 47452 4690
rect 47400 4626 47452 4632
rect 47308 3936 47360 3942
rect 47308 3878 47360 3884
rect 47216 3732 47268 3738
rect 47216 3674 47268 3680
rect 47124 3664 47176 3670
rect 47124 3606 47176 3612
rect 47032 2848 47084 2854
rect 47032 2790 47084 2796
rect 46940 1896 46992 1902
rect 46940 1838 46992 1844
rect 47044 800 47072 2790
rect 47228 1034 47256 3674
rect 47308 3528 47360 3534
rect 47308 3470 47360 3476
rect 47136 1006 47256 1034
rect 47136 800 47164 1006
rect 47320 800 47348 3470
rect 47412 3194 47440 4626
rect 47504 4010 47532 6802
rect 47596 4214 47624 7278
rect 47688 5914 47716 10406
rect 47780 9926 47808 12406
rect 47768 9920 47820 9926
rect 47768 9862 47820 9868
rect 47676 5908 47728 5914
rect 47676 5850 47728 5856
rect 47676 4480 47728 4486
rect 47676 4422 47728 4428
rect 47584 4208 47636 4214
rect 47584 4150 47636 4156
rect 47584 4072 47636 4078
rect 47584 4014 47636 4020
rect 47492 4004 47544 4010
rect 47492 3946 47544 3952
rect 47492 3460 47544 3466
rect 47492 3402 47544 3408
rect 47400 3188 47452 3194
rect 47400 3130 47452 3136
rect 47504 800 47532 3402
rect 47596 3233 47624 4014
rect 47688 3670 47716 4422
rect 47676 3664 47728 3670
rect 47676 3606 47728 3612
rect 47676 3460 47728 3466
rect 47676 3402 47728 3408
rect 47582 3224 47638 3233
rect 47582 3159 47638 3168
rect 47688 1748 47716 3402
rect 47780 3058 47808 9862
rect 48608 9450 48636 14486
rect 48700 14414 48728 46922
rect 48792 14482 48820 54062
rect 48780 14476 48832 14482
rect 48780 14418 48832 14424
rect 48688 14408 48740 14414
rect 48688 14350 48740 14356
rect 48884 12434 48912 57938
rect 48964 44260 49016 44266
rect 48964 44202 49016 44208
rect 48976 30598 49004 44202
rect 48964 30592 49016 30598
rect 48964 30534 49016 30540
rect 48976 30258 49004 30534
rect 48964 30252 49016 30258
rect 48964 30194 49016 30200
rect 48884 12406 49096 12434
rect 48688 12096 48740 12102
rect 48688 12038 48740 12044
rect 48596 9444 48648 9450
rect 48596 9386 48648 9392
rect 48412 9036 48464 9042
rect 48412 8978 48464 8984
rect 48424 8838 48452 8978
rect 48412 8832 48464 8838
rect 48412 8774 48464 8780
rect 48424 8634 48452 8774
rect 48412 8628 48464 8634
rect 48412 8570 48464 8576
rect 48136 8356 48188 8362
rect 48136 8298 48188 8304
rect 48504 8356 48556 8362
rect 48504 8298 48556 8304
rect 47860 7744 47912 7750
rect 47860 7686 47912 7692
rect 47872 6186 47900 7686
rect 48044 6724 48096 6730
rect 48044 6666 48096 6672
rect 47860 6180 47912 6186
rect 47860 6122 47912 6128
rect 47952 6180 48004 6186
rect 47952 6122 48004 6128
rect 47860 5908 47912 5914
rect 47860 5850 47912 5856
rect 47872 3913 47900 5850
rect 47964 5234 47992 6122
rect 47952 5228 48004 5234
rect 47952 5170 48004 5176
rect 48056 4690 48084 6666
rect 48148 5778 48176 8298
rect 48412 7880 48464 7886
rect 48412 7822 48464 7828
rect 48320 7744 48372 7750
rect 48320 7686 48372 7692
rect 48228 7200 48280 7206
rect 48228 7142 48280 7148
rect 48136 5772 48188 5778
rect 48136 5714 48188 5720
rect 48136 5024 48188 5030
rect 48136 4966 48188 4972
rect 48148 4690 48176 4966
rect 48044 4684 48096 4690
rect 47964 4644 48044 4672
rect 47858 3904 47914 3913
rect 47858 3839 47914 3848
rect 47768 3052 47820 3058
rect 47768 2994 47820 3000
rect 47766 2952 47822 2961
rect 47766 2887 47822 2896
rect 47860 2916 47912 2922
rect 47596 1720 47716 1748
rect 47596 800 47624 1720
rect 47780 800 47808 2887
rect 47860 2858 47912 2864
rect 47872 800 47900 2858
rect 47964 1970 47992 4644
rect 48044 4626 48096 4632
rect 48136 4684 48188 4690
rect 48136 4626 48188 4632
rect 48044 4140 48096 4146
rect 48044 4082 48096 4088
rect 47952 1964 48004 1970
rect 47952 1906 48004 1912
rect 48056 800 48084 4082
rect 48136 3664 48188 3670
rect 48136 3606 48188 3612
rect 48148 800 48176 3606
rect 48240 3602 48268 7142
rect 48332 5370 48360 7686
rect 48320 5364 48372 5370
rect 48320 5306 48372 5312
rect 48320 5228 48372 5234
rect 48320 5170 48372 5176
rect 48228 3596 48280 3602
rect 48228 3538 48280 3544
rect 48228 3052 48280 3058
rect 48228 2994 48280 3000
rect 48240 1426 48268 2994
rect 48332 2582 48360 5170
rect 48424 4214 48452 7822
rect 48516 5778 48544 8298
rect 48596 7812 48648 7818
rect 48596 7754 48648 7760
rect 48504 5772 48556 5778
rect 48504 5714 48556 5720
rect 48516 4457 48544 5714
rect 48608 5166 48636 7754
rect 48596 5160 48648 5166
rect 48596 5102 48648 5108
rect 48502 4448 48558 4457
rect 48502 4383 48558 4392
rect 48412 4208 48464 4214
rect 48412 4150 48464 4156
rect 48424 3505 48452 4150
rect 48608 4128 48636 5102
rect 48516 4100 48636 4128
rect 48516 3738 48544 4100
rect 48596 4004 48648 4010
rect 48596 3946 48648 3952
rect 48504 3732 48556 3738
rect 48504 3674 48556 3680
rect 48410 3496 48466 3505
rect 48410 3431 48466 3440
rect 48504 3052 48556 3058
rect 48504 2994 48556 3000
rect 48516 2650 48544 2994
rect 48504 2644 48556 2650
rect 48504 2586 48556 2592
rect 48320 2576 48372 2582
rect 48320 2518 48372 2524
rect 48502 2544 48558 2553
rect 48502 2479 48558 2488
rect 48228 1420 48280 1426
rect 48228 1362 48280 1368
rect 48516 1306 48544 2479
rect 48424 1278 48544 1306
rect 48320 1216 48372 1222
rect 48320 1158 48372 1164
rect 48332 800 48360 1158
rect 48424 800 48452 1278
rect 48608 800 48636 3946
rect 48700 3097 48728 12038
rect 48872 9444 48924 9450
rect 48872 9386 48924 9392
rect 48780 9376 48832 9382
rect 48780 9318 48832 9324
rect 48792 3126 48820 9318
rect 48780 3120 48832 3126
rect 48686 3088 48742 3097
rect 48780 3062 48832 3068
rect 48686 3023 48742 3032
rect 48688 2984 48740 2990
rect 48884 2972 48912 9386
rect 49068 8838 49096 12406
rect 49160 9382 49188 62766
rect 50080 62762 50108 63174
rect 50068 62756 50120 62762
rect 50068 62698 50120 62704
rect 49220 62588 49516 62608
rect 49276 62586 49300 62588
rect 49356 62586 49380 62588
rect 49436 62586 49460 62588
rect 49298 62534 49300 62586
rect 49362 62534 49374 62586
rect 49436 62534 49438 62586
rect 49276 62532 49300 62534
rect 49356 62532 49380 62534
rect 49436 62532 49460 62534
rect 49220 62512 49516 62532
rect 49608 62416 49660 62422
rect 49608 62358 49660 62364
rect 49220 61500 49516 61520
rect 49276 61498 49300 61500
rect 49356 61498 49380 61500
rect 49436 61498 49460 61500
rect 49298 61446 49300 61498
rect 49362 61446 49374 61498
rect 49436 61446 49438 61498
rect 49276 61444 49300 61446
rect 49356 61444 49380 61446
rect 49436 61444 49460 61446
rect 49220 61424 49516 61444
rect 49220 60412 49516 60432
rect 49276 60410 49300 60412
rect 49356 60410 49380 60412
rect 49436 60410 49460 60412
rect 49298 60358 49300 60410
rect 49362 60358 49374 60410
rect 49436 60358 49438 60410
rect 49276 60356 49300 60358
rect 49356 60356 49380 60358
rect 49436 60356 49460 60358
rect 49220 60336 49516 60356
rect 49620 60110 49648 62358
rect 49608 60104 49660 60110
rect 49608 60046 49660 60052
rect 49220 59324 49516 59344
rect 49276 59322 49300 59324
rect 49356 59322 49380 59324
rect 49436 59322 49460 59324
rect 49298 59270 49300 59322
rect 49362 59270 49374 59322
rect 49436 59270 49438 59322
rect 49276 59268 49300 59270
rect 49356 59268 49380 59270
rect 49436 59268 49460 59270
rect 49220 59248 49516 59268
rect 49220 58236 49516 58256
rect 49276 58234 49300 58236
rect 49356 58234 49380 58236
rect 49436 58234 49460 58236
rect 49298 58182 49300 58234
rect 49362 58182 49374 58234
rect 49436 58182 49438 58234
rect 49276 58180 49300 58182
rect 49356 58180 49380 58182
rect 49436 58180 49460 58182
rect 49220 58160 49516 58180
rect 49220 57148 49516 57168
rect 49276 57146 49300 57148
rect 49356 57146 49380 57148
rect 49436 57146 49460 57148
rect 49298 57094 49300 57146
rect 49362 57094 49374 57146
rect 49436 57094 49438 57146
rect 49276 57092 49300 57094
rect 49356 57092 49380 57094
rect 49436 57092 49460 57094
rect 49220 57072 49516 57092
rect 49220 56060 49516 56080
rect 49276 56058 49300 56060
rect 49356 56058 49380 56060
rect 49436 56058 49460 56060
rect 49298 56006 49300 56058
rect 49362 56006 49374 56058
rect 49436 56006 49438 56058
rect 49276 56004 49300 56006
rect 49356 56004 49380 56006
rect 49436 56004 49460 56006
rect 49220 55984 49516 56004
rect 49220 54972 49516 54992
rect 49276 54970 49300 54972
rect 49356 54970 49380 54972
rect 49436 54970 49460 54972
rect 49298 54918 49300 54970
rect 49362 54918 49374 54970
rect 49436 54918 49438 54970
rect 49276 54916 49300 54918
rect 49356 54916 49380 54918
rect 49436 54916 49460 54918
rect 49220 54896 49516 54916
rect 49220 53884 49516 53904
rect 49276 53882 49300 53884
rect 49356 53882 49380 53884
rect 49436 53882 49460 53884
rect 49298 53830 49300 53882
rect 49362 53830 49374 53882
rect 49436 53830 49438 53882
rect 49276 53828 49300 53830
rect 49356 53828 49380 53830
rect 49436 53828 49460 53830
rect 49220 53808 49516 53828
rect 49220 52796 49516 52816
rect 49276 52794 49300 52796
rect 49356 52794 49380 52796
rect 49436 52794 49460 52796
rect 49298 52742 49300 52794
rect 49362 52742 49374 52794
rect 49436 52742 49438 52794
rect 49276 52740 49300 52742
rect 49356 52740 49380 52742
rect 49436 52740 49460 52742
rect 49220 52720 49516 52740
rect 49220 51708 49516 51728
rect 49276 51706 49300 51708
rect 49356 51706 49380 51708
rect 49436 51706 49460 51708
rect 49298 51654 49300 51706
rect 49362 51654 49374 51706
rect 49436 51654 49438 51706
rect 49276 51652 49300 51654
rect 49356 51652 49380 51654
rect 49436 51652 49460 51654
rect 49220 51632 49516 51652
rect 49608 50720 49660 50726
rect 49608 50662 49660 50668
rect 49220 50620 49516 50640
rect 49276 50618 49300 50620
rect 49356 50618 49380 50620
rect 49436 50618 49460 50620
rect 49298 50566 49300 50618
rect 49362 50566 49374 50618
rect 49436 50566 49438 50618
rect 49276 50564 49300 50566
rect 49356 50564 49380 50566
rect 49436 50564 49460 50566
rect 49220 50544 49516 50564
rect 49220 49532 49516 49552
rect 49276 49530 49300 49532
rect 49356 49530 49380 49532
rect 49436 49530 49460 49532
rect 49298 49478 49300 49530
rect 49362 49478 49374 49530
rect 49436 49478 49438 49530
rect 49276 49476 49300 49478
rect 49356 49476 49380 49478
rect 49436 49476 49460 49478
rect 49220 49456 49516 49476
rect 49220 48444 49516 48464
rect 49276 48442 49300 48444
rect 49356 48442 49380 48444
rect 49436 48442 49460 48444
rect 49298 48390 49300 48442
rect 49362 48390 49374 48442
rect 49436 48390 49438 48442
rect 49276 48388 49300 48390
rect 49356 48388 49380 48390
rect 49436 48388 49460 48390
rect 49220 48368 49516 48388
rect 49220 47356 49516 47376
rect 49276 47354 49300 47356
rect 49356 47354 49380 47356
rect 49436 47354 49460 47356
rect 49298 47302 49300 47354
rect 49362 47302 49374 47354
rect 49436 47302 49438 47354
rect 49276 47300 49300 47302
rect 49356 47300 49380 47302
rect 49436 47300 49460 47302
rect 49220 47280 49516 47300
rect 49220 46268 49516 46288
rect 49276 46266 49300 46268
rect 49356 46266 49380 46268
rect 49436 46266 49460 46268
rect 49298 46214 49300 46266
rect 49362 46214 49374 46266
rect 49436 46214 49438 46266
rect 49276 46212 49300 46214
rect 49356 46212 49380 46214
rect 49436 46212 49460 46214
rect 49220 46192 49516 46212
rect 49220 45180 49516 45200
rect 49276 45178 49300 45180
rect 49356 45178 49380 45180
rect 49436 45178 49460 45180
rect 49298 45126 49300 45178
rect 49362 45126 49374 45178
rect 49436 45126 49438 45178
rect 49276 45124 49300 45126
rect 49356 45124 49380 45126
rect 49436 45124 49460 45126
rect 49220 45104 49516 45124
rect 49620 44742 49648 50662
rect 49608 44736 49660 44742
rect 49608 44678 49660 44684
rect 49620 44266 49648 44678
rect 49608 44260 49660 44266
rect 49608 44202 49660 44208
rect 49220 44092 49516 44112
rect 49276 44090 49300 44092
rect 49356 44090 49380 44092
rect 49436 44090 49460 44092
rect 49298 44038 49300 44090
rect 49362 44038 49374 44090
rect 49436 44038 49438 44090
rect 49276 44036 49300 44038
rect 49356 44036 49380 44038
rect 49436 44036 49460 44038
rect 49220 44016 49516 44036
rect 49220 43004 49516 43024
rect 49276 43002 49300 43004
rect 49356 43002 49380 43004
rect 49436 43002 49460 43004
rect 49298 42950 49300 43002
rect 49362 42950 49374 43002
rect 49436 42950 49438 43002
rect 49276 42948 49300 42950
rect 49356 42948 49380 42950
rect 49436 42948 49460 42950
rect 49220 42928 49516 42948
rect 49976 42356 50028 42362
rect 49976 42298 50028 42304
rect 49220 41916 49516 41936
rect 49276 41914 49300 41916
rect 49356 41914 49380 41916
rect 49436 41914 49460 41916
rect 49298 41862 49300 41914
rect 49362 41862 49374 41914
rect 49436 41862 49438 41914
rect 49276 41860 49300 41862
rect 49356 41860 49380 41862
rect 49436 41860 49460 41862
rect 49220 41840 49516 41860
rect 49220 40828 49516 40848
rect 49276 40826 49300 40828
rect 49356 40826 49380 40828
rect 49436 40826 49460 40828
rect 49298 40774 49300 40826
rect 49362 40774 49374 40826
rect 49436 40774 49438 40826
rect 49276 40772 49300 40774
rect 49356 40772 49380 40774
rect 49436 40772 49460 40774
rect 49220 40752 49516 40772
rect 49220 39740 49516 39760
rect 49276 39738 49300 39740
rect 49356 39738 49380 39740
rect 49436 39738 49460 39740
rect 49298 39686 49300 39738
rect 49362 39686 49374 39738
rect 49436 39686 49438 39738
rect 49276 39684 49300 39686
rect 49356 39684 49380 39686
rect 49436 39684 49460 39686
rect 49220 39664 49516 39684
rect 49220 38652 49516 38672
rect 49276 38650 49300 38652
rect 49356 38650 49380 38652
rect 49436 38650 49460 38652
rect 49298 38598 49300 38650
rect 49362 38598 49374 38650
rect 49436 38598 49438 38650
rect 49276 38596 49300 38598
rect 49356 38596 49380 38598
rect 49436 38596 49460 38598
rect 49220 38576 49516 38596
rect 49220 37564 49516 37584
rect 49276 37562 49300 37564
rect 49356 37562 49380 37564
rect 49436 37562 49460 37564
rect 49298 37510 49300 37562
rect 49362 37510 49374 37562
rect 49436 37510 49438 37562
rect 49276 37508 49300 37510
rect 49356 37508 49380 37510
rect 49436 37508 49460 37510
rect 49220 37488 49516 37508
rect 49220 36476 49516 36496
rect 49276 36474 49300 36476
rect 49356 36474 49380 36476
rect 49436 36474 49460 36476
rect 49298 36422 49300 36474
rect 49362 36422 49374 36474
rect 49436 36422 49438 36474
rect 49276 36420 49300 36422
rect 49356 36420 49380 36422
rect 49436 36420 49460 36422
rect 49220 36400 49516 36420
rect 49220 35388 49516 35408
rect 49276 35386 49300 35388
rect 49356 35386 49380 35388
rect 49436 35386 49460 35388
rect 49298 35334 49300 35386
rect 49362 35334 49374 35386
rect 49436 35334 49438 35386
rect 49276 35332 49300 35334
rect 49356 35332 49380 35334
rect 49436 35332 49460 35334
rect 49220 35312 49516 35332
rect 49220 34300 49516 34320
rect 49276 34298 49300 34300
rect 49356 34298 49380 34300
rect 49436 34298 49460 34300
rect 49298 34246 49300 34298
rect 49362 34246 49374 34298
rect 49436 34246 49438 34298
rect 49276 34244 49300 34246
rect 49356 34244 49380 34246
rect 49436 34244 49460 34246
rect 49220 34224 49516 34244
rect 49220 33212 49516 33232
rect 49276 33210 49300 33212
rect 49356 33210 49380 33212
rect 49436 33210 49460 33212
rect 49298 33158 49300 33210
rect 49362 33158 49374 33210
rect 49436 33158 49438 33210
rect 49276 33156 49300 33158
rect 49356 33156 49380 33158
rect 49436 33156 49460 33158
rect 49220 33136 49516 33156
rect 49884 32496 49936 32502
rect 49884 32438 49936 32444
rect 49220 32124 49516 32144
rect 49276 32122 49300 32124
rect 49356 32122 49380 32124
rect 49436 32122 49460 32124
rect 49298 32070 49300 32122
rect 49362 32070 49374 32122
rect 49436 32070 49438 32122
rect 49276 32068 49300 32070
rect 49356 32068 49380 32070
rect 49436 32068 49460 32070
rect 49220 32048 49516 32068
rect 49896 31822 49924 32438
rect 49884 31816 49936 31822
rect 49884 31758 49936 31764
rect 49220 31036 49516 31056
rect 49276 31034 49300 31036
rect 49356 31034 49380 31036
rect 49436 31034 49460 31036
rect 49298 30982 49300 31034
rect 49362 30982 49374 31034
rect 49436 30982 49438 31034
rect 49276 30980 49300 30982
rect 49356 30980 49380 30982
rect 49436 30980 49460 30982
rect 49220 30960 49516 30980
rect 49220 29948 49516 29968
rect 49276 29946 49300 29948
rect 49356 29946 49380 29948
rect 49436 29946 49460 29948
rect 49298 29894 49300 29946
rect 49362 29894 49374 29946
rect 49436 29894 49438 29946
rect 49276 29892 49300 29894
rect 49356 29892 49380 29894
rect 49436 29892 49460 29894
rect 49220 29872 49516 29892
rect 49220 28860 49516 28880
rect 49276 28858 49300 28860
rect 49356 28858 49380 28860
rect 49436 28858 49460 28860
rect 49298 28806 49300 28858
rect 49362 28806 49374 28858
rect 49436 28806 49438 28858
rect 49276 28804 49300 28806
rect 49356 28804 49380 28806
rect 49436 28804 49460 28806
rect 49220 28784 49516 28804
rect 49220 27772 49516 27792
rect 49276 27770 49300 27772
rect 49356 27770 49380 27772
rect 49436 27770 49460 27772
rect 49298 27718 49300 27770
rect 49362 27718 49374 27770
rect 49436 27718 49438 27770
rect 49276 27716 49300 27718
rect 49356 27716 49380 27718
rect 49436 27716 49460 27718
rect 49220 27696 49516 27716
rect 49220 26684 49516 26704
rect 49276 26682 49300 26684
rect 49356 26682 49380 26684
rect 49436 26682 49460 26684
rect 49298 26630 49300 26682
rect 49362 26630 49374 26682
rect 49436 26630 49438 26682
rect 49276 26628 49300 26630
rect 49356 26628 49380 26630
rect 49436 26628 49460 26630
rect 49220 26608 49516 26628
rect 49896 26586 49924 31758
rect 49884 26580 49936 26586
rect 49884 26522 49936 26528
rect 49332 26444 49384 26450
rect 49332 26386 49384 26392
rect 49608 26444 49660 26450
rect 49608 26386 49660 26392
rect 49344 26330 49372 26386
rect 49344 26314 49464 26330
rect 49344 26308 49476 26314
rect 49344 26302 49424 26308
rect 49424 26250 49476 26256
rect 49620 26246 49648 26386
rect 49896 26314 49924 26522
rect 49884 26308 49936 26314
rect 49884 26250 49936 26256
rect 49608 26240 49660 26246
rect 49608 26182 49660 26188
rect 49220 25596 49516 25616
rect 49276 25594 49300 25596
rect 49356 25594 49380 25596
rect 49436 25594 49460 25596
rect 49298 25542 49300 25594
rect 49362 25542 49374 25594
rect 49436 25542 49438 25594
rect 49276 25540 49300 25542
rect 49356 25540 49380 25542
rect 49436 25540 49460 25542
rect 49220 25520 49516 25540
rect 49220 24508 49516 24528
rect 49276 24506 49300 24508
rect 49356 24506 49380 24508
rect 49436 24506 49460 24508
rect 49298 24454 49300 24506
rect 49362 24454 49374 24506
rect 49436 24454 49438 24506
rect 49276 24452 49300 24454
rect 49356 24452 49380 24454
rect 49436 24452 49460 24454
rect 49220 24432 49516 24452
rect 49220 23420 49516 23440
rect 49276 23418 49300 23420
rect 49356 23418 49380 23420
rect 49436 23418 49460 23420
rect 49298 23366 49300 23418
rect 49362 23366 49374 23418
rect 49436 23366 49438 23418
rect 49276 23364 49300 23366
rect 49356 23364 49380 23366
rect 49436 23364 49460 23366
rect 49220 23344 49516 23364
rect 49220 22332 49516 22352
rect 49276 22330 49300 22332
rect 49356 22330 49380 22332
rect 49436 22330 49460 22332
rect 49298 22278 49300 22330
rect 49362 22278 49374 22330
rect 49436 22278 49438 22330
rect 49276 22276 49300 22278
rect 49356 22276 49380 22278
rect 49436 22276 49460 22278
rect 49220 22256 49516 22276
rect 49220 21244 49516 21264
rect 49276 21242 49300 21244
rect 49356 21242 49380 21244
rect 49436 21242 49460 21244
rect 49298 21190 49300 21242
rect 49362 21190 49374 21242
rect 49436 21190 49438 21242
rect 49276 21188 49300 21190
rect 49356 21188 49380 21190
rect 49436 21188 49460 21190
rect 49220 21168 49516 21188
rect 49220 20156 49516 20176
rect 49276 20154 49300 20156
rect 49356 20154 49380 20156
rect 49436 20154 49460 20156
rect 49298 20102 49300 20154
rect 49362 20102 49374 20154
rect 49436 20102 49438 20154
rect 49276 20100 49300 20102
rect 49356 20100 49380 20102
rect 49436 20100 49460 20102
rect 49220 20080 49516 20100
rect 49220 19068 49516 19088
rect 49276 19066 49300 19068
rect 49356 19066 49380 19068
rect 49436 19066 49460 19068
rect 49298 19014 49300 19066
rect 49362 19014 49374 19066
rect 49436 19014 49438 19066
rect 49276 19012 49300 19014
rect 49356 19012 49380 19014
rect 49436 19012 49460 19014
rect 49220 18992 49516 19012
rect 49220 17980 49516 18000
rect 49276 17978 49300 17980
rect 49356 17978 49380 17980
rect 49436 17978 49460 17980
rect 49298 17926 49300 17978
rect 49362 17926 49374 17978
rect 49436 17926 49438 17978
rect 49276 17924 49300 17926
rect 49356 17924 49380 17926
rect 49436 17924 49460 17926
rect 49220 17904 49516 17924
rect 49220 16892 49516 16912
rect 49276 16890 49300 16892
rect 49356 16890 49380 16892
rect 49436 16890 49460 16892
rect 49298 16838 49300 16890
rect 49362 16838 49374 16890
rect 49436 16838 49438 16890
rect 49276 16836 49300 16838
rect 49356 16836 49380 16838
rect 49436 16836 49460 16838
rect 49220 16816 49516 16836
rect 49220 15804 49516 15824
rect 49276 15802 49300 15804
rect 49356 15802 49380 15804
rect 49436 15802 49460 15804
rect 49298 15750 49300 15802
rect 49362 15750 49374 15802
rect 49436 15750 49438 15802
rect 49276 15748 49300 15750
rect 49356 15748 49380 15750
rect 49436 15748 49460 15750
rect 49220 15728 49516 15748
rect 49220 14716 49516 14736
rect 49276 14714 49300 14716
rect 49356 14714 49380 14716
rect 49436 14714 49460 14716
rect 49298 14662 49300 14714
rect 49362 14662 49374 14714
rect 49436 14662 49438 14714
rect 49276 14660 49300 14662
rect 49356 14660 49380 14662
rect 49436 14660 49460 14662
rect 49220 14640 49516 14660
rect 49220 13628 49516 13648
rect 49276 13626 49300 13628
rect 49356 13626 49380 13628
rect 49436 13626 49460 13628
rect 49298 13574 49300 13626
rect 49362 13574 49374 13626
rect 49436 13574 49438 13626
rect 49276 13572 49300 13574
rect 49356 13572 49380 13574
rect 49436 13572 49460 13574
rect 49220 13552 49516 13572
rect 49220 12540 49516 12560
rect 49276 12538 49300 12540
rect 49356 12538 49380 12540
rect 49436 12538 49460 12540
rect 49298 12486 49300 12538
rect 49362 12486 49374 12538
rect 49436 12486 49438 12538
rect 49276 12484 49300 12486
rect 49356 12484 49380 12486
rect 49436 12484 49460 12486
rect 49220 12464 49516 12484
rect 49220 11452 49516 11472
rect 49276 11450 49300 11452
rect 49356 11450 49380 11452
rect 49436 11450 49460 11452
rect 49298 11398 49300 11450
rect 49362 11398 49374 11450
rect 49436 11398 49438 11450
rect 49276 11396 49300 11398
rect 49356 11396 49380 11398
rect 49436 11396 49460 11398
rect 49220 11376 49516 11396
rect 49220 10364 49516 10384
rect 49276 10362 49300 10364
rect 49356 10362 49380 10364
rect 49436 10362 49460 10364
rect 49298 10310 49300 10362
rect 49362 10310 49374 10362
rect 49436 10310 49438 10362
rect 49276 10308 49300 10310
rect 49356 10308 49380 10310
rect 49436 10308 49460 10310
rect 49220 10288 49516 10308
rect 49148 9376 49200 9382
rect 49148 9318 49200 9324
rect 49608 9376 49660 9382
rect 49608 9318 49660 9324
rect 49220 9276 49516 9296
rect 49276 9274 49300 9276
rect 49356 9274 49380 9276
rect 49436 9274 49460 9276
rect 49298 9222 49300 9274
rect 49362 9222 49374 9274
rect 49436 9222 49438 9274
rect 49276 9220 49300 9222
rect 49356 9220 49380 9222
rect 49436 9220 49460 9222
rect 49220 9200 49516 9220
rect 49056 8832 49108 8838
rect 49056 8774 49108 8780
rect 49056 8356 49108 8362
rect 49056 8298 49108 8304
rect 48964 7200 49016 7206
rect 48964 7142 49016 7148
rect 48976 3602 49004 7142
rect 49068 5778 49096 8298
rect 49220 8188 49516 8208
rect 49276 8186 49300 8188
rect 49356 8186 49380 8188
rect 49436 8186 49460 8188
rect 49298 8134 49300 8186
rect 49362 8134 49374 8186
rect 49436 8134 49438 8186
rect 49276 8132 49300 8134
rect 49356 8132 49380 8134
rect 49436 8132 49460 8134
rect 49220 8112 49516 8132
rect 49148 7200 49200 7206
rect 49148 7142 49200 7148
rect 49056 5772 49108 5778
rect 49056 5714 49108 5720
rect 49068 4146 49096 5714
rect 49056 4140 49108 4146
rect 49056 4082 49108 4088
rect 49160 4026 49188 7142
rect 49220 7100 49516 7120
rect 49276 7098 49300 7100
rect 49356 7098 49380 7100
rect 49436 7098 49460 7100
rect 49298 7046 49300 7098
rect 49362 7046 49374 7098
rect 49436 7046 49438 7098
rect 49276 7044 49300 7046
rect 49356 7044 49380 7046
rect 49436 7044 49460 7046
rect 49220 7024 49516 7044
rect 49220 6012 49516 6032
rect 49276 6010 49300 6012
rect 49356 6010 49380 6012
rect 49436 6010 49460 6012
rect 49298 5958 49300 6010
rect 49362 5958 49374 6010
rect 49436 5958 49438 6010
rect 49276 5956 49300 5958
rect 49356 5956 49380 5958
rect 49436 5956 49460 5958
rect 49220 5936 49516 5956
rect 49220 4924 49516 4944
rect 49276 4922 49300 4924
rect 49356 4922 49380 4924
rect 49436 4922 49460 4924
rect 49298 4870 49300 4922
rect 49362 4870 49374 4922
rect 49436 4870 49438 4922
rect 49276 4868 49300 4870
rect 49356 4868 49380 4870
rect 49436 4868 49460 4870
rect 49220 4848 49516 4868
rect 49620 4706 49648 9318
rect 49988 8838 50016 42298
rect 50080 23186 50108 62698
rect 50436 59968 50488 59974
rect 50436 59910 50488 59916
rect 50252 57928 50304 57934
rect 50252 57870 50304 57876
rect 50264 57254 50292 57870
rect 50252 57248 50304 57254
rect 50252 57190 50304 57196
rect 50264 42702 50292 57190
rect 50448 50726 50476 59910
rect 50436 50720 50488 50726
rect 50436 50662 50488 50668
rect 50252 42696 50304 42702
rect 50252 42638 50304 42644
rect 50160 35624 50212 35630
rect 50160 35566 50212 35572
rect 50068 23180 50120 23186
rect 50068 23122 50120 23128
rect 50080 19990 50108 23122
rect 50068 19984 50120 19990
rect 50068 19926 50120 19932
rect 50172 12434 50200 35566
rect 50264 29646 50292 42638
rect 50712 29776 50764 29782
rect 50712 29718 50764 29724
rect 50252 29640 50304 29646
rect 50252 29582 50304 29588
rect 50264 26234 50292 29582
rect 50264 26206 50660 26234
rect 50344 19712 50396 19718
rect 50344 19654 50396 19660
rect 50172 12406 50292 12434
rect 50264 9382 50292 12406
rect 50252 9376 50304 9382
rect 50252 9318 50304 9324
rect 49700 8832 49752 8838
rect 49700 8774 49752 8780
rect 49976 8832 50028 8838
rect 49976 8774 50028 8780
rect 49240 4684 49292 4690
rect 49240 4626 49292 4632
rect 49528 4678 49648 4706
rect 49252 4214 49280 4626
rect 49240 4208 49292 4214
rect 49240 4150 49292 4156
rect 49240 4072 49292 4078
rect 49160 4020 49240 4026
rect 49160 4014 49292 4020
rect 49160 3998 49280 4014
rect 49056 3936 49108 3942
rect 49528 3924 49556 4678
rect 49056 3878 49108 3884
rect 49160 3896 49556 3924
rect 48964 3596 49016 3602
rect 48964 3538 49016 3544
rect 48688 2926 48740 2932
rect 48792 2944 48912 2972
rect 48700 2582 48728 2926
rect 48688 2576 48740 2582
rect 48792 2564 48820 2944
rect 48964 2848 49016 2854
rect 49068 2825 49096 3878
rect 49160 3720 49188 3896
rect 49220 3836 49516 3856
rect 49276 3834 49300 3836
rect 49356 3834 49380 3836
rect 49436 3834 49460 3836
rect 49298 3782 49300 3834
rect 49362 3782 49374 3834
rect 49436 3782 49438 3834
rect 49276 3780 49300 3782
rect 49356 3780 49380 3782
rect 49436 3780 49460 3782
rect 49220 3760 49516 3780
rect 49160 3692 49280 3720
rect 49148 3528 49200 3534
rect 49148 3470 49200 3476
rect 48964 2790 49016 2796
rect 49054 2816 49110 2825
rect 48872 2576 48924 2582
rect 48792 2536 48872 2564
rect 48688 2518 48740 2524
rect 48872 2518 48924 2524
rect 48870 2408 48926 2417
rect 48870 2343 48926 2352
rect 48688 1012 48740 1018
rect 48688 954 48740 960
rect 48700 800 48728 954
rect 48884 800 48912 2343
rect 48976 1018 49004 2790
rect 49054 2751 49110 2760
rect 49160 1442 49188 3470
rect 49252 2922 49280 3692
rect 49240 2916 49292 2922
rect 49240 2858 49292 2864
rect 49608 2916 49660 2922
rect 49608 2858 49660 2864
rect 49220 2748 49516 2768
rect 49276 2746 49300 2748
rect 49356 2746 49380 2748
rect 49436 2746 49460 2748
rect 49298 2694 49300 2746
rect 49362 2694 49374 2746
rect 49436 2694 49438 2746
rect 49276 2692 49300 2694
rect 49356 2692 49380 2694
rect 49436 2692 49460 2694
rect 49220 2672 49516 2692
rect 49240 2508 49292 2514
rect 49240 2450 49292 2456
rect 49068 1414 49188 1442
rect 48964 1012 49016 1018
rect 48964 954 49016 960
rect 49068 800 49096 1414
rect 49252 898 49280 2450
rect 49422 2272 49478 2281
rect 49422 2207 49478 2216
rect 49332 2100 49384 2106
rect 49332 2042 49384 2048
rect 49160 870 49280 898
rect 49160 800 49188 870
rect 49344 800 49372 2042
rect 49436 800 49464 2207
rect 49620 800 49648 2858
rect 49712 2582 49740 8774
rect 50160 7336 50212 7342
rect 50160 7278 50212 7284
rect 49976 7268 50028 7274
rect 49976 7210 50028 7216
rect 49884 7200 49936 7206
rect 49884 7142 49936 7148
rect 49792 6656 49844 6662
rect 49792 6598 49844 6604
rect 49804 4146 49832 6598
rect 49792 4140 49844 4146
rect 49792 4082 49844 4088
rect 49896 4078 49924 7142
rect 49988 6254 50016 7210
rect 50068 6656 50120 6662
rect 50068 6598 50120 6604
rect 49976 6248 50028 6254
rect 49976 6190 50028 6196
rect 49884 4072 49936 4078
rect 49882 4040 49884 4049
rect 49936 4040 49938 4049
rect 49882 3975 49938 3984
rect 49882 3904 49938 3913
rect 49882 3839 49938 3848
rect 49792 3120 49844 3126
rect 49792 3062 49844 3068
rect 49804 2650 49832 3062
rect 49792 2644 49844 2650
rect 49792 2586 49844 2592
rect 49700 2576 49752 2582
rect 49700 2518 49752 2524
rect 49790 2544 49846 2553
rect 49790 2479 49846 2488
rect 49804 2446 49832 2479
rect 49792 2440 49844 2446
rect 49792 2382 49844 2388
rect 49700 1420 49752 1426
rect 49700 1362 49752 1368
rect 49712 800 49740 1362
rect 49896 800 49924 3839
rect 49988 2961 50016 6190
rect 50080 3602 50108 6598
rect 50172 5778 50200 7278
rect 50160 5772 50212 5778
rect 50160 5714 50212 5720
rect 50172 3942 50200 5714
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 50160 3732 50212 3738
rect 50160 3674 50212 3680
rect 50068 3596 50120 3602
rect 50068 3538 50120 3544
rect 50068 3392 50120 3398
rect 50068 3334 50120 3340
rect 49974 2952 50030 2961
rect 49974 2887 50030 2896
rect 49976 2848 50028 2854
rect 49976 2790 50028 2796
rect 49988 800 50016 2790
rect 50080 2582 50108 3334
rect 50068 2576 50120 2582
rect 50068 2518 50120 2524
rect 50172 1426 50200 3674
rect 50264 2990 50292 9318
rect 50356 9042 50384 19654
rect 50528 18964 50580 18970
rect 50528 18906 50580 18912
rect 50344 9036 50396 9042
rect 50344 8978 50396 8984
rect 50436 8832 50488 8838
rect 50436 8774 50488 8780
rect 50344 7744 50396 7750
rect 50344 7686 50396 7692
rect 50356 5166 50384 7686
rect 50344 5160 50396 5166
rect 50344 5102 50396 5108
rect 50344 4684 50396 4690
rect 50344 4626 50396 4632
rect 50356 4282 50384 4626
rect 50344 4276 50396 4282
rect 50344 4218 50396 4224
rect 50344 3460 50396 3466
rect 50344 3402 50396 3408
rect 50252 2984 50304 2990
rect 50252 2926 50304 2932
rect 50356 2774 50384 3402
rect 50264 2746 50384 2774
rect 50160 1420 50212 1426
rect 50160 1362 50212 1368
rect 50160 1284 50212 1290
rect 50160 1226 50212 1232
rect 50172 800 50200 1226
rect 50264 800 50292 2746
rect 50448 2582 50476 8774
rect 50540 5302 50568 18906
rect 50632 15910 50660 26206
rect 50724 16726 50752 29718
rect 50816 18834 50844 66982
rect 54220 66396 54516 66416
rect 54276 66394 54300 66396
rect 54356 66394 54380 66396
rect 54436 66394 54460 66396
rect 54298 66342 54300 66394
rect 54362 66342 54374 66394
rect 54436 66342 54438 66394
rect 54276 66340 54300 66342
rect 54356 66340 54380 66342
rect 54436 66340 54460 66342
rect 54220 66320 54516 66340
rect 54220 65308 54516 65328
rect 54276 65306 54300 65308
rect 54356 65306 54380 65308
rect 54436 65306 54460 65308
rect 54298 65254 54300 65306
rect 54362 65254 54374 65306
rect 54436 65254 54438 65306
rect 54276 65252 54300 65254
rect 54356 65252 54380 65254
rect 54436 65252 54460 65254
rect 54220 65232 54516 65252
rect 54220 64220 54516 64240
rect 54276 64218 54300 64220
rect 54356 64218 54380 64220
rect 54436 64218 54460 64220
rect 54298 64166 54300 64218
rect 54362 64166 54374 64218
rect 54436 64166 54438 64218
rect 54276 64164 54300 64166
rect 54356 64164 54380 64166
rect 54436 64164 54460 64166
rect 54220 64144 54516 64164
rect 54220 63132 54516 63152
rect 54276 63130 54300 63132
rect 54356 63130 54380 63132
rect 54436 63130 54460 63132
rect 54298 63078 54300 63130
rect 54362 63078 54374 63130
rect 54436 63078 54438 63130
rect 54276 63076 54300 63078
rect 54356 63076 54380 63078
rect 54436 63076 54460 63078
rect 54220 63056 54516 63076
rect 51448 62688 51500 62694
rect 51448 62630 51500 62636
rect 51460 60722 51488 62630
rect 54220 62044 54516 62064
rect 54276 62042 54300 62044
rect 54356 62042 54380 62044
rect 54436 62042 54460 62044
rect 54298 61990 54300 62042
rect 54362 61990 54374 62042
rect 54436 61990 54438 62042
rect 54276 61988 54300 61990
rect 54356 61988 54380 61990
rect 54436 61988 54460 61990
rect 54220 61968 54516 61988
rect 54220 60956 54516 60976
rect 54276 60954 54300 60956
rect 54356 60954 54380 60956
rect 54436 60954 54460 60956
rect 54298 60902 54300 60954
rect 54362 60902 54374 60954
rect 54436 60902 54438 60954
rect 54276 60900 54300 60902
rect 54356 60900 54380 60902
rect 54436 60900 54460 60902
rect 54220 60880 54516 60900
rect 51448 60716 51500 60722
rect 51448 60658 51500 60664
rect 51460 60246 51488 60658
rect 51448 60240 51500 60246
rect 51448 60182 51500 60188
rect 50988 60172 51040 60178
rect 50988 60114 51040 60120
rect 52368 60172 52420 60178
rect 52368 60114 52420 60120
rect 51000 59974 51028 60114
rect 51632 60104 51684 60110
rect 51632 60046 51684 60052
rect 50988 59968 51040 59974
rect 50988 59910 51040 59916
rect 51644 59430 51672 60046
rect 52092 59968 52144 59974
rect 52092 59910 52144 59916
rect 51632 59424 51684 59430
rect 51632 59366 51684 59372
rect 51448 57520 51500 57526
rect 51448 57462 51500 57468
rect 51356 42152 51408 42158
rect 51356 42094 51408 42100
rect 50896 40724 50948 40730
rect 50896 40666 50948 40672
rect 50804 18828 50856 18834
rect 50804 18770 50856 18776
rect 50712 16720 50764 16726
rect 50712 16662 50764 16668
rect 50620 15904 50672 15910
rect 50620 15846 50672 15852
rect 50632 8634 50660 15846
rect 50724 8634 50752 16662
rect 50908 9110 50936 40666
rect 51264 36032 51316 36038
rect 51264 35974 51316 35980
rect 51276 11150 51304 35974
rect 51264 11144 51316 11150
rect 51264 11086 51316 11092
rect 51368 10742 51396 42094
rect 51356 10736 51408 10742
rect 51356 10678 51408 10684
rect 50896 9104 50948 9110
rect 50896 9046 50948 9052
rect 51356 9104 51408 9110
rect 51356 9046 51408 9052
rect 50620 8628 50672 8634
rect 50620 8570 50672 8576
rect 50712 8628 50764 8634
rect 50712 8570 50764 8576
rect 50528 5296 50580 5302
rect 50528 5238 50580 5244
rect 50632 5166 50660 8570
rect 50896 7744 50948 7750
rect 50896 7686 50948 7692
rect 50804 7200 50856 7206
rect 50804 7142 50856 7148
rect 50712 6656 50764 6662
rect 50712 6598 50764 6604
rect 50528 5160 50580 5166
rect 50528 5102 50580 5108
rect 50620 5160 50672 5166
rect 50620 5102 50672 5108
rect 50540 3398 50568 5102
rect 50620 4140 50672 4146
rect 50620 4082 50672 4088
rect 50528 3392 50580 3398
rect 50528 3334 50580 3340
rect 50528 3120 50580 3126
rect 50528 3062 50580 3068
rect 50436 2576 50488 2582
rect 50436 2518 50488 2524
rect 50540 1170 50568 3062
rect 50448 1142 50568 1170
rect 50448 800 50476 1142
rect 50632 1034 50660 4082
rect 50724 4078 50752 6598
rect 50816 4690 50844 7142
rect 50908 6254 50936 7686
rect 51264 6656 51316 6662
rect 51264 6598 51316 6604
rect 50896 6248 50948 6254
rect 50896 6190 50948 6196
rect 50804 4684 50856 4690
rect 50804 4626 50856 4632
rect 50712 4072 50764 4078
rect 50712 4014 50764 4020
rect 50804 4072 50856 4078
rect 50804 4014 50856 4020
rect 50724 3913 50752 4014
rect 50710 3904 50766 3913
rect 50710 3839 50766 3848
rect 50816 3482 50844 4014
rect 50540 1006 50660 1034
rect 50724 3454 50844 3482
rect 50540 800 50568 1006
rect 50724 800 50752 3454
rect 50804 3392 50856 3398
rect 50804 3334 50856 3340
rect 50816 1290 50844 3334
rect 50908 3233 50936 6190
rect 51172 5772 51224 5778
rect 51172 5714 51224 5720
rect 51080 5228 51132 5234
rect 51080 5170 51132 5176
rect 51092 4128 51120 5170
rect 51184 4146 51212 5714
rect 51000 4100 51120 4128
rect 51172 4140 51224 4146
rect 50894 3224 50950 3233
rect 50894 3159 50950 3168
rect 50896 3052 50948 3058
rect 50896 2994 50948 3000
rect 50804 1284 50856 1290
rect 50804 1226 50856 1232
rect 50908 800 50936 2994
rect 51000 800 51028 4100
rect 51172 4082 51224 4088
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 51092 3398 51120 3878
rect 51276 3602 51304 6598
rect 51368 5098 51396 9046
rect 51460 8838 51488 57462
rect 51644 55894 51672 59366
rect 51632 55888 51684 55894
rect 51632 55830 51684 55836
rect 52000 53032 52052 53038
rect 52000 52974 52052 52980
rect 51816 14272 51868 14278
rect 51816 14214 51868 14220
rect 51448 8832 51500 8838
rect 51448 8774 51500 8780
rect 51632 8832 51684 8838
rect 51632 8774 51684 8780
rect 51448 8628 51500 8634
rect 51500 8588 51580 8616
rect 51448 8570 51500 8576
rect 51448 7744 51500 7750
rect 51448 7686 51500 7692
rect 51356 5092 51408 5098
rect 51356 5034 51408 5040
rect 51460 4690 51488 7686
rect 51552 5030 51580 8588
rect 51540 5024 51592 5030
rect 51540 4966 51592 4972
rect 51448 4684 51500 4690
rect 51448 4626 51500 4632
rect 51460 3738 51488 4626
rect 51540 4004 51592 4010
rect 51540 3946 51592 3952
rect 51448 3732 51500 3738
rect 51448 3674 51500 3680
rect 51264 3596 51316 3602
rect 51264 3538 51316 3544
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 51080 3392 51132 3398
rect 51080 3334 51132 3340
rect 51172 3392 51224 3398
rect 51172 3334 51224 3340
rect 51078 3224 51134 3233
rect 51078 3159 51134 3168
rect 51092 2106 51120 3159
rect 51080 2100 51132 2106
rect 51080 2042 51132 2048
rect 51184 800 51212 3334
rect 51368 2990 51396 3470
rect 51448 3460 51500 3466
rect 51448 3402 51500 3408
rect 51356 2984 51408 2990
rect 51356 2926 51408 2932
rect 51264 2848 51316 2854
rect 51264 2790 51316 2796
rect 51276 800 51304 2790
rect 51460 800 51488 3402
rect 51552 800 51580 3946
rect 51644 2582 51672 8774
rect 51828 8634 51856 14214
rect 51908 13320 51960 13326
rect 51908 13262 51960 13268
rect 51920 8634 51948 13262
rect 52012 8838 52040 52974
rect 52104 41682 52132 59910
rect 52380 59430 52408 60114
rect 53196 59968 53248 59974
rect 53196 59910 53248 59916
rect 52368 59424 52420 59430
rect 52368 59366 52420 59372
rect 53012 53032 53064 53038
rect 53012 52974 53064 52980
rect 53024 52902 53052 52974
rect 53012 52896 53064 52902
rect 53012 52838 53064 52844
rect 52092 41676 52144 41682
rect 52092 41618 52144 41624
rect 53024 29578 53052 52838
rect 53012 29572 53064 29578
rect 53012 29514 53064 29520
rect 52552 20868 52604 20874
rect 52552 20810 52604 20816
rect 52564 12434 52592 20810
rect 52472 12406 52592 12434
rect 52472 8838 52500 12406
rect 53012 11824 53064 11830
rect 53012 11766 53064 11772
rect 53024 8838 53052 11766
rect 53208 11762 53236 59910
rect 54220 59868 54516 59888
rect 54276 59866 54300 59868
rect 54356 59866 54380 59868
rect 54436 59866 54460 59868
rect 54298 59814 54300 59866
rect 54362 59814 54374 59866
rect 54436 59814 54438 59866
rect 54276 59812 54300 59814
rect 54356 59812 54380 59814
rect 54436 59812 54460 59814
rect 54220 59792 54516 59812
rect 54220 58780 54516 58800
rect 54276 58778 54300 58780
rect 54356 58778 54380 58780
rect 54436 58778 54460 58780
rect 54298 58726 54300 58778
rect 54362 58726 54374 58778
rect 54436 58726 54438 58778
rect 54276 58724 54300 58726
rect 54356 58724 54380 58726
rect 54436 58724 54460 58726
rect 54220 58704 54516 58724
rect 54220 57692 54516 57712
rect 54276 57690 54300 57692
rect 54356 57690 54380 57692
rect 54436 57690 54460 57692
rect 54298 57638 54300 57690
rect 54362 57638 54374 57690
rect 54436 57638 54438 57690
rect 54276 57636 54300 57638
rect 54356 57636 54380 57638
rect 54436 57636 54460 57638
rect 54220 57616 54516 57636
rect 54220 56604 54516 56624
rect 54276 56602 54300 56604
rect 54356 56602 54380 56604
rect 54436 56602 54460 56604
rect 54298 56550 54300 56602
rect 54362 56550 54374 56602
rect 54436 56550 54438 56602
rect 54276 56548 54300 56550
rect 54356 56548 54380 56550
rect 54436 56548 54460 56550
rect 54220 56528 54516 56548
rect 54220 55516 54516 55536
rect 54276 55514 54300 55516
rect 54356 55514 54380 55516
rect 54436 55514 54460 55516
rect 54298 55462 54300 55514
rect 54362 55462 54374 55514
rect 54436 55462 54438 55514
rect 54276 55460 54300 55462
rect 54356 55460 54380 55462
rect 54436 55460 54460 55462
rect 54220 55440 54516 55460
rect 54220 54428 54516 54448
rect 54276 54426 54300 54428
rect 54356 54426 54380 54428
rect 54436 54426 54460 54428
rect 54298 54374 54300 54426
rect 54362 54374 54374 54426
rect 54436 54374 54438 54426
rect 54276 54372 54300 54374
rect 54356 54372 54380 54374
rect 54436 54372 54460 54374
rect 54220 54352 54516 54372
rect 53932 53440 53984 53446
rect 53932 53382 53984 53388
rect 53944 53174 53972 53382
rect 54220 53340 54516 53360
rect 54276 53338 54300 53340
rect 54356 53338 54380 53340
rect 54436 53338 54460 53340
rect 54298 53286 54300 53338
rect 54362 53286 54374 53338
rect 54436 53286 54438 53338
rect 54276 53284 54300 53286
rect 54356 53284 54380 53286
rect 54436 53284 54460 53286
rect 54220 53264 54516 53284
rect 53932 53168 53984 53174
rect 53932 53110 53984 53116
rect 53840 52896 53892 52902
rect 53840 52838 53892 52844
rect 53852 52562 53880 52838
rect 53840 52556 53892 52562
rect 53840 52498 53892 52504
rect 53944 51814 53972 53110
rect 54576 53032 54628 53038
rect 54576 52974 54628 52980
rect 54668 53032 54720 53038
rect 54668 52974 54720 52980
rect 54588 52494 54616 52974
rect 54680 52562 54708 52974
rect 54668 52556 54720 52562
rect 54668 52498 54720 52504
rect 54024 52488 54076 52494
rect 54024 52430 54076 52436
rect 54576 52488 54628 52494
rect 54576 52430 54628 52436
rect 53932 51808 53984 51814
rect 53932 51750 53984 51756
rect 54036 50386 54064 52430
rect 54220 52252 54516 52272
rect 54276 52250 54300 52252
rect 54356 52250 54380 52252
rect 54436 52250 54460 52252
rect 54298 52198 54300 52250
rect 54362 52198 54374 52250
rect 54436 52198 54438 52250
rect 54276 52196 54300 52198
rect 54356 52196 54380 52198
rect 54436 52196 54460 52198
rect 54220 52176 54516 52196
rect 54220 51164 54516 51184
rect 54276 51162 54300 51164
rect 54356 51162 54380 51164
rect 54436 51162 54460 51164
rect 54298 51110 54300 51162
rect 54362 51110 54374 51162
rect 54436 51110 54438 51162
rect 54276 51108 54300 51110
rect 54356 51108 54380 51110
rect 54436 51108 54460 51110
rect 54220 51088 54516 51108
rect 54024 50380 54076 50386
rect 54024 50322 54076 50328
rect 54220 50076 54516 50096
rect 54276 50074 54300 50076
rect 54356 50074 54380 50076
rect 54436 50074 54460 50076
rect 54298 50022 54300 50074
rect 54362 50022 54374 50074
rect 54436 50022 54438 50074
rect 54276 50020 54300 50022
rect 54356 50020 54380 50022
rect 54436 50020 54460 50022
rect 54220 50000 54516 50020
rect 54220 48988 54516 49008
rect 54276 48986 54300 48988
rect 54356 48986 54380 48988
rect 54436 48986 54460 48988
rect 54298 48934 54300 48986
rect 54362 48934 54374 48986
rect 54436 48934 54438 48986
rect 54276 48932 54300 48934
rect 54356 48932 54380 48934
rect 54436 48932 54460 48934
rect 54220 48912 54516 48932
rect 54220 47900 54516 47920
rect 54276 47898 54300 47900
rect 54356 47898 54380 47900
rect 54436 47898 54460 47900
rect 54298 47846 54300 47898
rect 54362 47846 54374 47898
rect 54436 47846 54438 47898
rect 54276 47844 54300 47846
rect 54356 47844 54380 47846
rect 54436 47844 54460 47846
rect 54220 47824 54516 47844
rect 54220 46812 54516 46832
rect 54276 46810 54300 46812
rect 54356 46810 54380 46812
rect 54436 46810 54460 46812
rect 54298 46758 54300 46810
rect 54362 46758 54374 46810
rect 54436 46758 54438 46810
rect 54276 46756 54300 46758
rect 54356 46756 54380 46758
rect 54436 46756 54460 46758
rect 54220 46736 54516 46756
rect 54220 45724 54516 45744
rect 54276 45722 54300 45724
rect 54356 45722 54380 45724
rect 54436 45722 54460 45724
rect 54298 45670 54300 45722
rect 54362 45670 54374 45722
rect 54436 45670 54438 45722
rect 54276 45668 54300 45670
rect 54356 45668 54380 45670
rect 54436 45668 54460 45670
rect 54220 45648 54516 45668
rect 54220 44636 54516 44656
rect 54276 44634 54300 44636
rect 54356 44634 54380 44636
rect 54436 44634 54460 44636
rect 54298 44582 54300 44634
rect 54362 44582 54374 44634
rect 54436 44582 54438 44634
rect 54276 44580 54300 44582
rect 54356 44580 54380 44582
rect 54436 44580 54460 44582
rect 54220 44560 54516 44580
rect 54220 43548 54516 43568
rect 54276 43546 54300 43548
rect 54356 43546 54380 43548
rect 54436 43546 54460 43548
rect 54298 43494 54300 43546
rect 54362 43494 54374 43546
rect 54436 43494 54438 43546
rect 54276 43492 54300 43494
rect 54356 43492 54380 43494
rect 54436 43492 54460 43494
rect 54220 43472 54516 43492
rect 54220 42460 54516 42480
rect 54276 42458 54300 42460
rect 54356 42458 54380 42460
rect 54436 42458 54460 42460
rect 54298 42406 54300 42458
rect 54362 42406 54374 42458
rect 54436 42406 54438 42458
rect 54276 42404 54300 42406
rect 54356 42404 54380 42406
rect 54436 42404 54460 42406
rect 54220 42384 54516 42404
rect 53472 42016 53524 42022
rect 53472 41958 53524 41964
rect 53288 19712 53340 19718
rect 53288 19654 53340 19660
rect 53300 12850 53328 19654
rect 53288 12844 53340 12850
rect 53288 12786 53340 12792
rect 53484 12434 53512 41958
rect 54220 41372 54516 41392
rect 54276 41370 54300 41372
rect 54356 41370 54380 41372
rect 54436 41370 54460 41372
rect 54298 41318 54300 41370
rect 54362 41318 54374 41370
rect 54436 41318 54438 41370
rect 54276 41316 54300 41318
rect 54356 41316 54380 41318
rect 54436 41316 54460 41318
rect 54220 41296 54516 41316
rect 54220 40284 54516 40304
rect 54276 40282 54300 40284
rect 54356 40282 54380 40284
rect 54436 40282 54460 40284
rect 54298 40230 54300 40282
rect 54362 40230 54374 40282
rect 54436 40230 54438 40282
rect 54276 40228 54300 40230
rect 54356 40228 54380 40230
rect 54436 40228 54460 40230
rect 54220 40208 54516 40228
rect 54220 39196 54516 39216
rect 54276 39194 54300 39196
rect 54356 39194 54380 39196
rect 54436 39194 54460 39196
rect 54298 39142 54300 39194
rect 54362 39142 54374 39194
rect 54436 39142 54438 39194
rect 54276 39140 54300 39142
rect 54356 39140 54380 39142
rect 54436 39140 54460 39142
rect 54220 39120 54516 39140
rect 54220 38108 54516 38128
rect 54276 38106 54300 38108
rect 54356 38106 54380 38108
rect 54436 38106 54460 38108
rect 54298 38054 54300 38106
rect 54362 38054 54374 38106
rect 54436 38054 54438 38106
rect 54276 38052 54300 38054
rect 54356 38052 54380 38054
rect 54436 38052 54460 38054
rect 54220 38032 54516 38052
rect 54220 37020 54516 37040
rect 54276 37018 54300 37020
rect 54356 37018 54380 37020
rect 54436 37018 54460 37020
rect 54298 36966 54300 37018
rect 54362 36966 54374 37018
rect 54436 36966 54438 37018
rect 54276 36964 54300 36966
rect 54356 36964 54380 36966
rect 54436 36964 54460 36966
rect 54220 36944 54516 36964
rect 54220 35932 54516 35952
rect 54276 35930 54300 35932
rect 54356 35930 54380 35932
rect 54436 35930 54460 35932
rect 54298 35878 54300 35930
rect 54362 35878 54374 35930
rect 54436 35878 54438 35930
rect 54276 35876 54300 35878
rect 54356 35876 54380 35878
rect 54436 35876 54460 35878
rect 54220 35856 54516 35876
rect 54220 34844 54516 34864
rect 54276 34842 54300 34844
rect 54356 34842 54380 34844
rect 54436 34842 54460 34844
rect 54298 34790 54300 34842
rect 54362 34790 54374 34842
rect 54436 34790 54438 34842
rect 54276 34788 54300 34790
rect 54356 34788 54380 34790
rect 54436 34788 54460 34790
rect 54220 34768 54516 34788
rect 54220 33756 54516 33776
rect 54276 33754 54300 33756
rect 54356 33754 54380 33756
rect 54436 33754 54460 33756
rect 54298 33702 54300 33754
rect 54362 33702 54374 33754
rect 54436 33702 54438 33754
rect 54276 33700 54300 33702
rect 54356 33700 54380 33702
rect 54436 33700 54460 33702
rect 54220 33680 54516 33700
rect 54220 32668 54516 32688
rect 54276 32666 54300 32668
rect 54356 32666 54380 32668
rect 54436 32666 54460 32668
rect 54298 32614 54300 32666
rect 54362 32614 54374 32666
rect 54436 32614 54438 32666
rect 54276 32612 54300 32614
rect 54356 32612 54380 32614
rect 54436 32612 54460 32614
rect 54220 32592 54516 32612
rect 54220 31580 54516 31600
rect 54276 31578 54300 31580
rect 54356 31578 54380 31580
rect 54436 31578 54460 31580
rect 54298 31526 54300 31578
rect 54362 31526 54374 31578
rect 54436 31526 54438 31578
rect 54276 31524 54300 31526
rect 54356 31524 54380 31526
rect 54436 31524 54460 31526
rect 54220 31504 54516 31524
rect 54220 30492 54516 30512
rect 54276 30490 54300 30492
rect 54356 30490 54380 30492
rect 54436 30490 54460 30492
rect 54298 30438 54300 30490
rect 54362 30438 54374 30490
rect 54436 30438 54438 30490
rect 54276 30436 54300 30438
rect 54356 30436 54380 30438
rect 54436 30436 54460 30438
rect 54220 30416 54516 30436
rect 54772 29714 54800 66982
rect 56508 66836 56560 66842
rect 56508 66778 56560 66784
rect 55220 65000 55272 65006
rect 55220 64942 55272 64948
rect 55036 62144 55088 62150
rect 55036 62086 55088 62092
rect 54760 29708 54812 29714
rect 54760 29650 54812 29656
rect 54220 29404 54516 29424
rect 54276 29402 54300 29404
rect 54356 29402 54380 29404
rect 54436 29402 54460 29404
rect 54298 29350 54300 29402
rect 54362 29350 54374 29402
rect 54436 29350 54438 29402
rect 54276 29348 54300 29350
rect 54356 29348 54380 29350
rect 54436 29348 54460 29350
rect 54220 29328 54516 29348
rect 54220 28316 54516 28336
rect 54276 28314 54300 28316
rect 54356 28314 54380 28316
rect 54436 28314 54460 28316
rect 54298 28262 54300 28314
rect 54362 28262 54374 28314
rect 54436 28262 54438 28314
rect 54276 28260 54300 28262
rect 54356 28260 54380 28262
rect 54436 28260 54460 28262
rect 54220 28240 54516 28260
rect 54220 27228 54516 27248
rect 54276 27226 54300 27228
rect 54356 27226 54380 27228
rect 54436 27226 54460 27228
rect 54298 27174 54300 27226
rect 54362 27174 54374 27226
rect 54436 27174 54438 27226
rect 54276 27172 54300 27174
rect 54356 27172 54380 27174
rect 54436 27172 54460 27174
rect 54220 27152 54516 27172
rect 54576 27056 54628 27062
rect 54576 26998 54628 27004
rect 53840 26988 53892 26994
rect 53840 26930 53892 26936
rect 53852 23594 53880 26930
rect 54220 26140 54516 26160
rect 54276 26138 54300 26140
rect 54356 26138 54380 26140
rect 54436 26138 54460 26140
rect 54298 26086 54300 26138
rect 54362 26086 54374 26138
rect 54436 26086 54438 26138
rect 54276 26084 54300 26086
rect 54356 26084 54380 26086
rect 54436 26084 54460 26086
rect 54220 26064 54516 26084
rect 54220 25052 54516 25072
rect 54276 25050 54300 25052
rect 54356 25050 54380 25052
rect 54436 25050 54460 25052
rect 54298 24998 54300 25050
rect 54362 24998 54374 25050
rect 54436 24998 54438 25050
rect 54276 24996 54300 24998
rect 54356 24996 54380 24998
rect 54436 24996 54460 24998
rect 54220 24976 54516 24996
rect 54116 24064 54168 24070
rect 54116 24006 54168 24012
rect 54128 23866 54156 24006
rect 54220 23964 54516 23984
rect 54276 23962 54300 23964
rect 54356 23962 54380 23964
rect 54436 23962 54460 23964
rect 54298 23910 54300 23962
rect 54362 23910 54374 23962
rect 54436 23910 54438 23962
rect 54276 23908 54300 23910
rect 54356 23908 54380 23910
rect 54436 23908 54460 23910
rect 54220 23888 54516 23908
rect 54116 23860 54168 23866
rect 54116 23802 54168 23808
rect 54392 23656 54444 23662
rect 54392 23598 54444 23604
rect 53840 23588 53892 23594
rect 53840 23530 53892 23536
rect 54404 23526 54432 23598
rect 53932 23520 53984 23526
rect 53932 23462 53984 23468
rect 54392 23520 54444 23526
rect 54392 23462 54444 23468
rect 53944 23254 53972 23462
rect 53932 23248 53984 23254
rect 53932 23190 53984 23196
rect 54116 23044 54168 23050
rect 54116 22986 54168 22992
rect 53932 17128 53984 17134
rect 53932 17070 53984 17076
rect 53748 14952 53800 14958
rect 53748 14894 53800 14900
rect 53392 12406 53512 12434
rect 53196 11756 53248 11762
rect 53196 11698 53248 11704
rect 52000 8832 52052 8838
rect 52000 8774 52052 8780
rect 52460 8832 52512 8838
rect 52460 8774 52512 8780
rect 53012 8832 53064 8838
rect 53012 8774 53064 8780
rect 51816 8628 51868 8634
rect 51816 8570 51868 8576
rect 51908 8628 51960 8634
rect 51908 8570 51960 8576
rect 51724 7268 51776 7274
rect 51724 7210 51776 7216
rect 51736 5778 51764 7210
rect 51816 6656 51868 6662
rect 51816 6598 51868 6604
rect 51724 5772 51776 5778
rect 51724 5714 51776 5720
rect 51724 5636 51776 5642
rect 51724 5578 51776 5584
rect 51736 3466 51764 5578
rect 51828 3602 51856 6598
rect 51920 5166 51948 8570
rect 52012 5642 52040 8774
rect 52276 8356 52328 8362
rect 52276 8298 52328 8304
rect 52092 7744 52144 7750
rect 52092 7686 52144 7692
rect 52000 5636 52052 5642
rect 52000 5578 52052 5584
rect 52104 5166 52132 7686
rect 52184 7200 52236 7206
rect 52184 7142 52236 7148
rect 51908 5160 51960 5166
rect 51908 5102 51960 5108
rect 52092 5160 52144 5166
rect 52092 5102 52144 5108
rect 52000 5024 52052 5030
rect 52000 4966 52052 4972
rect 51908 4820 51960 4826
rect 51908 4762 51960 4768
rect 51816 3596 51868 3602
rect 51816 3538 51868 3544
rect 51724 3460 51776 3466
rect 51724 3402 51776 3408
rect 51828 3398 51856 3538
rect 51816 3392 51868 3398
rect 51816 3334 51868 3340
rect 51724 3052 51776 3058
rect 51724 2994 51776 3000
rect 51632 2576 51684 2582
rect 51632 2518 51684 2524
rect 51736 800 51764 2994
rect 51920 2990 51948 4762
rect 52012 3670 52040 4966
rect 52196 4690 52224 7142
rect 52288 4826 52316 8298
rect 52368 7744 52420 7750
rect 52368 7686 52420 7692
rect 52380 5778 52408 7686
rect 52368 5772 52420 5778
rect 52368 5714 52420 5720
rect 52368 5636 52420 5642
rect 52368 5578 52420 5584
rect 52276 4820 52328 4826
rect 52276 4762 52328 4768
rect 52380 4706 52408 5578
rect 52184 4684 52236 4690
rect 52184 4626 52236 4632
rect 52288 4678 52408 4706
rect 52092 4072 52144 4078
rect 52092 4014 52144 4020
rect 52000 3664 52052 3670
rect 52000 3606 52052 3612
rect 51908 2984 51960 2990
rect 51908 2926 51960 2932
rect 51816 2916 51868 2922
rect 51816 2858 51868 2864
rect 51828 800 51856 2858
rect 52104 2774 52132 4014
rect 52196 3942 52224 4626
rect 52184 3936 52236 3942
rect 52184 3878 52236 3884
rect 52288 3534 52316 4678
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52012 2746 52132 2774
rect 52012 800 52040 2746
rect 52274 2544 52330 2553
rect 52184 2508 52236 2514
rect 52274 2479 52330 2488
rect 52184 2450 52236 2456
rect 52092 2372 52144 2378
rect 52092 2314 52144 2320
rect 52104 800 52132 2314
rect 52196 1222 52224 2450
rect 52184 1216 52236 1222
rect 52184 1158 52236 1164
rect 52288 800 52316 2479
rect 52380 800 52408 3334
rect 52472 2990 52500 8774
rect 52828 7744 52880 7750
rect 52828 7686 52880 7692
rect 52552 6656 52604 6662
rect 52552 6598 52604 6604
rect 52564 4078 52592 6598
rect 52644 6112 52696 6118
rect 52644 6054 52696 6060
rect 52656 4146 52684 6054
rect 52840 5778 52868 7686
rect 52920 7200 52972 7206
rect 52920 7142 52972 7148
rect 52828 5772 52880 5778
rect 52828 5714 52880 5720
rect 52840 5658 52868 5714
rect 52932 5710 52960 7142
rect 52748 5630 52868 5658
rect 52920 5704 52972 5710
rect 52920 5646 52972 5652
rect 52644 4140 52696 4146
rect 52644 4082 52696 4088
rect 52552 4072 52604 4078
rect 52552 4014 52604 4020
rect 52552 3460 52604 3466
rect 52552 3402 52604 3408
rect 52460 2984 52512 2990
rect 52460 2926 52512 2932
rect 52564 800 52592 3402
rect 52748 800 52776 5630
rect 52828 4684 52880 4690
rect 52828 4626 52880 4632
rect 52840 800 52868 4626
rect 52932 2922 52960 5646
rect 53024 3602 53052 8774
rect 53392 8362 53420 12406
rect 53380 8356 53432 8362
rect 53380 8298 53432 8304
rect 53196 6656 53248 6662
rect 53196 6598 53248 6604
rect 53104 5704 53156 5710
rect 53104 5646 53156 5652
rect 53012 3596 53064 3602
rect 53012 3538 53064 3544
rect 52920 2916 52972 2922
rect 52920 2858 52972 2864
rect 53012 2916 53064 2922
rect 53012 2858 53064 2864
rect 53024 800 53052 2858
rect 53116 800 53144 5646
rect 53208 4690 53236 6598
rect 53288 6112 53340 6118
rect 53288 6054 53340 6060
rect 53196 4684 53248 4690
rect 53196 4626 53248 4632
rect 53300 4570 53328 6054
rect 53208 4542 53328 4570
rect 53208 3398 53236 4542
rect 53392 3670 53420 8298
rect 53760 7750 53788 14894
rect 53840 13796 53892 13802
rect 53840 13738 53892 13744
rect 53852 12986 53880 13738
rect 53840 12980 53892 12986
rect 53840 12922 53892 12928
rect 53944 12646 53972 17070
rect 53932 12640 53984 12646
rect 53932 12582 53984 12588
rect 54128 8838 54156 22986
rect 54220 22876 54516 22896
rect 54276 22874 54300 22876
rect 54356 22874 54380 22876
rect 54436 22874 54460 22876
rect 54298 22822 54300 22874
rect 54362 22822 54374 22874
rect 54436 22822 54438 22874
rect 54276 22820 54300 22822
rect 54356 22820 54380 22822
rect 54436 22820 54460 22822
rect 54220 22800 54516 22820
rect 54220 21788 54516 21808
rect 54276 21786 54300 21788
rect 54356 21786 54380 21788
rect 54436 21786 54460 21788
rect 54298 21734 54300 21786
rect 54362 21734 54374 21786
rect 54436 21734 54438 21786
rect 54276 21732 54300 21734
rect 54356 21732 54380 21734
rect 54436 21732 54460 21734
rect 54220 21712 54516 21732
rect 54220 20700 54516 20720
rect 54276 20698 54300 20700
rect 54356 20698 54380 20700
rect 54436 20698 54460 20700
rect 54298 20646 54300 20698
rect 54362 20646 54374 20698
rect 54436 20646 54438 20698
rect 54276 20644 54300 20646
rect 54356 20644 54380 20646
rect 54436 20644 54460 20646
rect 54220 20624 54516 20644
rect 54220 19612 54516 19632
rect 54276 19610 54300 19612
rect 54356 19610 54380 19612
rect 54436 19610 54460 19612
rect 54298 19558 54300 19610
rect 54362 19558 54374 19610
rect 54436 19558 54438 19610
rect 54276 19556 54300 19558
rect 54356 19556 54380 19558
rect 54436 19556 54460 19558
rect 54220 19536 54516 19556
rect 54220 18524 54516 18544
rect 54276 18522 54300 18524
rect 54356 18522 54380 18524
rect 54436 18522 54460 18524
rect 54298 18470 54300 18522
rect 54362 18470 54374 18522
rect 54436 18470 54438 18522
rect 54276 18468 54300 18470
rect 54356 18468 54380 18470
rect 54436 18468 54460 18470
rect 54220 18448 54516 18468
rect 54220 17436 54516 17456
rect 54276 17434 54300 17436
rect 54356 17434 54380 17436
rect 54436 17434 54460 17436
rect 54298 17382 54300 17434
rect 54362 17382 54374 17434
rect 54436 17382 54438 17434
rect 54276 17380 54300 17382
rect 54356 17380 54380 17382
rect 54436 17380 54460 17382
rect 54220 17360 54516 17380
rect 54220 16348 54516 16368
rect 54276 16346 54300 16348
rect 54356 16346 54380 16348
rect 54436 16346 54460 16348
rect 54298 16294 54300 16346
rect 54362 16294 54374 16346
rect 54436 16294 54438 16346
rect 54276 16292 54300 16294
rect 54356 16292 54380 16294
rect 54436 16292 54460 16294
rect 54220 16272 54516 16292
rect 54220 15260 54516 15280
rect 54276 15258 54300 15260
rect 54356 15258 54380 15260
rect 54436 15258 54460 15260
rect 54298 15206 54300 15258
rect 54362 15206 54374 15258
rect 54436 15206 54438 15258
rect 54276 15204 54300 15206
rect 54356 15204 54380 15206
rect 54436 15204 54460 15206
rect 54220 15184 54516 15204
rect 54220 14172 54516 14192
rect 54276 14170 54300 14172
rect 54356 14170 54380 14172
rect 54436 14170 54460 14172
rect 54298 14118 54300 14170
rect 54362 14118 54374 14170
rect 54436 14118 54438 14170
rect 54276 14116 54300 14118
rect 54356 14116 54380 14118
rect 54436 14116 54460 14118
rect 54220 14096 54516 14116
rect 54220 13084 54516 13104
rect 54276 13082 54300 13084
rect 54356 13082 54380 13084
rect 54436 13082 54460 13084
rect 54298 13030 54300 13082
rect 54362 13030 54374 13082
rect 54436 13030 54438 13082
rect 54276 13028 54300 13030
rect 54356 13028 54380 13030
rect 54436 13028 54460 13030
rect 54220 13008 54516 13028
rect 54588 12434 54616 26998
rect 54760 24132 54812 24138
rect 54760 24074 54812 24080
rect 54772 23526 54800 24074
rect 54760 23520 54812 23526
rect 54760 23462 54812 23468
rect 54944 17060 54996 17066
rect 54944 17002 54996 17008
rect 54956 12434 54984 17002
rect 54588 12406 54708 12434
rect 54220 11996 54516 12016
rect 54276 11994 54300 11996
rect 54356 11994 54380 11996
rect 54436 11994 54460 11996
rect 54298 11942 54300 11994
rect 54362 11942 54374 11994
rect 54436 11942 54438 11994
rect 54276 11940 54300 11942
rect 54356 11940 54380 11942
rect 54436 11940 54460 11942
rect 54220 11920 54516 11940
rect 54220 10908 54516 10928
rect 54276 10906 54300 10908
rect 54356 10906 54380 10908
rect 54436 10906 54460 10908
rect 54298 10854 54300 10906
rect 54362 10854 54374 10906
rect 54436 10854 54438 10906
rect 54276 10852 54300 10854
rect 54356 10852 54380 10854
rect 54436 10852 54460 10854
rect 54220 10832 54516 10852
rect 54220 9820 54516 9840
rect 54276 9818 54300 9820
rect 54356 9818 54380 9820
rect 54436 9818 54460 9820
rect 54298 9766 54300 9818
rect 54362 9766 54374 9818
rect 54436 9766 54438 9818
rect 54276 9764 54300 9766
rect 54356 9764 54380 9766
rect 54436 9764 54460 9766
rect 54220 9744 54516 9764
rect 54116 8832 54168 8838
rect 54116 8774 54168 8780
rect 54024 8628 54076 8634
rect 54024 8570 54076 8576
rect 53472 7744 53524 7750
rect 53472 7686 53524 7692
rect 53748 7744 53800 7750
rect 53748 7686 53800 7692
rect 53380 3664 53432 3670
rect 53380 3606 53432 3612
rect 53288 3528 53340 3534
rect 53288 3470 53340 3476
rect 53196 3392 53248 3398
rect 53196 3334 53248 3340
rect 53300 800 53328 3470
rect 53380 3460 53432 3466
rect 53380 3402 53432 3408
rect 53392 800 53420 3402
rect 53484 2582 53512 7686
rect 53840 7268 53892 7274
rect 53840 7210 53892 7216
rect 53748 7200 53800 7206
rect 53748 7142 53800 7148
rect 53760 5166 53788 7142
rect 53748 5160 53800 5166
rect 53748 5102 53800 5108
rect 53760 5001 53788 5102
rect 53852 5098 53880 7210
rect 53932 6656 53984 6662
rect 53932 6598 53984 6604
rect 53840 5092 53892 5098
rect 53840 5034 53892 5040
rect 53746 4992 53802 5001
rect 53746 4927 53802 4936
rect 53852 4842 53880 5034
rect 53576 4814 53880 4842
rect 53472 2576 53524 2582
rect 53472 2518 53524 2524
rect 53576 800 53604 4814
rect 53944 4690 53972 6598
rect 53932 4684 53984 4690
rect 53852 4644 53932 4672
rect 53852 4128 53880 4644
rect 53932 4626 53984 4632
rect 53932 4480 53984 4486
rect 53932 4422 53984 4428
rect 53668 4100 53880 4128
rect 53668 800 53696 4100
rect 53944 4060 53972 4422
rect 53852 4032 53972 4060
rect 53748 4004 53800 4010
rect 53748 3946 53800 3952
rect 53760 3398 53788 3946
rect 53748 3392 53800 3398
rect 53748 3334 53800 3340
rect 53852 3210 53880 4032
rect 53932 3936 53984 3942
rect 53932 3878 53984 3884
rect 53760 3182 53880 3210
rect 53760 2582 53788 3182
rect 53840 3052 53892 3058
rect 53840 2994 53892 3000
rect 53748 2576 53800 2582
rect 53748 2518 53800 2524
rect 53852 800 53880 2994
rect 53944 1034 53972 3878
rect 54036 2990 54064 8570
rect 54128 3670 54156 8774
rect 54220 8732 54516 8752
rect 54276 8730 54300 8732
rect 54356 8730 54380 8732
rect 54436 8730 54460 8732
rect 54298 8678 54300 8730
rect 54362 8678 54374 8730
rect 54436 8678 54438 8730
rect 54276 8676 54300 8678
rect 54356 8676 54380 8678
rect 54436 8676 54460 8678
rect 54220 8656 54516 8676
rect 54680 8362 54708 12406
rect 54864 12406 54984 12434
rect 54668 8356 54720 8362
rect 54668 8298 54720 8304
rect 54220 7644 54516 7664
rect 54276 7642 54300 7644
rect 54356 7642 54380 7644
rect 54436 7642 54460 7644
rect 54298 7590 54300 7642
rect 54362 7590 54374 7642
rect 54436 7590 54438 7642
rect 54276 7588 54300 7590
rect 54356 7588 54380 7590
rect 54436 7588 54460 7590
rect 54220 7568 54516 7588
rect 54576 6656 54628 6662
rect 54576 6598 54628 6604
rect 54220 6556 54516 6576
rect 54276 6554 54300 6556
rect 54356 6554 54380 6556
rect 54436 6554 54460 6556
rect 54298 6502 54300 6554
rect 54362 6502 54374 6554
rect 54436 6502 54438 6554
rect 54276 6500 54300 6502
rect 54356 6500 54380 6502
rect 54436 6500 54460 6502
rect 54220 6480 54516 6500
rect 54220 5468 54516 5488
rect 54276 5466 54300 5468
rect 54356 5466 54380 5468
rect 54436 5466 54460 5468
rect 54298 5414 54300 5466
rect 54362 5414 54374 5466
rect 54436 5414 54438 5466
rect 54276 5412 54300 5414
rect 54356 5412 54380 5414
rect 54436 5412 54460 5414
rect 54220 5392 54516 5412
rect 54588 4690 54616 6598
rect 54576 4684 54628 4690
rect 54576 4626 54628 4632
rect 54220 4380 54516 4400
rect 54276 4378 54300 4380
rect 54356 4378 54380 4380
rect 54436 4378 54460 4380
rect 54298 4326 54300 4378
rect 54362 4326 54374 4378
rect 54436 4326 54438 4378
rect 54276 4324 54300 4326
rect 54356 4324 54380 4326
rect 54436 4324 54460 4326
rect 54220 4304 54516 4324
rect 54116 3664 54168 3670
rect 54116 3606 54168 3612
rect 54116 3460 54168 3466
rect 54116 3402 54168 3408
rect 54024 2984 54076 2990
rect 54024 2926 54076 2932
rect 54128 1442 54156 3402
rect 54220 3292 54516 3312
rect 54276 3290 54300 3292
rect 54356 3290 54380 3292
rect 54436 3290 54460 3292
rect 54298 3238 54300 3290
rect 54362 3238 54374 3290
rect 54436 3238 54438 3290
rect 54276 3236 54300 3238
rect 54356 3236 54380 3238
rect 54436 3236 54460 3238
rect 54220 3216 54516 3236
rect 54208 3120 54260 3126
rect 54208 3062 54260 3068
rect 54220 2650 54248 3062
rect 54484 2848 54536 2854
rect 54484 2790 54536 2796
rect 54208 2644 54260 2650
rect 54208 2586 54260 2592
rect 54496 2582 54524 2790
rect 54484 2576 54536 2582
rect 54484 2518 54536 2524
rect 54220 2204 54516 2224
rect 54276 2202 54300 2204
rect 54356 2202 54380 2204
rect 54436 2202 54460 2204
rect 54298 2150 54300 2202
rect 54362 2150 54374 2202
rect 54436 2150 54438 2202
rect 54276 2148 54300 2150
rect 54356 2148 54380 2150
rect 54436 2148 54460 2150
rect 54220 2128 54516 2148
rect 54390 2000 54446 2009
rect 54390 1935 54446 1944
rect 54128 1414 54340 1442
rect 53944 1006 54156 1034
rect 53932 944 53984 950
rect 53932 886 53984 892
rect 53944 800 53972 886
rect 54128 800 54156 1006
rect 54312 800 54340 1414
rect 54404 800 54432 1935
rect 54588 800 54616 4626
rect 54680 2990 54708 8298
rect 54864 7750 54892 12406
rect 55048 8634 55076 62086
rect 55128 57792 55180 57798
rect 55128 57734 55180 57740
rect 55140 14074 55168 57734
rect 55128 14068 55180 14074
rect 55128 14010 55180 14016
rect 55036 8628 55088 8634
rect 55036 8570 55088 8576
rect 55232 8362 55260 64942
rect 56520 60178 56548 66778
rect 57808 66706 57836 67050
rect 62580 67040 62632 67046
rect 62580 66982 62632 66988
rect 64604 67040 64656 67046
rect 64604 66982 64656 66988
rect 59220 66940 59516 66960
rect 59276 66938 59300 66940
rect 59356 66938 59380 66940
rect 59436 66938 59460 66940
rect 59298 66886 59300 66938
rect 59362 66886 59374 66938
rect 59436 66886 59438 66938
rect 59276 66884 59300 66886
rect 59356 66884 59380 66886
rect 59436 66884 59460 66886
rect 59220 66864 59516 66884
rect 57796 66700 57848 66706
rect 57796 66642 57848 66648
rect 62592 66638 62620 66982
rect 62580 66632 62632 66638
rect 62580 66574 62632 66580
rect 64220 66396 64516 66416
rect 64276 66394 64300 66396
rect 64356 66394 64380 66396
rect 64436 66394 64460 66396
rect 64298 66342 64300 66394
rect 64362 66342 64374 66394
rect 64436 66342 64438 66394
rect 64276 66340 64300 66342
rect 64356 66340 64380 66342
rect 64436 66340 64460 66342
rect 64220 66320 64516 66340
rect 61476 66292 61528 66298
rect 61476 66234 61528 66240
rect 59220 65852 59516 65872
rect 59276 65850 59300 65852
rect 59356 65850 59380 65852
rect 59436 65850 59460 65852
rect 59298 65798 59300 65850
rect 59362 65798 59374 65850
rect 59436 65798 59438 65850
rect 59276 65796 59300 65798
rect 59356 65796 59380 65798
rect 59436 65796 59460 65798
rect 59220 65776 59516 65796
rect 56784 65408 56836 65414
rect 56784 65350 56836 65356
rect 56508 60172 56560 60178
rect 56508 60114 56560 60120
rect 55588 53440 55640 53446
rect 55588 53382 55640 53388
rect 55864 53440 55916 53446
rect 55864 53382 55916 53388
rect 55600 53038 55628 53382
rect 55588 53032 55640 53038
rect 55588 52974 55640 52980
rect 55600 52698 55628 52974
rect 55588 52692 55640 52698
rect 55588 52634 55640 52640
rect 55312 52488 55364 52494
rect 55312 52430 55364 52436
rect 55324 43994 55352 52430
rect 55312 43988 55364 43994
rect 55312 43930 55364 43936
rect 55680 38752 55732 38758
rect 55680 38694 55732 38700
rect 55312 33856 55364 33862
rect 55312 33798 55364 33804
rect 55324 13394 55352 33798
rect 55692 31958 55720 38694
rect 55680 31952 55732 31958
rect 55680 31894 55732 31900
rect 55404 21412 55456 21418
rect 55404 21354 55456 21360
rect 55312 13388 55364 13394
rect 55312 13330 55364 13336
rect 55220 8356 55272 8362
rect 55220 8298 55272 8304
rect 54852 7744 54904 7750
rect 54852 7686 54904 7692
rect 54760 6112 54812 6118
rect 54760 6054 54812 6060
rect 54772 4078 54800 6054
rect 54864 4486 54892 7686
rect 55036 7200 55088 7206
rect 55036 7142 55088 7148
rect 54944 6656 54996 6662
rect 54944 6598 54996 6604
rect 54956 5710 54984 6598
rect 55048 5778 55076 7142
rect 55128 6112 55180 6118
rect 55128 6054 55180 6060
rect 55036 5772 55088 5778
rect 55036 5714 55088 5720
rect 54944 5704 54996 5710
rect 54944 5646 54996 5652
rect 54944 5160 54996 5166
rect 54944 5102 54996 5108
rect 54956 5001 54984 5102
rect 54942 4992 54998 5001
rect 54942 4927 54998 4936
rect 54852 4480 54904 4486
rect 54852 4422 54904 4428
rect 54852 4140 54904 4146
rect 54852 4082 54904 4088
rect 54760 4072 54812 4078
rect 54760 4014 54812 4020
rect 54772 3534 54800 4014
rect 54760 3528 54812 3534
rect 54760 3470 54812 3476
rect 54668 2984 54720 2990
rect 54668 2926 54720 2932
rect 54760 2848 54812 2854
rect 54680 2808 54760 2836
rect 54680 800 54708 2808
rect 54760 2790 54812 2796
rect 54864 800 54892 4082
rect 54944 4004 54996 4010
rect 54944 3946 54996 3952
rect 54956 800 54984 3946
rect 55048 950 55076 5714
rect 55140 4078 55168 6054
rect 55128 4072 55180 4078
rect 55128 4014 55180 4020
rect 55128 3460 55180 3466
rect 55128 3402 55180 3408
rect 55036 944 55088 950
rect 55036 886 55088 892
rect 55140 800 55168 3402
rect 55232 2922 55260 8298
rect 55416 8090 55444 21354
rect 55876 14278 55904 53382
rect 55956 50856 56008 50862
rect 55956 50798 56008 50804
rect 55968 14482 55996 50798
rect 56048 43988 56100 43994
rect 56048 43930 56100 43936
rect 56060 43790 56088 43930
rect 56048 43784 56100 43790
rect 56048 43726 56100 43732
rect 56060 34950 56088 43726
rect 56048 34944 56100 34950
rect 56048 34886 56100 34892
rect 56232 31884 56284 31890
rect 56232 31826 56284 31832
rect 56244 21622 56272 31826
rect 56416 25764 56468 25770
rect 56416 25706 56468 25712
rect 56232 21616 56284 21622
rect 56232 21558 56284 21564
rect 56428 21162 56456 25706
rect 56508 23520 56560 23526
rect 56508 23462 56560 23468
rect 56520 23118 56548 23462
rect 56508 23112 56560 23118
rect 56508 23054 56560 23060
rect 56520 22642 56548 23054
rect 56508 22636 56560 22642
rect 56508 22578 56560 22584
rect 56428 21134 56548 21162
rect 56048 17536 56100 17542
rect 56048 17478 56100 17484
rect 55956 14476 56008 14482
rect 55956 14418 56008 14424
rect 55864 14272 55916 14278
rect 55864 14214 55916 14220
rect 55680 13252 55732 13258
rect 55680 13194 55732 13200
rect 55692 8362 55720 13194
rect 55680 8356 55732 8362
rect 55680 8298 55732 8304
rect 55404 8084 55456 8090
rect 55324 8044 55404 8072
rect 55220 2916 55272 2922
rect 55220 2858 55272 2864
rect 55324 2582 55352 8044
rect 55404 8026 55456 8032
rect 55496 7200 55548 7206
rect 55496 7142 55548 7148
rect 55404 6656 55456 6662
rect 55404 6598 55456 6604
rect 55416 5166 55444 6598
rect 55508 5778 55536 7142
rect 55588 6112 55640 6118
rect 55588 6054 55640 6060
rect 55496 5772 55548 5778
rect 55496 5714 55548 5720
rect 55404 5160 55456 5166
rect 55404 5102 55456 5108
rect 55404 4684 55456 4690
rect 55404 4626 55456 4632
rect 55312 2576 55364 2582
rect 55312 2518 55364 2524
rect 55220 1420 55272 1426
rect 55220 1362 55272 1368
rect 55232 800 55260 1362
rect 55416 800 55444 4626
rect 55508 4146 55536 5714
rect 55496 4140 55548 4146
rect 55496 4082 55548 4088
rect 55600 4078 55628 6054
rect 55588 4072 55640 4078
rect 55588 4014 55640 4020
rect 55588 3936 55640 3942
rect 55588 3878 55640 3884
rect 55496 3052 55548 3058
rect 55496 2994 55548 3000
rect 55508 800 55536 2994
rect 55600 1426 55628 3878
rect 55692 3670 55720 8298
rect 56060 8090 56088 17478
rect 56140 16652 56192 16658
rect 56140 16594 56192 16600
rect 56152 16250 56180 16594
rect 56520 16522 56548 21134
rect 56508 16516 56560 16522
rect 56508 16458 56560 16464
rect 56140 16244 56192 16250
rect 56140 16186 56192 16192
rect 56152 15910 56180 16186
rect 56140 15904 56192 15910
rect 56140 15846 56192 15852
rect 56048 8084 56100 8090
rect 56048 8026 56100 8032
rect 55956 7948 56008 7954
rect 55956 7890 56008 7896
rect 55968 7750 55996 7890
rect 55956 7744 56008 7750
rect 55956 7686 56008 7692
rect 55864 6248 55916 6254
rect 55864 6190 55916 6196
rect 55772 5092 55824 5098
rect 55772 5034 55824 5040
rect 55680 3664 55732 3670
rect 55680 3606 55732 3612
rect 55784 3482 55812 5034
rect 55876 4214 55904 6190
rect 55968 5273 55996 7686
rect 55954 5264 56010 5273
rect 55954 5199 56010 5208
rect 55956 5160 56008 5166
rect 55956 5102 56008 5108
rect 55864 4208 55916 4214
rect 55864 4150 55916 4156
rect 55864 4072 55916 4078
rect 55864 4014 55916 4020
rect 55692 3454 55812 3482
rect 55588 1420 55640 1426
rect 55588 1362 55640 1368
rect 55692 800 55720 3454
rect 55876 3380 55904 4014
rect 55968 3942 55996 5102
rect 55956 3936 56008 3942
rect 55956 3878 56008 3884
rect 55954 3768 56010 3777
rect 55954 3703 56010 3712
rect 55784 3352 55904 3380
rect 55784 800 55812 3352
rect 55968 3210 55996 3703
rect 55876 3182 55996 3210
rect 55876 2582 55904 3182
rect 56060 2922 56088 8026
rect 56796 7546 56824 65350
rect 59220 64764 59516 64784
rect 59276 64762 59300 64764
rect 59356 64762 59380 64764
rect 59436 64762 59460 64764
rect 59298 64710 59300 64762
rect 59362 64710 59374 64762
rect 59436 64710 59438 64762
rect 59276 64708 59300 64710
rect 59356 64708 59380 64710
rect 59436 64708 59460 64710
rect 59220 64688 59516 64708
rect 59220 63676 59516 63696
rect 59276 63674 59300 63676
rect 59356 63674 59380 63676
rect 59436 63674 59460 63676
rect 59298 63622 59300 63674
rect 59362 63622 59374 63674
rect 59436 63622 59438 63674
rect 59276 63620 59300 63622
rect 59356 63620 59380 63622
rect 59436 63620 59460 63622
rect 59220 63600 59516 63620
rect 59220 62588 59516 62608
rect 59276 62586 59300 62588
rect 59356 62586 59380 62588
rect 59436 62586 59460 62588
rect 59298 62534 59300 62586
rect 59362 62534 59374 62586
rect 59436 62534 59438 62586
rect 59276 62532 59300 62534
rect 59356 62532 59380 62534
rect 59436 62532 59460 62534
rect 59220 62512 59516 62532
rect 59220 61500 59516 61520
rect 59276 61498 59300 61500
rect 59356 61498 59380 61500
rect 59436 61498 59460 61500
rect 59298 61446 59300 61498
rect 59362 61446 59374 61498
rect 59436 61446 59438 61498
rect 59276 61444 59300 61446
rect 59356 61444 59380 61446
rect 59436 61444 59460 61446
rect 59220 61424 59516 61444
rect 59220 60412 59516 60432
rect 59276 60410 59300 60412
rect 59356 60410 59380 60412
rect 59436 60410 59460 60412
rect 59298 60358 59300 60410
rect 59362 60358 59374 60410
rect 59436 60358 59438 60410
rect 59276 60356 59300 60358
rect 59356 60356 59380 60358
rect 59436 60356 59460 60358
rect 59220 60336 59516 60356
rect 58624 60104 58676 60110
rect 58624 60046 58676 60052
rect 58636 57798 58664 60046
rect 58716 59424 58768 59430
rect 58716 59366 58768 59372
rect 58624 57792 58676 57798
rect 58624 57734 58676 57740
rect 58636 45558 58664 57734
rect 58624 45552 58676 45558
rect 58624 45494 58676 45500
rect 58636 44946 58664 45494
rect 58728 45014 58756 59366
rect 59220 59324 59516 59344
rect 59276 59322 59300 59324
rect 59356 59322 59380 59324
rect 59436 59322 59460 59324
rect 59298 59270 59300 59322
rect 59362 59270 59374 59322
rect 59436 59270 59438 59322
rect 59276 59268 59300 59270
rect 59356 59268 59380 59270
rect 59436 59268 59460 59270
rect 59220 59248 59516 59268
rect 59220 58236 59516 58256
rect 59276 58234 59300 58236
rect 59356 58234 59380 58236
rect 59436 58234 59460 58236
rect 59298 58182 59300 58234
rect 59362 58182 59374 58234
rect 59436 58182 59438 58234
rect 59276 58180 59300 58182
rect 59356 58180 59380 58182
rect 59436 58180 59460 58182
rect 59220 58160 59516 58180
rect 59220 57148 59516 57168
rect 59276 57146 59300 57148
rect 59356 57146 59380 57148
rect 59436 57146 59460 57148
rect 59298 57094 59300 57146
rect 59362 57094 59374 57146
rect 59436 57094 59438 57146
rect 59276 57092 59300 57094
rect 59356 57092 59380 57094
rect 59436 57092 59460 57094
rect 59220 57072 59516 57092
rect 59220 56060 59516 56080
rect 59276 56058 59300 56060
rect 59356 56058 59380 56060
rect 59436 56058 59460 56060
rect 59298 56006 59300 56058
rect 59362 56006 59374 56058
rect 59436 56006 59438 56058
rect 59276 56004 59300 56006
rect 59356 56004 59380 56006
rect 59436 56004 59460 56006
rect 59220 55984 59516 56004
rect 59220 54972 59516 54992
rect 59276 54970 59300 54972
rect 59356 54970 59380 54972
rect 59436 54970 59460 54972
rect 59298 54918 59300 54970
rect 59362 54918 59374 54970
rect 59436 54918 59438 54970
rect 59276 54916 59300 54918
rect 59356 54916 59380 54918
rect 59436 54916 59460 54918
rect 59220 54896 59516 54916
rect 59220 53884 59516 53904
rect 59276 53882 59300 53884
rect 59356 53882 59380 53884
rect 59436 53882 59460 53884
rect 59298 53830 59300 53882
rect 59362 53830 59374 53882
rect 59436 53830 59438 53882
rect 59276 53828 59300 53830
rect 59356 53828 59380 53830
rect 59436 53828 59460 53830
rect 59220 53808 59516 53828
rect 59220 52796 59516 52816
rect 59276 52794 59300 52796
rect 59356 52794 59380 52796
rect 59436 52794 59460 52796
rect 59298 52742 59300 52794
rect 59362 52742 59374 52794
rect 59436 52742 59438 52794
rect 59276 52740 59300 52742
rect 59356 52740 59380 52742
rect 59436 52740 59460 52742
rect 59220 52720 59516 52740
rect 59220 51708 59516 51728
rect 59276 51706 59300 51708
rect 59356 51706 59380 51708
rect 59436 51706 59460 51708
rect 59298 51654 59300 51706
rect 59362 51654 59374 51706
rect 59436 51654 59438 51706
rect 59276 51652 59300 51654
rect 59356 51652 59380 51654
rect 59436 51652 59460 51654
rect 59220 51632 59516 51652
rect 59220 50620 59516 50640
rect 59276 50618 59300 50620
rect 59356 50618 59380 50620
rect 59436 50618 59460 50620
rect 59298 50566 59300 50618
rect 59362 50566 59374 50618
rect 59436 50566 59438 50618
rect 59276 50564 59300 50566
rect 59356 50564 59380 50566
rect 59436 50564 59460 50566
rect 59220 50544 59516 50564
rect 59220 49532 59516 49552
rect 59276 49530 59300 49532
rect 59356 49530 59380 49532
rect 59436 49530 59460 49532
rect 59298 49478 59300 49530
rect 59362 49478 59374 49530
rect 59436 49478 59438 49530
rect 59276 49476 59300 49478
rect 59356 49476 59380 49478
rect 59436 49476 59460 49478
rect 59220 49456 59516 49476
rect 59220 48444 59516 48464
rect 59276 48442 59300 48444
rect 59356 48442 59380 48444
rect 59436 48442 59460 48444
rect 59298 48390 59300 48442
rect 59362 48390 59374 48442
rect 59436 48390 59438 48442
rect 59276 48388 59300 48390
rect 59356 48388 59380 48390
rect 59436 48388 59460 48390
rect 59220 48368 59516 48388
rect 59220 47356 59516 47376
rect 59276 47354 59300 47356
rect 59356 47354 59380 47356
rect 59436 47354 59460 47356
rect 59298 47302 59300 47354
rect 59362 47302 59374 47354
rect 59436 47302 59438 47354
rect 59276 47300 59300 47302
rect 59356 47300 59380 47302
rect 59436 47300 59460 47302
rect 59220 47280 59516 47300
rect 60740 46504 60792 46510
rect 60740 46446 60792 46452
rect 59220 46268 59516 46288
rect 59276 46266 59300 46268
rect 59356 46266 59380 46268
rect 59436 46266 59460 46268
rect 59298 46214 59300 46266
rect 59362 46214 59374 46266
rect 59436 46214 59438 46266
rect 59276 46212 59300 46214
rect 59356 46212 59380 46214
rect 59436 46212 59460 46214
rect 59220 46192 59516 46212
rect 59220 45180 59516 45200
rect 59276 45178 59300 45180
rect 59356 45178 59380 45180
rect 59436 45178 59460 45180
rect 59298 45126 59300 45178
rect 59362 45126 59374 45178
rect 59436 45126 59438 45178
rect 59276 45124 59300 45126
rect 59356 45124 59380 45126
rect 59436 45124 59460 45126
rect 59220 45104 59516 45124
rect 58716 45008 58768 45014
rect 58716 44950 58768 44956
rect 58624 44940 58676 44946
rect 58624 44882 58676 44888
rect 57704 41472 57756 41478
rect 57704 41414 57756 41420
rect 58636 41414 58664 44882
rect 57336 33448 57388 33454
rect 57336 33390 57388 33396
rect 57244 26308 57296 26314
rect 57244 26250 57296 26256
rect 56968 23112 57020 23118
rect 56968 23054 57020 23060
rect 56980 22438 57008 23054
rect 56968 22432 57020 22438
rect 56968 22374 57020 22380
rect 57256 8090 57284 26250
rect 57348 8294 57376 33390
rect 57428 26852 57480 26858
rect 57428 26794 57480 26800
rect 57336 8288 57388 8294
rect 57336 8230 57388 8236
rect 57440 8090 57468 26794
rect 57716 11626 57744 41414
rect 58544 41386 58664 41414
rect 57888 34944 57940 34950
rect 57888 34886 57940 34892
rect 57900 34746 57928 34886
rect 57888 34740 57940 34746
rect 57888 34682 57940 34688
rect 58440 25832 58492 25838
rect 58440 25774 58492 25780
rect 58452 23322 58480 25774
rect 58544 24818 58572 41386
rect 58728 35766 58756 44950
rect 58808 44940 58860 44946
rect 58808 44882 58860 44888
rect 58820 44538 58848 44882
rect 60004 44804 60056 44810
rect 60004 44746 60056 44752
rect 58808 44532 58860 44538
rect 58808 44474 58860 44480
rect 59220 44092 59516 44112
rect 59276 44090 59300 44092
rect 59356 44090 59380 44092
rect 59436 44090 59460 44092
rect 59298 44038 59300 44090
rect 59362 44038 59374 44090
rect 59436 44038 59438 44090
rect 59276 44036 59300 44038
rect 59356 44036 59380 44038
rect 59436 44036 59460 44038
rect 59220 44016 59516 44036
rect 59220 43004 59516 43024
rect 59276 43002 59300 43004
rect 59356 43002 59380 43004
rect 59436 43002 59460 43004
rect 59298 42950 59300 43002
rect 59362 42950 59374 43002
rect 59436 42950 59438 43002
rect 59276 42948 59300 42950
rect 59356 42948 59380 42950
rect 59436 42948 59460 42950
rect 59220 42928 59516 42948
rect 59220 41916 59516 41936
rect 59276 41914 59300 41916
rect 59356 41914 59380 41916
rect 59436 41914 59460 41916
rect 59298 41862 59300 41914
rect 59362 41862 59374 41914
rect 59436 41862 59438 41914
rect 59276 41860 59300 41862
rect 59356 41860 59380 41862
rect 59436 41860 59460 41862
rect 59220 41840 59516 41860
rect 59220 40828 59516 40848
rect 59276 40826 59300 40828
rect 59356 40826 59380 40828
rect 59436 40826 59460 40828
rect 59298 40774 59300 40826
rect 59362 40774 59374 40826
rect 59436 40774 59438 40826
rect 59276 40772 59300 40774
rect 59356 40772 59380 40774
rect 59436 40772 59460 40774
rect 59220 40752 59516 40772
rect 59220 39740 59516 39760
rect 59276 39738 59300 39740
rect 59356 39738 59380 39740
rect 59436 39738 59460 39740
rect 59298 39686 59300 39738
rect 59362 39686 59374 39738
rect 59436 39686 59438 39738
rect 59276 39684 59300 39686
rect 59356 39684 59380 39686
rect 59436 39684 59460 39686
rect 59220 39664 59516 39684
rect 59220 38652 59516 38672
rect 59276 38650 59300 38652
rect 59356 38650 59380 38652
rect 59436 38650 59460 38652
rect 59298 38598 59300 38650
rect 59362 38598 59374 38650
rect 59436 38598 59438 38650
rect 59276 38596 59300 38598
rect 59356 38596 59380 38598
rect 59436 38596 59460 38598
rect 59220 38576 59516 38596
rect 59220 37564 59516 37584
rect 59276 37562 59300 37564
rect 59356 37562 59380 37564
rect 59436 37562 59460 37564
rect 59298 37510 59300 37562
rect 59362 37510 59374 37562
rect 59436 37510 59438 37562
rect 59276 37508 59300 37510
rect 59356 37508 59380 37510
rect 59436 37508 59460 37510
rect 59220 37488 59516 37508
rect 59220 36476 59516 36496
rect 59276 36474 59300 36476
rect 59356 36474 59380 36476
rect 59436 36474 59460 36476
rect 59298 36422 59300 36474
rect 59362 36422 59374 36474
rect 59436 36422 59438 36474
rect 59276 36420 59300 36422
rect 59356 36420 59380 36422
rect 59436 36420 59460 36422
rect 59220 36400 59516 36420
rect 59544 36236 59596 36242
rect 59544 36178 59596 36184
rect 58716 35760 58768 35766
rect 58716 35702 58768 35708
rect 58728 31958 58756 35702
rect 59220 35388 59516 35408
rect 59276 35386 59300 35388
rect 59356 35386 59380 35388
rect 59436 35386 59460 35388
rect 59298 35334 59300 35386
rect 59362 35334 59374 35386
rect 59436 35334 59438 35386
rect 59276 35332 59300 35334
rect 59356 35332 59380 35334
rect 59436 35332 59460 35334
rect 59220 35312 59516 35332
rect 59220 34300 59516 34320
rect 59276 34298 59300 34300
rect 59356 34298 59380 34300
rect 59436 34298 59460 34300
rect 59298 34246 59300 34298
rect 59362 34246 59374 34298
rect 59436 34246 59438 34298
rect 59276 34244 59300 34246
rect 59356 34244 59380 34246
rect 59436 34244 59460 34246
rect 59220 34224 59516 34244
rect 59220 33212 59516 33232
rect 59276 33210 59300 33212
rect 59356 33210 59380 33212
rect 59436 33210 59460 33212
rect 59298 33158 59300 33210
rect 59362 33158 59374 33210
rect 59436 33158 59438 33210
rect 59276 33156 59300 33158
rect 59356 33156 59380 33158
rect 59436 33156 59460 33158
rect 59220 33136 59516 33156
rect 59220 32124 59516 32144
rect 59276 32122 59300 32124
rect 59356 32122 59380 32124
rect 59436 32122 59460 32124
rect 59298 32070 59300 32122
rect 59362 32070 59374 32122
rect 59436 32070 59438 32122
rect 59276 32068 59300 32070
rect 59356 32068 59380 32070
rect 59436 32068 59460 32070
rect 59220 32048 59516 32068
rect 58716 31952 58768 31958
rect 58716 31894 58768 31900
rect 59220 31036 59516 31056
rect 59276 31034 59300 31036
rect 59356 31034 59380 31036
rect 59436 31034 59460 31036
rect 59298 30982 59300 31034
rect 59362 30982 59374 31034
rect 59436 30982 59438 31034
rect 59276 30980 59300 30982
rect 59356 30980 59380 30982
rect 59436 30980 59460 30982
rect 59220 30960 59516 30980
rect 59220 29948 59516 29968
rect 59276 29946 59300 29948
rect 59356 29946 59380 29948
rect 59436 29946 59460 29948
rect 59298 29894 59300 29946
rect 59362 29894 59374 29946
rect 59436 29894 59438 29946
rect 59276 29892 59300 29894
rect 59356 29892 59380 29894
rect 59436 29892 59460 29894
rect 59220 29872 59516 29892
rect 59220 28860 59516 28880
rect 59276 28858 59300 28860
rect 59356 28858 59380 28860
rect 59436 28858 59460 28860
rect 59298 28806 59300 28858
rect 59362 28806 59374 28858
rect 59436 28806 59438 28858
rect 59276 28804 59300 28806
rect 59356 28804 59380 28806
rect 59436 28804 59460 28806
rect 59220 28784 59516 28804
rect 59220 27772 59516 27792
rect 59276 27770 59300 27772
rect 59356 27770 59380 27772
rect 59436 27770 59460 27772
rect 59298 27718 59300 27770
rect 59362 27718 59374 27770
rect 59436 27718 59438 27770
rect 59276 27716 59300 27718
rect 59356 27716 59380 27718
rect 59436 27716 59460 27718
rect 59220 27696 59516 27716
rect 59220 26684 59516 26704
rect 59276 26682 59300 26684
rect 59356 26682 59380 26684
rect 59436 26682 59460 26684
rect 59298 26630 59300 26682
rect 59362 26630 59374 26682
rect 59436 26630 59438 26682
rect 59276 26628 59300 26630
rect 59356 26628 59380 26630
rect 59436 26628 59460 26630
rect 59220 26608 59516 26628
rect 59220 25596 59516 25616
rect 59276 25594 59300 25596
rect 59356 25594 59380 25596
rect 59436 25594 59460 25596
rect 59298 25542 59300 25594
rect 59362 25542 59374 25594
rect 59436 25542 59438 25594
rect 59276 25540 59300 25542
rect 59356 25540 59380 25542
rect 59436 25540 59460 25542
rect 59220 25520 59516 25540
rect 58532 24812 58584 24818
rect 58532 24754 58584 24760
rect 59220 24508 59516 24528
rect 59276 24506 59300 24508
rect 59356 24506 59380 24508
rect 59436 24506 59460 24508
rect 59298 24454 59300 24506
rect 59362 24454 59374 24506
rect 59436 24454 59438 24506
rect 59276 24452 59300 24454
rect 59356 24452 59380 24454
rect 59436 24452 59460 24454
rect 59220 24432 59516 24452
rect 59220 23420 59516 23440
rect 59276 23418 59300 23420
rect 59356 23418 59380 23420
rect 59436 23418 59460 23420
rect 59298 23366 59300 23418
rect 59362 23366 59374 23418
rect 59436 23366 59438 23418
rect 59276 23364 59300 23366
rect 59356 23364 59380 23366
rect 59436 23364 59460 23366
rect 59220 23344 59516 23364
rect 58440 23316 58492 23322
rect 58440 23258 58492 23264
rect 59220 22332 59516 22352
rect 59276 22330 59300 22332
rect 59356 22330 59380 22332
rect 59436 22330 59460 22332
rect 59298 22278 59300 22330
rect 59362 22278 59374 22330
rect 59436 22278 59438 22330
rect 59276 22276 59300 22278
rect 59356 22276 59380 22278
rect 59436 22276 59460 22278
rect 59220 22256 59516 22276
rect 59220 21244 59516 21264
rect 59276 21242 59300 21244
rect 59356 21242 59380 21244
rect 59436 21242 59460 21244
rect 59298 21190 59300 21242
rect 59362 21190 59374 21242
rect 59436 21190 59438 21242
rect 59276 21188 59300 21190
rect 59356 21188 59380 21190
rect 59436 21188 59460 21190
rect 59220 21168 59516 21188
rect 57980 21004 58032 21010
rect 57980 20946 58032 20952
rect 57704 11620 57756 11626
rect 57704 11562 57756 11568
rect 57520 8288 57572 8294
rect 57520 8230 57572 8236
rect 57244 8084 57296 8090
rect 57428 8084 57480 8090
rect 57296 8044 57376 8072
rect 57244 8026 57296 8032
rect 56784 7540 56836 7546
rect 57152 7540 57204 7546
rect 56836 7500 57008 7528
rect 56784 7482 56836 7488
rect 56232 7200 56284 7206
rect 56232 7142 56284 7148
rect 56140 6112 56192 6118
rect 56140 6054 56192 6060
rect 56152 4690 56180 6054
rect 56244 5098 56272 7142
rect 56324 6656 56376 6662
rect 56324 6598 56376 6604
rect 56336 5166 56364 6598
rect 56416 6180 56468 6186
rect 56416 6122 56468 6128
rect 56428 5778 56456 6122
rect 56876 6112 56928 6118
rect 56876 6054 56928 6060
rect 56416 5772 56468 5778
rect 56416 5714 56468 5720
rect 56324 5160 56376 5166
rect 56324 5102 56376 5108
rect 56232 5092 56284 5098
rect 56232 5034 56284 5040
rect 56140 4684 56192 4690
rect 56140 4626 56192 4632
rect 56428 4570 56456 5714
rect 56784 5568 56836 5574
rect 56784 5510 56836 5516
rect 56600 5160 56652 5166
rect 56600 5102 56652 5108
rect 56152 4542 56456 4570
rect 56048 2916 56100 2922
rect 56048 2858 56100 2864
rect 55956 2848 56008 2854
rect 55956 2790 56008 2796
rect 55864 2576 55916 2582
rect 55864 2518 55916 2524
rect 55968 800 55996 2790
rect 56152 800 56180 4542
rect 56232 4480 56284 4486
rect 56232 4422 56284 4428
rect 56244 4282 56272 4422
rect 56232 4276 56284 4282
rect 56232 4218 56284 4224
rect 56324 4140 56376 4146
rect 56324 4082 56376 4088
rect 56232 4004 56284 4010
rect 56232 3946 56284 3952
rect 56244 800 56272 3946
rect 56336 2922 56364 4082
rect 56416 3460 56468 3466
rect 56416 3402 56468 3408
rect 56324 2916 56376 2922
rect 56324 2858 56376 2864
rect 56428 800 56456 3402
rect 56612 2774 56640 5102
rect 56692 4684 56744 4690
rect 56692 4626 56744 4632
rect 56520 2746 56640 2774
rect 56520 800 56548 2746
rect 56704 800 56732 4626
rect 56796 4078 56824 5510
rect 56888 4690 56916 6054
rect 56876 4684 56928 4690
rect 56876 4626 56928 4632
rect 56876 4480 56928 4486
rect 56876 4422 56928 4428
rect 56784 4072 56836 4078
rect 56784 4014 56836 4020
rect 56784 2984 56836 2990
rect 56784 2926 56836 2932
rect 56796 800 56824 2926
rect 56888 1442 56916 4422
rect 56980 2582 57008 7500
rect 57152 7482 57204 7488
rect 57060 4684 57112 4690
rect 57060 4626 57112 4632
rect 56968 2576 57020 2582
rect 56968 2518 57020 2524
rect 56888 1414 57008 1442
rect 56980 800 57008 1414
rect 57072 800 57100 4626
rect 57164 3670 57192 7482
rect 57244 6656 57296 6662
rect 57244 6598 57296 6604
rect 57256 5166 57284 6598
rect 57244 5160 57296 5166
rect 57244 5102 57296 5108
rect 57152 3664 57204 3670
rect 57152 3606 57204 3612
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 57256 800 57284 3402
rect 57348 2922 57376 8044
rect 57428 8026 57480 8032
rect 57440 3670 57468 8026
rect 57532 7546 57560 8230
rect 57992 7546 58020 20946
rect 59220 20156 59516 20176
rect 59276 20154 59300 20156
rect 59356 20154 59380 20156
rect 59436 20154 59460 20156
rect 59298 20102 59300 20154
rect 59362 20102 59374 20154
rect 59436 20102 59438 20154
rect 59276 20100 59300 20102
rect 59356 20100 59380 20102
rect 59436 20100 59460 20102
rect 59220 20080 59516 20100
rect 59220 19068 59516 19088
rect 59276 19066 59300 19068
rect 59356 19066 59380 19068
rect 59436 19066 59460 19068
rect 59298 19014 59300 19066
rect 59362 19014 59374 19066
rect 59436 19014 59438 19066
rect 59276 19012 59300 19014
rect 59356 19012 59380 19014
rect 59436 19012 59460 19014
rect 59220 18992 59516 19012
rect 59220 17980 59516 18000
rect 59276 17978 59300 17980
rect 59356 17978 59380 17980
rect 59436 17978 59460 17980
rect 59298 17926 59300 17978
rect 59362 17926 59374 17978
rect 59436 17926 59438 17978
rect 59276 17924 59300 17926
rect 59356 17924 59380 17926
rect 59436 17924 59460 17926
rect 59220 17904 59516 17924
rect 59220 16892 59516 16912
rect 59276 16890 59300 16892
rect 59356 16890 59380 16892
rect 59436 16890 59460 16892
rect 59298 16838 59300 16890
rect 59362 16838 59374 16890
rect 59436 16838 59438 16890
rect 59276 16836 59300 16838
rect 59356 16836 59380 16838
rect 59436 16836 59460 16838
rect 59220 16816 59516 16836
rect 59556 16574 59584 36178
rect 60016 35834 60044 44746
rect 60188 42628 60240 42634
rect 60188 42570 60240 42576
rect 60004 35828 60056 35834
rect 60004 35770 60056 35776
rect 59556 16546 59676 16574
rect 59220 15804 59516 15824
rect 59276 15802 59300 15804
rect 59356 15802 59380 15804
rect 59436 15802 59460 15804
rect 59298 15750 59300 15802
rect 59362 15750 59374 15802
rect 59436 15750 59438 15802
rect 59276 15748 59300 15750
rect 59356 15748 59380 15750
rect 59436 15748 59460 15750
rect 59220 15728 59516 15748
rect 59220 14716 59516 14736
rect 59276 14714 59300 14716
rect 59356 14714 59380 14716
rect 59436 14714 59460 14716
rect 59298 14662 59300 14714
rect 59362 14662 59374 14714
rect 59436 14662 59438 14714
rect 59276 14660 59300 14662
rect 59356 14660 59380 14662
rect 59436 14660 59460 14662
rect 59220 14640 59516 14660
rect 58440 14272 58492 14278
rect 58440 14214 58492 14220
rect 57520 7540 57572 7546
rect 57520 7482 57572 7488
rect 57980 7540 58032 7546
rect 58032 7500 58204 7528
rect 57980 7482 58032 7488
rect 57612 6724 57664 6730
rect 57612 6666 57664 6672
rect 57520 6112 57572 6118
rect 57520 6054 57572 6060
rect 57532 4690 57560 6054
rect 57624 5166 57652 6666
rect 57888 6656 57940 6662
rect 57888 6598 57940 6604
rect 57704 5568 57756 5574
rect 57704 5510 57756 5516
rect 57612 5160 57664 5166
rect 57612 5102 57664 5108
rect 57520 4684 57572 4690
rect 57520 4626 57572 4632
rect 57428 3664 57480 3670
rect 57428 3606 57480 3612
rect 57336 2916 57388 2922
rect 57336 2858 57388 2864
rect 57624 2774 57652 5102
rect 57716 4078 57744 5510
rect 57900 4690 57928 6598
rect 57888 4684 57940 4690
rect 57888 4626 57940 4632
rect 57900 4486 57928 4626
rect 57888 4480 57940 4486
rect 57888 4422 57940 4428
rect 57704 4072 57756 4078
rect 57704 4014 57756 4020
rect 57980 3596 58032 3602
rect 57980 3538 58032 3544
rect 57796 3528 57848 3534
rect 57796 3470 57848 3476
rect 57348 2746 57652 2774
rect 57348 800 57376 2746
rect 57520 2644 57572 2650
rect 57520 2586 57572 2592
rect 57532 800 57560 2586
rect 57612 2372 57664 2378
rect 57612 2314 57664 2320
rect 57624 800 57652 2314
rect 57808 800 57836 3470
rect 57992 800 58020 3538
rect 58176 2582 58204 7500
rect 58256 4072 58308 4078
rect 58256 4014 58308 4020
rect 58164 2576 58216 2582
rect 58164 2518 58216 2524
rect 58072 2372 58124 2378
rect 58072 2314 58124 2320
rect 58084 800 58112 2314
rect 58268 800 58296 4014
rect 58348 2984 58400 2990
rect 58348 2926 58400 2932
rect 58360 800 58388 2926
rect 58452 2310 58480 14214
rect 59220 13628 59516 13648
rect 59276 13626 59300 13628
rect 59356 13626 59380 13628
rect 59436 13626 59460 13628
rect 59298 13574 59300 13626
rect 59362 13574 59374 13626
rect 59436 13574 59438 13626
rect 59276 13572 59300 13574
rect 59356 13572 59380 13574
rect 59436 13572 59460 13574
rect 59220 13552 59516 13572
rect 59220 12540 59516 12560
rect 59276 12538 59300 12540
rect 59356 12538 59380 12540
rect 59436 12538 59460 12540
rect 59298 12486 59300 12538
rect 59362 12486 59374 12538
rect 59436 12486 59438 12538
rect 59276 12484 59300 12486
rect 59356 12484 59380 12486
rect 59436 12484 59460 12486
rect 59220 12464 59516 12484
rect 59220 11452 59516 11472
rect 59276 11450 59300 11452
rect 59356 11450 59380 11452
rect 59436 11450 59460 11452
rect 59298 11398 59300 11450
rect 59362 11398 59374 11450
rect 59436 11398 59438 11450
rect 59276 11396 59300 11398
rect 59356 11396 59380 11398
rect 59436 11396 59460 11398
rect 59220 11376 59516 11396
rect 59220 10364 59516 10384
rect 59276 10362 59300 10364
rect 59356 10362 59380 10364
rect 59436 10362 59460 10364
rect 59298 10310 59300 10362
rect 59362 10310 59374 10362
rect 59436 10310 59438 10362
rect 59276 10308 59300 10310
rect 59356 10308 59380 10310
rect 59436 10308 59460 10310
rect 59220 10288 59516 10308
rect 59220 9276 59516 9296
rect 59276 9274 59300 9276
rect 59356 9274 59380 9276
rect 59436 9274 59460 9276
rect 59298 9222 59300 9274
rect 59362 9222 59374 9274
rect 59436 9222 59438 9274
rect 59276 9220 59300 9222
rect 59356 9220 59380 9222
rect 59436 9220 59460 9222
rect 59220 9200 59516 9220
rect 59220 8188 59516 8208
rect 59276 8186 59300 8188
rect 59356 8186 59380 8188
rect 59436 8186 59460 8188
rect 59298 8134 59300 8186
rect 59362 8134 59374 8186
rect 59436 8134 59438 8186
rect 59276 8132 59300 8134
rect 59356 8132 59380 8134
rect 59436 8132 59460 8134
rect 59220 8112 59516 8132
rect 59544 7200 59596 7206
rect 59544 7142 59596 7148
rect 59220 7100 59516 7120
rect 59276 7098 59300 7100
rect 59356 7098 59380 7100
rect 59436 7098 59460 7100
rect 59298 7046 59300 7098
rect 59362 7046 59374 7098
rect 59436 7046 59438 7098
rect 59276 7044 59300 7046
rect 59356 7044 59380 7046
rect 59436 7044 59460 7046
rect 59220 7024 59516 7044
rect 58900 6112 58952 6118
rect 58900 6054 58952 6060
rect 58808 5568 58860 5574
rect 58808 5510 58860 5516
rect 58716 5024 58768 5030
rect 58716 4966 58768 4972
rect 58624 4684 58676 4690
rect 58624 4626 58676 4632
rect 58532 3392 58584 3398
rect 58532 3334 58584 3340
rect 58544 2650 58572 3334
rect 58532 2644 58584 2650
rect 58532 2586 58584 2592
rect 58544 2514 58572 2586
rect 58532 2508 58584 2514
rect 58532 2450 58584 2456
rect 58440 2304 58492 2310
rect 58440 2246 58492 2252
rect 58532 2304 58584 2310
rect 58532 2246 58584 2252
rect 58544 800 58572 2246
rect 58636 800 58664 4626
rect 58728 3602 58756 4966
rect 58820 4078 58848 5510
rect 58912 4690 58940 6054
rect 59220 6012 59516 6032
rect 59276 6010 59300 6012
rect 59356 6010 59380 6012
rect 59436 6010 59460 6012
rect 59298 5958 59300 6010
rect 59362 5958 59374 6010
rect 59436 5958 59438 6010
rect 59276 5956 59300 5958
rect 59356 5956 59380 5958
rect 59436 5956 59460 5958
rect 59220 5936 59516 5956
rect 59556 5681 59584 7142
rect 59648 6866 59676 16546
rect 60200 7546 60228 42570
rect 60372 35624 60424 35630
rect 60372 35566 60424 35572
rect 60384 35222 60412 35566
rect 60372 35216 60424 35222
rect 60372 35158 60424 35164
rect 60464 28008 60516 28014
rect 60464 27950 60516 27956
rect 60476 9450 60504 27950
rect 60464 9444 60516 9450
rect 60464 9386 60516 9392
rect 60752 7546 60780 46446
rect 60832 43240 60884 43246
rect 60832 43182 60884 43188
rect 60844 7750 60872 43182
rect 60924 35760 60976 35766
rect 60924 35702 60976 35708
rect 60936 35494 60964 35702
rect 60924 35488 60976 35494
rect 60924 35430 60976 35436
rect 60924 27328 60976 27334
rect 60924 27270 60976 27276
rect 60936 21010 60964 27270
rect 60924 21004 60976 21010
rect 60924 20946 60976 20952
rect 61488 18426 61516 66234
rect 64220 65308 64516 65328
rect 64276 65306 64300 65308
rect 64356 65306 64380 65308
rect 64436 65306 64460 65308
rect 64298 65254 64300 65306
rect 64362 65254 64374 65306
rect 64436 65254 64438 65306
rect 64276 65252 64300 65254
rect 64356 65252 64380 65254
rect 64436 65252 64460 65254
rect 64220 65232 64516 65252
rect 64220 64220 64516 64240
rect 64276 64218 64300 64220
rect 64356 64218 64380 64220
rect 64436 64218 64460 64220
rect 64298 64166 64300 64218
rect 64362 64166 64374 64218
rect 64436 64166 64438 64218
rect 64276 64164 64300 64166
rect 64356 64164 64380 64166
rect 64436 64164 64460 64166
rect 64220 64144 64516 64164
rect 64220 63132 64516 63152
rect 64276 63130 64300 63132
rect 64356 63130 64380 63132
rect 64436 63130 64460 63132
rect 64298 63078 64300 63130
rect 64362 63078 64374 63130
rect 64436 63078 64438 63130
rect 64276 63076 64300 63078
rect 64356 63076 64380 63078
rect 64436 63076 64460 63078
rect 64220 63056 64516 63076
rect 62764 63028 62816 63034
rect 62764 62970 62816 62976
rect 62776 55078 62804 62970
rect 64220 62044 64516 62064
rect 64276 62042 64300 62044
rect 64356 62042 64380 62044
rect 64436 62042 64460 62044
rect 64298 61990 64300 62042
rect 64362 61990 64374 62042
rect 64436 61990 64438 62042
rect 64276 61988 64300 61990
rect 64356 61988 64380 61990
rect 64436 61988 64460 61990
rect 64220 61968 64516 61988
rect 64220 60956 64516 60976
rect 64276 60954 64300 60956
rect 64356 60954 64380 60956
rect 64436 60954 64460 60956
rect 64298 60902 64300 60954
rect 64362 60902 64374 60954
rect 64436 60902 64438 60954
rect 64276 60900 64300 60902
rect 64356 60900 64380 60902
rect 64436 60900 64460 60902
rect 64220 60880 64516 60900
rect 64220 59868 64516 59888
rect 64276 59866 64300 59868
rect 64356 59866 64380 59868
rect 64436 59866 64460 59868
rect 64298 59814 64300 59866
rect 64362 59814 64374 59866
rect 64436 59814 64438 59866
rect 64276 59812 64300 59814
rect 64356 59812 64380 59814
rect 64436 59812 64460 59814
rect 64220 59792 64516 59812
rect 64144 58880 64196 58886
rect 64144 58822 64196 58828
rect 63960 57588 64012 57594
rect 63960 57530 64012 57536
rect 62764 55072 62816 55078
rect 62764 55014 62816 55020
rect 62120 54528 62172 54534
rect 62120 54470 62172 54476
rect 61568 35828 61620 35834
rect 61568 35770 61620 35776
rect 61580 35630 61608 35770
rect 61568 35624 61620 35630
rect 61568 35566 61620 35572
rect 61844 32020 61896 32026
rect 61844 31962 61896 31968
rect 61660 19372 61712 19378
rect 61660 19314 61712 19320
rect 61476 18420 61528 18426
rect 61476 18362 61528 18368
rect 61384 8900 61436 8906
rect 61384 8842 61436 8848
rect 61396 8634 61424 8842
rect 61384 8628 61436 8634
rect 61384 8570 61436 8576
rect 60832 7744 60884 7750
rect 60832 7686 60884 7692
rect 60188 7540 60240 7546
rect 60188 7482 60240 7488
rect 60740 7540 60792 7546
rect 60740 7482 60792 7488
rect 59636 6860 59688 6866
rect 59636 6802 59688 6808
rect 59542 5672 59598 5681
rect 59542 5607 59598 5616
rect 59544 5024 59596 5030
rect 59544 4966 59596 4972
rect 59220 4924 59516 4944
rect 59276 4922 59300 4924
rect 59356 4922 59380 4924
rect 59436 4922 59460 4924
rect 59298 4870 59300 4922
rect 59362 4870 59374 4922
rect 59436 4870 59438 4922
rect 59276 4868 59300 4870
rect 59356 4868 59380 4870
rect 59436 4868 59460 4870
rect 59220 4848 59516 4868
rect 59360 4752 59412 4758
rect 59360 4694 59412 4700
rect 58900 4684 58952 4690
rect 58900 4626 58952 4632
rect 59372 4486 59400 4694
rect 59360 4480 59412 4486
rect 59360 4422 59412 4428
rect 58808 4072 58860 4078
rect 59176 4072 59228 4078
rect 58808 4014 58860 4020
rect 59096 4032 59176 4060
rect 58992 3936 59044 3942
rect 58992 3878 59044 3884
rect 58716 3596 58768 3602
rect 58716 3538 58768 3544
rect 58808 3596 58860 3602
rect 58808 3538 58860 3544
rect 58820 800 58848 3538
rect 59004 2922 59032 3878
rect 58992 2916 59044 2922
rect 58992 2858 59044 2864
rect 58900 2440 58952 2446
rect 58900 2382 58952 2388
rect 58912 800 58940 2382
rect 59004 1358 59032 2858
rect 58992 1352 59044 1358
rect 58992 1294 59044 1300
rect 59096 800 59124 4032
rect 59176 4014 59228 4020
rect 59220 3836 59516 3856
rect 59276 3834 59300 3836
rect 59356 3834 59380 3836
rect 59436 3834 59460 3836
rect 59298 3782 59300 3834
rect 59362 3782 59374 3834
rect 59436 3782 59438 3834
rect 59276 3780 59300 3782
rect 59356 3780 59380 3782
rect 59436 3780 59460 3782
rect 59220 3760 59516 3780
rect 59556 3670 59584 4966
rect 59544 3664 59596 3670
rect 59544 3606 59596 3612
rect 59220 2748 59516 2768
rect 59276 2746 59300 2748
rect 59356 2746 59380 2748
rect 59436 2746 59460 2748
rect 59298 2694 59300 2746
rect 59362 2694 59374 2746
rect 59436 2694 59438 2746
rect 59276 2692 59300 2694
rect 59356 2692 59380 2694
rect 59436 2692 59460 2694
rect 59220 2672 59516 2692
rect 59648 2582 59676 6802
rect 60188 6656 60240 6662
rect 60188 6598 60240 6604
rect 60372 6656 60424 6662
rect 60372 6598 60424 6604
rect 59912 6180 59964 6186
rect 59912 6122 59964 6128
rect 59820 6112 59872 6118
rect 59820 6054 59872 6060
rect 59728 4684 59780 4690
rect 59728 4626 59780 4632
rect 59360 2576 59412 2582
rect 59360 2518 59412 2524
rect 59636 2576 59688 2582
rect 59636 2518 59688 2524
rect 59176 1352 59228 1358
rect 59176 1294 59228 1300
rect 59188 800 59216 1294
rect 59372 800 59400 2518
rect 59740 1442 59768 4626
rect 59832 4078 59860 6054
rect 59924 5166 59952 6122
rect 60096 6112 60148 6118
rect 60096 6054 60148 6060
rect 60004 5568 60056 5574
rect 60004 5510 60056 5516
rect 59912 5160 59964 5166
rect 59912 5102 59964 5108
rect 59820 4072 59872 4078
rect 59820 4014 59872 4020
rect 59820 2916 59872 2922
rect 59820 2858 59872 2864
rect 59556 1414 59768 1442
rect 59556 800 59584 1414
rect 59832 1170 59860 2858
rect 59648 1142 59860 1170
rect 59648 800 59676 1142
rect 59820 1080 59872 1086
rect 59820 1022 59872 1028
rect 59832 800 59860 1022
rect 59924 800 59952 5102
rect 60016 3602 60044 5510
rect 60108 4690 60136 6054
rect 60096 4684 60148 4690
rect 60096 4626 60148 4632
rect 60200 4622 60228 6598
rect 60280 5568 60332 5574
rect 60280 5510 60332 5516
rect 60188 4616 60240 4622
rect 60188 4558 60240 4564
rect 60004 3596 60056 3602
rect 60004 3538 60056 3544
rect 60096 3596 60148 3602
rect 60096 3538 60148 3544
rect 60108 800 60136 3538
rect 60292 2990 60320 5510
rect 60384 5166 60412 6598
rect 60646 5672 60702 5681
rect 60556 5636 60608 5642
rect 60646 5607 60702 5616
rect 60556 5578 60608 5584
rect 60464 5568 60516 5574
rect 60464 5510 60516 5516
rect 60372 5160 60424 5166
rect 60372 5102 60424 5108
rect 60280 2984 60332 2990
rect 60280 2926 60332 2932
rect 60188 2372 60240 2378
rect 60188 2314 60240 2320
rect 60200 800 60228 2314
rect 60384 800 60412 5102
rect 60476 4078 60504 5510
rect 60464 4072 60516 4078
rect 60464 4014 60516 4020
rect 60476 800 60504 4014
rect 60568 3602 60596 5578
rect 60660 4758 60688 5607
rect 60844 5234 60872 7686
rect 61672 7546 61700 19314
rect 61856 12434 61884 31962
rect 61856 12406 61976 12434
rect 61948 7750 61976 12406
rect 62132 11830 62160 54470
rect 62776 53122 62804 55014
rect 62776 53094 62896 53122
rect 62868 53038 62896 53094
rect 62856 53032 62908 53038
rect 62856 52974 62908 52980
rect 62764 52964 62816 52970
rect 62764 52906 62816 52912
rect 62396 52692 62448 52698
rect 62396 52634 62448 52640
rect 62408 43858 62436 52634
rect 62776 49774 62804 52906
rect 62868 52698 62896 52974
rect 62856 52692 62908 52698
rect 62856 52634 62908 52640
rect 62764 49768 62816 49774
rect 62764 49710 62816 49716
rect 63684 46436 63736 46442
rect 63684 46378 63736 46384
rect 62396 43852 62448 43858
rect 62396 43794 62448 43800
rect 62304 41540 62356 41546
rect 62304 41482 62356 41488
rect 62212 37732 62264 37738
rect 62212 37674 62264 37680
rect 62120 11824 62172 11830
rect 62120 11766 62172 11772
rect 62224 8362 62252 37674
rect 62316 8906 62344 41482
rect 62408 32502 62436 43794
rect 63316 38888 63368 38894
rect 63316 38830 63368 38836
rect 62948 33448 63000 33454
rect 62948 33390 63000 33396
rect 62856 33380 62908 33386
rect 62856 33322 62908 33328
rect 62396 32496 62448 32502
rect 62396 32438 62448 32444
rect 62672 26308 62724 26314
rect 62672 26250 62724 26256
rect 62396 23248 62448 23254
rect 62396 23190 62448 23196
rect 62408 12434 62436 23190
rect 62684 21554 62712 26250
rect 62672 21548 62724 21554
rect 62672 21490 62724 21496
rect 62408 12406 62528 12434
rect 62304 8900 62356 8906
rect 62304 8842 62356 8848
rect 62212 8356 62264 8362
rect 62212 8298 62264 8304
rect 61936 7744 61988 7750
rect 61936 7686 61988 7692
rect 61108 7540 61160 7546
rect 61108 7482 61160 7488
rect 61660 7540 61712 7546
rect 61660 7482 61712 7488
rect 61844 7540 61896 7546
rect 61844 7482 61896 7488
rect 60832 5228 60884 5234
rect 60832 5170 60884 5176
rect 60740 5160 60792 5166
rect 60740 5102 60792 5108
rect 60648 4752 60700 4758
rect 60648 4694 60700 4700
rect 60648 4616 60700 4622
rect 60648 4558 60700 4564
rect 60556 3596 60608 3602
rect 60556 3538 60608 3544
rect 60660 2774 60688 4558
rect 60568 2746 60688 2774
rect 60568 2582 60596 2746
rect 60648 2644 60700 2650
rect 60648 2586 60700 2592
rect 60556 2576 60608 2582
rect 60556 2518 60608 2524
rect 60660 800 60688 2586
rect 60752 800 60780 5102
rect 60924 3596 60976 3602
rect 60924 3538 60976 3544
rect 60936 800 60964 3538
rect 61016 2916 61068 2922
rect 61016 2858 61068 2864
rect 61028 800 61056 2858
rect 61120 2582 61148 7482
rect 61200 7472 61252 7478
rect 61200 7414 61252 7420
rect 61212 2990 61240 7414
rect 61384 6656 61436 6662
rect 61384 6598 61436 6604
rect 61396 5166 61424 6598
rect 61660 6112 61712 6118
rect 61660 6054 61712 6060
rect 61384 5160 61436 5166
rect 61384 5102 61436 5108
rect 61292 5092 61344 5098
rect 61292 5034 61344 5040
rect 61200 2984 61252 2990
rect 61200 2926 61252 2932
rect 61304 2774 61332 5034
rect 61672 4078 61700 6054
rect 61752 5568 61804 5574
rect 61752 5510 61804 5516
rect 61384 4072 61436 4078
rect 61384 4014 61436 4020
rect 61660 4072 61712 4078
rect 61660 4014 61712 4020
rect 61212 2746 61332 2774
rect 61108 2576 61160 2582
rect 61108 2518 61160 2524
rect 61212 800 61240 2746
rect 61396 800 61424 4014
rect 61660 3732 61712 3738
rect 61660 3674 61712 3680
rect 61476 2372 61528 2378
rect 61476 2314 61528 2320
rect 61488 1426 61516 2314
rect 61568 2304 61620 2310
rect 61568 2246 61620 2252
rect 61476 1420 61528 1426
rect 61476 1362 61528 1368
rect 61580 1170 61608 2246
rect 61488 1142 61608 1170
rect 61488 800 61516 1142
rect 61672 800 61700 3674
rect 61764 3670 61792 5510
rect 61752 3664 61804 3670
rect 61752 3606 61804 3612
rect 61752 3528 61804 3534
rect 61752 3470 61804 3476
rect 61764 800 61792 3470
rect 61856 2582 61884 7482
rect 61844 2576 61896 2582
rect 61844 2518 61896 2524
rect 61948 2514 61976 7686
rect 62028 6656 62080 6662
rect 62028 6598 62080 6604
rect 62040 5166 62068 6598
rect 62028 5160 62080 5166
rect 62028 5102 62080 5108
rect 62120 5160 62172 5166
rect 62120 5102 62172 5108
rect 62132 2666 62160 5102
rect 62224 2990 62252 8298
rect 62500 7750 62528 12406
rect 62672 9376 62724 9382
rect 62672 9318 62724 9324
rect 62580 8356 62632 8362
rect 62580 8298 62632 8304
rect 62488 7744 62540 7750
rect 62488 7686 62540 7692
rect 62396 7200 62448 7206
rect 62396 7142 62448 7148
rect 62304 6112 62356 6118
rect 62304 6054 62356 6060
rect 62316 3602 62344 6054
rect 62408 4690 62436 7142
rect 62500 7002 62528 7686
rect 62488 6996 62540 7002
rect 62488 6938 62540 6944
rect 62592 5778 62620 8298
rect 62580 5772 62632 5778
rect 62580 5714 62632 5720
rect 62592 4706 62620 5714
rect 62684 4826 62712 9318
rect 62868 8838 62896 33322
rect 62960 13530 62988 33390
rect 62948 13524 63000 13530
rect 62948 13466 63000 13472
rect 63328 9382 63356 38830
rect 63500 24744 63552 24750
rect 63500 24686 63552 24692
rect 63512 17270 63540 24686
rect 63500 17264 63552 17270
rect 63500 17206 63552 17212
rect 63500 16448 63552 16454
rect 63500 16390 63552 16396
rect 63316 9376 63368 9382
rect 63316 9318 63368 9324
rect 63512 8838 63540 16390
rect 63592 9376 63644 9382
rect 63592 9318 63644 9324
rect 62856 8832 62908 8838
rect 62856 8774 62908 8780
rect 63132 8832 63184 8838
rect 63132 8774 63184 8780
rect 63500 8832 63552 8838
rect 63500 8774 63552 8780
rect 63040 7744 63092 7750
rect 63040 7686 63092 7692
rect 62764 7200 62816 7206
rect 62764 7142 62816 7148
rect 62776 5166 62804 7142
rect 62856 6656 62908 6662
rect 62856 6598 62908 6604
rect 62764 5160 62816 5166
rect 62764 5102 62816 5108
rect 62672 4820 62724 4826
rect 62672 4762 62724 4768
rect 62396 4684 62448 4690
rect 62396 4626 62448 4632
rect 62488 4684 62540 4690
rect 62592 4678 62804 4706
rect 62488 4626 62540 4632
rect 62408 3738 62436 4626
rect 62396 3732 62448 3738
rect 62396 3674 62448 3680
rect 62304 3596 62356 3602
rect 62304 3538 62356 3544
rect 62212 2984 62264 2990
rect 62212 2926 62264 2932
rect 62304 2916 62356 2922
rect 62304 2858 62356 2864
rect 62212 2848 62264 2854
rect 62212 2790 62264 2796
rect 62040 2638 62160 2666
rect 61936 2508 61988 2514
rect 61936 2450 61988 2456
rect 61936 1420 61988 1426
rect 61936 1362 61988 1368
rect 61948 800 61976 1362
rect 62040 800 62068 2638
rect 62224 800 62252 2790
rect 62316 800 62344 2858
rect 62500 800 62528 4626
rect 62580 4072 62632 4078
rect 62580 4014 62632 4020
rect 62592 800 62620 4014
rect 62776 3890 62804 4678
rect 62868 4078 62896 6598
rect 63052 5166 63080 7686
rect 63040 5160 63092 5166
rect 62960 5120 63040 5148
rect 62856 4072 62908 4078
rect 62856 4014 62908 4020
rect 62776 3862 62896 3890
rect 62672 3596 62724 3602
rect 62672 3538 62724 3544
rect 62684 2854 62712 3538
rect 62868 3194 62896 3862
rect 62856 3188 62908 3194
rect 62856 3130 62908 3136
rect 62764 3120 62816 3126
rect 62764 3062 62816 3068
rect 62672 2848 62724 2854
rect 62672 2790 62724 2796
rect 62776 800 62804 3062
rect 62960 2774 62988 5120
rect 63040 5102 63092 5108
rect 63040 4072 63092 4078
rect 63040 4014 63092 4020
rect 62868 2746 62988 2774
rect 62868 800 62896 2746
rect 63052 800 63080 4014
rect 63144 2922 63172 8774
rect 63316 7200 63368 7206
rect 63316 7142 63368 7148
rect 63500 7200 63552 7206
rect 63500 7142 63552 7148
rect 63224 6112 63276 6118
rect 63224 6054 63276 6060
rect 63236 3602 63264 6054
rect 63328 4690 63356 7142
rect 63408 6656 63460 6662
rect 63408 6598 63460 6604
rect 63316 4684 63368 4690
rect 63316 4626 63368 4632
rect 63420 4078 63448 6598
rect 63512 5778 63540 7142
rect 63500 5772 63552 5778
rect 63500 5714 63552 5720
rect 63408 4072 63460 4078
rect 63408 4014 63460 4020
rect 63512 3890 63540 5714
rect 63604 5302 63632 9318
rect 63696 9178 63724 46378
rect 63868 16992 63920 16998
rect 63868 16934 63920 16940
rect 63776 10124 63828 10130
rect 63776 10066 63828 10072
rect 63788 9874 63816 10066
rect 63880 10010 63908 16934
rect 63972 10130 64000 57530
rect 64052 29300 64104 29306
rect 64052 29242 64104 29248
rect 63960 10124 64012 10130
rect 63960 10066 64012 10072
rect 63880 9982 64000 10010
rect 63972 9926 64000 9982
rect 63960 9920 64012 9926
rect 63788 9846 63908 9874
rect 63960 9862 64012 9868
rect 63684 9172 63736 9178
rect 63684 9114 63736 9120
rect 63880 8838 63908 9846
rect 63776 8832 63828 8838
rect 63776 8774 63828 8780
rect 63868 8832 63920 8838
rect 63868 8774 63920 8780
rect 63684 6112 63736 6118
rect 63684 6054 63736 6060
rect 63592 5296 63644 5302
rect 63592 5238 63644 5244
rect 63592 5160 63644 5166
rect 63592 5102 63644 5108
rect 63604 4060 63632 5102
rect 63696 4214 63724 6054
rect 63684 4208 63736 4214
rect 63684 4150 63736 4156
rect 63604 4032 63724 4060
rect 63420 3862 63540 3890
rect 63592 3936 63644 3942
rect 63592 3878 63644 3884
rect 63224 3596 63276 3602
rect 63224 3538 63276 3544
rect 63224 3052 63276 3058
rect 63224 2994 63276 3000
rect 63132 2916 63184 2922
rect 63132 2858 63184 2864
rect 63236 800 63264 2994
rect 63420 2774 63448 3862
rect 63604 3754 63632 3878
rect 63328 2746 63448 2774
rect 63512 3726 63632 3754
rect 63328 800 63356 2746
rect 63408 2440 63460 2446
rect 63408 2382 63460 2388
rect 63420 1426 63448 2382
rect 63408 1420 63460 1426
rect 63408 1362 63460 1368
rect 63512 800 63540 3726
rect 63592 2916 63644 2922
rect 63592 2858 63644 2864
rect 63604 800 63632 2858
rect 63696 1442 63724 4032
rect 63788 2582 63816 8774
rect 63868 7744 63920 7750
rect 63868 7686 63920 7692
rect 63880 5166 63908 7686
rect 63868 5160 63920 5166
rect 63868 5102 63920 5108
rect 63868 4684 63920 4690
rect 63868 4626 63920 4632
rect 63776 2576 63828 2582
rect 63776 2518 63828 2524
rect 63696 1414 63816 1442
rect 63788 800 63816 1414
rect 63880 800 63908 4626
rect 63972 3738 64000 9862
rect 64064 9330 64092 29242
rect 64156 10538 64184 58822
rect 64220 58780 64516 58800
rect 64276 58778 64300 58780
rect 64356 58778 64380 58780
rect 64436 58778 64460 58780
rect 64298 58726 64300 58778
rect 64362 58726 64374 58778
rect 64436 58726 64438 58778
rect 64276 58724 64300 58726
rect 64356 58724 64380 58726
rect 64436 58724 64460 58726
rect 64220 58704 64516 58724
rect 64220 57692 64516 57712
rect 64276 57690 64300 57692
rect 64356 57690 64380 57692
rect 64436 57690 64460 57692
rect 64298 57638 64300 57690
rect 64362 57638 64374 57690
rect 64436 57638 64438 57690
rect 64276 57636 64300 57638
rect 64356 57636 64380 57638
rect 64436 57636 64460 57638
rect 64220 57616 64516 57636
rect 64220 56604 64516 56624
rect 64276 56602 64300 56604
rect 64356 56602 64380 56604
rect 64436 56602 64460 56604
rect 64298 56550 64300 56602
rect 64362 56550 64374 56602
rect 64436 56550 64438 56602
rect 64276 56548 64300 56550
rect 64356 56548 64380 56550
rect 64436 56548 64460 56550
rect 64220 56528 64516 56548
rect 64220 55516 64516 55536
rect 64276 55514 64300 55516
rect 64356 55514 64380 55516
rect 64436 55514 64460 55516
rect 64298 55462 64300 55514
rect 64362 55462 64374 55514
rect 64436 55462 64438 55514
rect 64276 55460 64300 55462
rect 64356 55460 64380 55462
rect 64436 55460 64460 55462
rect 64220 55440 64516 55460
rect 64220 54428 64516 54448
rect 64276 54426 64300 54428
rect 64356 54426 64380 54428
rect 64436 54426 64460 54428
rect 64298 54374 64300 54426
rect 64362 54374 64374 54426
rect 64436 54374 64438 54426
rect 64276 54372 64300 54374
rect 64356 54372 64380 54374
rect 64436 54372 64460 54374
rect 64220 54352 64516 54372
rect 64220 53340 64516 53360
rect 64276 53338 64300 53340
rect 64356 53338 64380 53340
rect 64436 53338 64460 53340
rect 64298 53286 64300 53338
rect 64362 53286 64374 53338
rect 64436 53286 64438 53338
rect 64276 53284 64300 53286
rect 64356 53284 64380 53286
rect 64436 53284 64460 53286
rect 64220 53264 64516 53284
rect 64220 52252 64516 52272
rect 64276 52250 64300 52252
rect 64356 52250 64380 52252
rect 64436 52250 64460 52252
rect 64298 52198 64300 52250
rect 64362 52198 64374 52250
rect 64436 52198 64438 52250
rect 64276 52196 64300 52198
rect 64356 52196 64380 52198
rect 64436 52196 64460 52198
rect 64220 52176 64516 52196
rect 64220 51164 64516 51184
rect 64276 51162 64300 51164
rect 64356 51162 64380 51164
rect 64436 51162 64460 51164
rect 64298 51110 64300 51162
rect 64362 51110 64374 51162
rect 64436 51110 64438 51162
rect 64276 51108 64300 51110
rect 64356 51108 64380 51110
rect 64436 51108 64460 51110
rect 64220 51088 64516 51108
rect 64220 50076 64516 50096
rect 64276 50074 64300 50076
rect 64356 50074 64380 50076
rect 64436 50074 64460 50076
rect 64298 50022 64300 50074
rect 64362 50022 64374 50074
rect 64436 50022 64438 50074
rect 64276 50020 64300 50022
rect 64356 50020 64380 50022
rect 64436 50020 64460 50022
rect 64220 50000 64516 50020
rect 64220 48988 64516 49008
rect 64276 48986 64300 48988
rect 64356 48986 64380 48988
rect 64436 48986 64460 48988
rect 64298 48934 64300 48986
rect 64362 48934 64374 48986
rect 64436 48934 64438 48986
rect 64276 48932 64300 48934
rect 64356 48932 64380 48934
rect 64436 48932 64460 48934
rect 64220 48912 64516 48932
rect 64220 47900 64516 47920
rect 64276 47898 64300 47900
rect 64356 47898 64380 47900
rect 64436 47898 64460 47900
rect 64298 47846 64300 47898
rect 64362 47846 64374 47898
rect 64436 47846 64438 47898
rect 64276 47844 64300 47846
rect 64356 47844 64380 47846
rect 64436 47844 64460 47846
rect 64220 47824 64516 47844
rect 64220 46812 64516 46832
rect 64276 46810 64300 46812
rect 64356 46810 64380 46812
rect 64436 46810 64460 46812
rect 64298 46758 64300 46810
rect 64362 46758 64374 46810
rect 64436 46758 64438 46810
rect 64276 46756 64300 46758
rect 64356 46756 64380 46758
rect 64436 46756 64460 46758
rect 64220 46736 64516 46756
rect 64220 45724 64516 45744
rect 64276 45722 64300 45724
rect 64356 45722 64380 45724
rect 64436 45722 64460 45724
rect 64298 45670 64300 45722
rect 64362 45670 64374 45722
rect 64436 45670 64438 45722
rect 64276 45668 64300 45670
rect 64356 45668 64380 45670
rect 64436 45668 64460 45670
rect 64220 45648 64516 45668
rect 64220 44636 64516 44656
rect 64276 44634 64300 44636
rect 64356 44634 64380 44636
rect 64436 44634 64460 44636
rect 64298 44582 64300 44634
rect 64362 44582 64374 44634
rect 64436 44582 64438 44634
rect 64276 44580 64300 44582
rect 64356 44580 64380 44582
rect 64436 44580 64460 44582
rect 64220 44560 64516 44580
rect 64220 43548 64516 43568
rect 64276 43546 64300 43548
rect 64356 43546 64380 43548
rect 64436 43546 64460 43548
rect 64298 43494 64300 43546
rect 64362 43494 64374 43546
rect 64436 43494 64438 43546
rect 64276 43492 64300 43494
rect 64356 43492 64380 43494
rect 64436 43492 64460 43494
rect 64220 43472 64516 43492
rect 64220 42460 64516 42480
rect 64276 42458 64300 42460
rect 64356 42458 64380 42460
rect 64436 42458 64460 42460
rect 64298 42406 64300 42458
rect 64362 42406 64374 42458
rect 64436 42406 64438 42458
rect 64276 42404 64300 42406
rect 64356 42404 64380 42406
rect 64436 42404 64460 42406
rect 64220 42384 64516 42404
rect 64220 41372 64516 41392
rect 64276 41370 64300 41372
rect 64356 41370 64380 41372
rect 64436 41370 64460 41372
rect 64298 41318 64300 41370
rect 64362 41318 64374 41370
rect 64436 41318 64438 41370
rect 64276 41316 64300 41318
rect 64356 41316 64380 41318
rect 64436 41316 64460 41318
rect 64220 41296 64516 41316
rect 64220 40284 64516 40304
rect 64276 40282 64300 40284
rect 64356 40282 64380 40284
rect 64436 40282 64460 40284
rect 64298 40230 64300 40282
rect 64362 40230 64374 40282
rect 64436 40230 64438 40282
rect 64276 40228 64300 40230
rect 64356 40228 64380 40230
rect 64436 40228 64460 40230
rect 64220 40208 64516 40228
rect 64220 39196 64516 39216
rect 64276 39194 64300 39196
rect 64356 39194 64380 39196
rect 64436 39194 64460 39196
rect 64298 39142 64300 39194
rect 64362 39142 64374 39194
rect 64436 39142 64438 39194
rect 64276 39140 64300 39142
rect 64356 39140 64380 39142
rect 64436 39140 64460 39142
rect 64220 39120 64516 39140
rect 64220 38108 64516 38128
rect 64276 38106 64300 38108
rect 64356 38106 64380 38108
rect 64436 38106 64460 38108
rect 64298 38054 64300 38106
rect 64362 38054 64374 38106
rect 64436 38054 64438 38106
rect 64276 38052 64300 38054
rect 64356 38052 64380 38054
rect 64436 38052 64460 38054
rect 64220 38032 64516 38052
rect 64220 37020 64516 37040
rect 64276 37018 64300 37020
rect 64356 37018 64380 37020
rect 64436 37018 64460 37020
rect 64298 36966 64300 37018
rect 64362 36966 64374 37018
rect 64436 36966 64438 37018
rect 64276 36964 64300 36966
rect 64356 36964 64380 36966
rect 64436 36964 64460 36966
rect 64220 36944 64516 36964
rect 64220 35932 64516 35952
rect 64276 35930 64300 35932
rect 64356 35930 64380 35932
rect 64436 35930 64460 35932
rect 64298 35878 64300 35930
rect 64362 35878 64374 35930
rect 64436 35878 64438 35930
rect 64276 35876 64300 35878
rect 64356 35876 64380 35878
rect 64436 35876 64460 35878
rect 64220 35856 64516 35876
rect 64220 34844 64516 34864
rect 64276 34842 64300 34844
rect 64356 34842 64380 34844
rect 64436 34842 64460 34844
rect 64298 34790 64300 34842
rect 64362 34790 64374 34842
rect 64436 34790 64438 34842
rect 64276 34788 64300 34790
rect 64356 34788 64380 34790
rect 64436 34788 64460 34790
rect 64220 34768 64516 34788
rect 64220 33756 64516 33776
rect 64276 33754 64300 33756
rect 64356 33754 64380 33756
rect 64436 33754 64460 33756
rect 64298 33702 64300 33754
rect 64362 33702 64374 33754
rect 64436 33702 64438 33754
rect 64276 33700 64300 33702
rect 64356 33700 64380 33702
rect 64436 33700 64460 33702
rect 64220 33680 64516 33700
rect 64220 32668 64516 32688
rect 64276 32666 64300 32668
rect 64356 32666 64380 32668
rect 64436 32666 64460 32668
rect 64298 32614 64300 32666
rect 64362 32614 64374 32666
rect 64436 32614 64438 32666
rect 64276 32612 64300 32614
rect 64356 32612 64380 32614
rect 64436 32612 64460 32614
rect 64220 32592 64516 32612
rect 64220 31580 64516 31600
rect 64276 31578 64300 31580
rect 64356 31578 64380 31580
rect 64436 31578 64460 31580
rect 64298 31526 64300 31578
rect 64362 31526 64374 31578
rect 64436 31526 64438 31578
rect 64276 31524 64300 31526
rect 64356 31524 64380 31526
rect 64436 31524 64460 31526
rect 64220 31504 64516 31524
rect 64220 30492 64516 30512
rect 64276 30490 64300 30492
rect 64356 30490 64380 30492
rect 64436 30490 64460 30492
rect 64298 30438 64300 30490
rect 64362 30438 64374 30490
rect 64436 30438 64438 30490
rect 64276 30436 64300 30438
rect 64356 30436 64380 30438
rect 64436 30436 64460 30438
rect 64220 30416 64516 30436
rect 64220 29404 64516 29424
rect 64276 29402 64300 29404
rect 64356 29402 64380 29404
rect 64436 29402 64460 29404
rect 64298 29350 64300 29402
rect 64362 29350 64374 29402
rect 64436 29350 64438 29402
rect 64276 29348 64300 29350
rect 64356 29348 64380 29350
rect 64436 29348 64460 29350
rect 64220 29328 64516 29348
rect 64220 28316 64516 28336
rect 64276 28314 64300 28316
rect 64356 28314 64380 28316
rect 64436 28314 64460 28316
rect 64298 28262 64300 28314
rect 64362 28262 64374 28314
rect 64436 28262 64438 28314
rect 64276 28260 64300 28262
rect 64356 28260 64380 28262
rect 64436 28260 64460 28262
rect 64220 28240 64516 28260
rect 64220 27228 64516 27248
rect 64276 27226 64300 27228
rect 64356 27226 64380 27228
rect 64436 27226 64460 27228
rect 64298 27174 64300 27226
rect 64362 27174 64374 27226
rect 64436 27174 64438 27226
rect 64276 27172 64300 27174
rect 64356 27172 64380 27174
rect 64436 27172 64460 27174
rect 64220 27152 64516 27172
rect 64220 26140 64516 26160
rect 64276 26138 64300 26140
rect 64356 26138 64380 26140
rect 64436 26138 64460 26140
rect 64298 26086 64300 26138
rect 64362 26086 64374 26138
rect 64436 26086 64438 26138
rect 64276 26084 64300 26086
rect 64356 26084 64380 26086
rect 64436 26084 64460 26086
rect 64220 26064 64516 26084
rect 64220 25052 64516 25072
rect 64276 25050 64300 25052
rect 64356 25050 64380 25052
rect 64436 25050 64460 25052
rect 64298 24998 64300 25050
rect 64362 24998 64374 25050
rect 64436 24998 64438 25050
rect 64276 24996 64300 24998
rect 64356 24996 64380 24998
rect 64436 24996 64460 24998
rect 64220 24976 64516 24996
rect 64220 23964 64516 23984
rect 64276 23962 64300 23964
rect 64356 23962 64380 23964
rect 64436 23962 64460 23964
rect 64298 23910 64300 23962
rect 64362 23910 64374 23962
rect 64436 23910 64438 23962
rect 64276 23908 64300 23910
rect 64356 23908 64380 23910
rect 64436 23908 64460 23910
rect 64220 23888 64516 23908
rect 64220 22876 64516 22896
rect 64276 22874 64300 22876
rect 64356 22874 64380 22876
rect 64436 22874 64460 22876
rect 64298 22822 64300 22874
rect 64362 22822 64374 22874
rect 64436 22822 64438 22874
rect 64276 22820 64300 22822
rect 64356 22820 64380 22822
rect 64436 22820 64460 22822
rect 64220 22800 64516 22820
rect 64616 22778 64644 66982
rect 64696 66020 64748 66026
rect 64696 65962 64748 65968
rect 64708 64394 64736 65962
rect 64696 64388 64748 64394
rect 64696 64330 64748 64336
rect 64696 62484 64748 62490
rect 64696 62426 64748 62432
rect 64604 22772 64656 22778
rect 64604 22714 64656 22720
rect 64220 21788 64516 21808
rect 64276 21786 64300 21788
rect 64356 21786 64380 21788
rect 64436 21786 64460 21788
rect 64298 21734 64300 21786
rect 64362 21734 64374 21786
rect 64436 21734 64438 21786
rect 64276 21732 64300 21734
rect 64356 21732 64380 21734
rect 64436 21732 64460 21734
rect 64220 21712 64516 21732
rect 64220 20700 64516 20720
rect 64276 20698 64300 20700
rect 64356 20698 64380 20700
rect 64436 20698 64460 20700
rect 64298 20646 64300 20698
rect 64362 20646 64374 20698
rect 64436 20646 64438 20698
rect 64276 20644 64300 20646
rect 64356 20644 64380 20646
rect 64436 20644 64460 20646
rect 64220 20624 64516 20644
rect 64220 19612 64516 19632
rect 64276 19610 64300 19612
rect 64356 19610 64380 19612
rect 64436 19610 64460 19612
rect 64298 19558 64300 19610
rect 64362 19558 64374 19610
rect 64436 19558 64438 19610
rect 64276 19556 64300 19558
rect 64356 19556 64380 19558
rect 64436 19556 64460 19558
rect 64220 19536 64516 19556
rect 64220 18524 64516 18544
rect 64276 18522 64300 18524
rect 64356 18522 64380 18524
rect 64436 18522 64460 18524
rect 64298 18470 64300 18522
rect 64362 18470 64374 18522
rect 64436 18470 64438 18522
rect 64276 18468 64300 18470
rect 64356 18468 64380 18470
rect 64436 18468 64460 18470
rect 64220 18448 64516 18468
rect 64220 17436 64516 17456
rect 64276 17434 64300 17436
rect 64356 17434 64380 17436
rect 64436 17434 64460 17436
rect 64298 17382 64300 17434
rect 64362 17382 64374 17434
rect 64436 17382 64438 17434
rect 64276 17380 64300 17382
rect 64356 17380 64380 17382
rect 64436 17380 64460 17382
rect 64220 17360 64516 17380
rect 64220 16348 64516 16368
rect 64276 16346 64300 16348
rect 64356 16346 64380 16348
rect 64436 16346 64460 16348
rect 64298 16294 64300 16346
rect 64362 16294 64374 16346
rect 64436 16294 64438 16346
rect 64276 16292 64300 16294
rect 64356 16292 64380 16294
rect 64436 16292 64460 16294
rect 64220 16272 64516 16292
rect 64220 15260 64516 15280
rect 64276 15258 64300 15260
rect 64356 15258 64380 15260
rect 64436 15258 64460 15260
rect 64298 15206 64300 15258
rect 64362 15206 64374 15258
rect 64436 15206 64438 15258
rect 64276 15204 64300 15206
rect 64356 15204 64380 15206
rect 64436 15204 64460 15206
rect 64220 15184 64516 15204
rect 64220 14172 64516 14192
rect 64276 14170 64300 14172
rect 64356 14170 64380 14172
rect 64436 14170 64460 14172
rect 64298 14118 64300 14170
rect 64362 14118 64374 14170
rect 64436 14118 64438 14170
rect 64276 14116 64300 14118
rect 64356 14116 64380 14118
rect 64436 14116 64460 14118
rect 64220 14096 64516 14116
rect 64220 13084 64516 13104
rect 64276 13082 64300 13084
rect 64356 13082 64380 13084
rect 64436 13082 64460 13084
rect 64298 13030 64300 13082
rect 64362 13030 64374 13082
rect 64436 13030 64438 13082
rect 64276 13028 64300 13030
rect 64356 13028 64380 13030
rect 64436 13028 64460 13030
rect 64220 13008 64516 13028
rect 64220 11996 64516 12016
rect 64276 11994 64300 11996
rect 64356 11994 64380 11996
rect 64436 11994 64460 11996
rect 64298 11942 64300 11994
rect 64362 11942 64374 11994
rect 64436 11942 64438 11994
rect 64276 11940 64300 11942
rect 64356 11940 64380 11942
rect 64436 11940 64460 11942
rect 64220 11920 64516 11940
rect 64220 10908 64516 10928
rect 64276 10906 64300 10908
rect 64356 10906 64380 10908
rect 64436 10906 64460 10908
rect 64298 10854 64300 10906
rect 64362 10854 64374 10906
rect 64436 10854 64438 10906
rect 64276 10852 64300 10854
rect 64356 10852 64380 10854
rect 64436 10852 64460 10854
rect 64220 10832 64516 10852
rect 64144 10532 64196 10538
rect 64144 10474 64196 10480
rect 64708 10470 64736 62426
rect 64800 39438 64828 67118
rect 67008 66842 67036 67118
rect 67560 66842 67588 67895
rect 66996 66836 67048 66842
rect 66996 66778 67048 66784
rect 67548 66836 67600 66842
rect 67548 66778 67600 66784
rect 66352 66700 66404 66706
rect 66352 66642 66404 66648
rect 65708 66496 65760 66502
rect 65708 66438 65760 66444
rect 66076 66496 66128 66502
rect 66076 66438 66128 66444
rect 65524 66156 65576 66162
rect 65524 66098 65576 66104
rect 65536 65754 65564 66098
rect 65524 65748 65576 65754
rect 65524 65690 65576 65696
rect 65432 65408 65484 65414
rect 65432 65350 65484 65356
rect 65064 62484 65116 62490
rect 65064 62426 65116 62432
rect 65076 58002 65104 62426
rect 65064 57996 65116 58002
rect 65064 57938 65116 57944
rect 65076 57798 65104 57938
rect 65064 57792 65116 57798
rect 65064 57734 65116 57740
rect 65444 55214 65472 65350
rect 65536 58070 65564 65690
rect 65524 58064 65576 58070
rect 65576 58012 65656 58018
rect 65524 58006 65656 58012
rect 65536 57990 65656 58006
rect 65352 55186 65472 55214
rect 65248 53032 65300 53038
rect 65248 52974 65300 52980
rect 64788 39432 64840 39438
rect 64788 39374 64840 39380
rect 65154 33552 65210 33561
rect 65154 33487 65210 33496
rect 64880 32768 64932 32774
rect 64880 32710 64932 32716
rect 64892 16574 64920 32710
rect 65168 32434 65196 33487
rect 65156 32428 65208 32434
rect 65156 32370 65208 32376
rect 64892 16546 65012 16574
rect 64696 10464 64748 10470
rect 64696 10406 64748 10412
rect 64880 10464 64932 10470
rect 64880 10406 64932 10412
rect 64220 9820 64516 9840
rect 64276 9818 64300 9820
rect 64356 9818 64380 9820
rect 64436 9818 64460 9820
rect 64298 9766 64300 9818
rect 64362 9766 64374 9818
rect 64436 9766 64438 9818
rect 64276 9764 64300 9766
rect 64356 9764 64380 9766
rect 64436 9764 64460 9766
rect 64220 9744 64516 9764
rect 64236 9376 64288 9382
rect 64064 9324 64236 9330
rect 64064 9318 64288 9324
rect 64064 9302 64276 9318
rect 64052 8832 64104 8838
rect 64052 8774 64104 8780
rect 64064 6730 64092 8774
rect 64156 6798 64184 9302
rect 64220 8732 64516 8752
rect 64276 8730 64300 8732
rect 64356 8730 64380 8732
rect 64436 8730 64460 8732
rect 64298 8678 64300 8730
rect 64362 8678 64374 8730
rect 64436 8678 64438 8730
rect 64276 8676 64300 8678
rect 64356 8676 64380 8678
rect 64436 8676 64460 8678
rect 64220 8656 64516 8676
rect 64604 8356 64656 8362
rect 64604 8298 64656 8304
rect 64220 7644 64516 7664
rect 64276 7642 64300 7644
rect 64356 7642 64380 7644
rect 64436 7642 64460 7644
rect 64298 7590 64300 7642
rect 64362 7590 64374 7642
rect 64436 7590 64438 7642
rect 64276 7588 64300 7590
rect 64356 7588 64380 7590
rect 64436 7588 64460 7590
rect 64220 7568 64516 7588
rect 64144 6792 64196 6798
rect 64144 6734 64196 6740
rect 64052 6724 64104 6730
rect 64052 6666 64104 6672
rect 64144 6656 64196 6662
rect 64144 6598 64196 6604
rect 64052 5772 64104 5778
rect 64052 5714 64104 5720
rect 64064 4570 64092 5714
rect 64156 4690 64184 6598
rect 64220 6556 64516 6576
rect 64276 6554 64300 6556
rect 64356 6554 64380 6556
rect 64436 6554 64460 6556
rect 64298 6502 64300 6554
rect 64362 6502 64374 6554
rect 64436 6502 64438 6554
rect 64276 6500 64300 6502
rect 64356 6500 64380 6502
rect 64436 6500 64460 6502
rect 64220 6480 64516 6500
rect 64512 6112 64564 6118
rect 64512 6054 64564 6060
rect 64524 5642 64552 6054
rect 64616 5778 64644 8298
rect 64696 8288 64748 8294
rect 64696 8230 64748 8236
rect 64708 6254 64736 8230
rect 64788 7200 64840 7206
rect 64788 7142 64840 7148
rect 64696 6248 64748 6254
rect 64696 6190 64748 6196
rect 64604 5772 64656 5778
rect 64604 5714 64656 5720
rect 64708 5658 64736 6190
rect 64512 5636 64564 5642
rect 64512 5578 64564 5584
rect 64616 5630 64736 5658
rect 64220 5468 64516 5488
rect 64276 5466 64300 5468
rect 64356 5466 64380 5468
rect 64436 5466 64460 5468
rect 64298 5414 64300 5466
rect 64362 5414 64374 5466
rect 64436 5414 64438 5466
rect 64276 5412 64300 5414
rect 64356 5412 64380 5414
rect 64436 5412 64460 5414
rect 64220 5392 64516 5412
rect 64236 5296 64288 5302
rect 64236 5238 64288 5244
rect 64144 4684 64196 4690
rect 64144 4626 64196 4632
rect 64064 4542 64184 4570
rect 64248 4554 64276 5238
rect 64052 4480 64104 4486
rect 64052 4422 64104 4428
rect 63960 3732 64012 3738
rect 63960 3674 64012 3680
rect 64064 3584 64092 4422
rect 63972 3556 64092 3584
rect 63972 2990 64000 3556
rect 64052 3460 64104 3466
rect 64052 3402 64104 3408
rect 63960 2984 64012 2990
rect 63960 2926 64012 2932
rect 64064 800 64092 3402
rect 64156 800 64184 4542
rect 64236 4548 64288 4554
rect 64236 4490 64288 4496
rect 64220 4380 64516 4400
rect 64276 4378 64300 4380
rect 64356 4378 64380 4380
rect 64436 4378 64460 4380
rect 64298 4326 64300 4378
rect 64362 4326 64374 4378
rect 64436 4326 64438 4378
rect 64276 4324 64300 4326
rect 64356 4324 64380 4326
rect 64436 4324 64460 4326
rect 64220 4304 64516 4324
rect 64220 3292 64516 3312
rect 64276 3290 64300 3292
rect 64356 3290 64380 3292
rect 64436 3290 64460 3292
rect 64298 3238 64300 3290
rect 64362 3238 64374 3290
rect 64436 3238 64438 3290
rect 64276 3236 64300 3238
rect 64356 3236 64380 3238
rect 64436 3236 64460 3238
rect 64220 3216 64516 3236
rect 64220 2204 64516 2224
rect 64276 2202 64300 2204
rect 64356 2202 64380 2204
rect 64436 2202 64460 2204
rect 64298 2150 64300 2202
rect 64362 2150 64374 2202
rect 64436 2150 64438 2202
rect 64276 2148 64300 2150
rect 64356 2148 64380 2150
rect 64436 2148 64460 2150
rect 64220 2128 64516 2148
rect 64326 2000 64382 2009
rect 64616 1986 64644 5630
rect 64696 5568 64748 5574
rect 64696 5510 64748 5516
rect 64708 4690 64736 5510
rect 64800 4690 64828 7142
rect 64696 4684 64748 4690
rect 64696 4626 64748 4632
rect 64788 4684 64840 4690
rect 64788 4626 64840 4632
rect 64708 4593 64736 4626
rect 64694 4584 64750 4593
rect 64694 4519 64750 4528
rect 64696 2916 64748 2922
rect 64696 2858 64748 2864
rect 64326 1935 64382 1944
rect 64524 1958 64644 1986
rect 64340 800 64368 1935
rect 64420 1284 64472 1290
rect 64420 1226 64472 1232
rect 64432 800 64460 1226
rect 64524 898 64552 1958
rect 64708 1290 64736 2858
rect 64696 1284 64748 1290
rect 64696 1226 64748 1232
rect 64524 870 64644 898
rect 64616 800 64644 870
rect 64800 800 64828 4626
rect 64892 3670 64920 10406
rect 64984 10198 65012 16546
rect 65260 12782 65288 52974
rect 65352 47598 65380 55186
rect 65432 49972 65484 49978
rect 65432 49914 65484 49920
rect 65340 47592 65392 47598
rect 65340 47534 65392 47540
rect 65340 41064 65392 41070
rect 65340 41006 65392 41012
rect 65352 14278 65380 41006
rect 65340 14272 65392 14278
rect 65340 14214 65392 14220
rect 65248 12776 65300 12782
rect 65248 12718 65300 12724
rect 65064 11824 65116 11830
rect 65064 11766 65116 11772
rect 64972 10192 65024 10198
rect 64972 10134 65024 10140
rect 65076 10010 65104 11766
rect 65444 11150 65472 49914
rect 65628 45490 65656 57990
rect 65616 45484 65668 45490
rect 65616 45426 65668 45432
rect 65524 42152 65576 42158
rect 65524 42094 65576 42100
rect 65432 11144 65484 11150
rect 65432 11086 65484 11092
rect 65536 10470 65564 42094
rect 65720 40730 65748 66438
rect 66088 66094 66116 66438
rect 65800 66088 65852 66094
rect 65800 66030 65852 66036
rect 66076 66088 66128 66094
rect 66076 66030 66128 66036
rect 65812 49094 65840 66030
rect 66168 65408 66220 65414
rect 66168 65350 66220 65356
rect 66180 65074 66208 65350
rect 66168 65068 66220 65074
rect 66168 65010 66220 65016
rect 66260 64932 66312 64938
rect 66260 64874 66312 64880
rect 66168 64320 66220 64326
rect 66168 64262 66220 64268
rect 66180 57254 66208 64262
rect 66272 59634 66300 64874
rect 66260 59628 66312 59634
rect 66260 59570 66312 59576
rect 66168 57248 66220 57254
rect 66168 57190 66220 57196
rect 66364 53106 66392 66642
rect 68098 66600 68154 66609
rect 68098 66535 68154 66544
rect 68112 66094 68140 66535
rect 68100 66088 68152 66094
rect 68100 66030 68152 66036
rect 66720 65952 66772 65958
rect 66720 65894 66772 65900
rect 66732 65618 66760 65894
rect 68112 65754 68140 66030
rect 68100 65748 68152 65754
rect 68100 65690 68152 65696
rect 66720 65612 66772 65618
rect 66720 65554 66772 65560
rect 67640 65544 67692 65550
rect 67640 65486 67692 65492
rect 67180 65136 67232 65142
rect 67180 65078 67232 65084
rect 66812 65000 66864 65006
rect 66812 64942 66864 64948
rect 66628 63232 66680 63238
rect 66628 63174 66680 63180
rect 66536 62688 66588 62694
rect 66536 62630 66588 62636
rect 66548 62422 66576 62630
rect 66536 62416 66588 62422
rect 66536 62358 66588 62364
rect 66640 62234 66668 63174
rect 66548 62206 66668 62234
rect 66352 53100 66404 53106
rect 66352 53042 66404 53048
rect 65984 52420 66036 52426
rect 65984 52362 66036 52368
rect 65800 49088 65852 49094
rect 65800 49030 65852 49036
rect 65708 40724 65760 40730
rect 65708 40666 65760 40672
rect 65892 35216 65944 35222
rect 65892 35158 65944 35164
rect 65800 17332 65852 17338
rect 65800 17274 65852 17280
rect 65524 10464 65576 10470
rect 65524 10406 65576 10412
rect 65708 10464 65760 10470
rect 65708 10406 65760 10412
rect 64984 9982 65104 10010
rect 64984 9926 65012 9982
rect 64972 9920 65024 9926
rect 64972 9862 65024 9868
rect 64880 3664 64932 3670
rect 64880 3606 64932 3612
rect 64880 3460 64932 3466
rect 64880 3402 64932 3408
rect 64892 800 64920 3402
rect 64984 2990 65012 9862
rect 65248 9376 65300 9382
rect 65248 9318 65300 9324
rect 65064 8832 65116 8838
rect 65064 8774 65116 8780
rect 65076 6254 65104 8774
rect 65156 7744 65208 7750
rect 65156 7686 65208 7692
rect 65064 6248 65116 6254
rect 65064 6190 65116 6196
rect 64972 2984 65024 2990
rect 64972 2926 65024 2932
rect 65076 800 65104 6190
rect 65168 5166 65196 7686
rect 65260 7410 65288 9318
rect 65524 8900 65576 8906
rect 65524 8842 65576 8848
rect 65432 8832 65484 8838
rect 65432 8774 65484 8780
rect 65340 7812 65392 7818
rect 65340 7754 65392 7760
rect 65248 7404 65300 7410
rect 65248 7346 65300 7352
rect 65352 6934 65380 7754
rect 65340 6928 65392 6934
rect 65246 6896 65302 6905
rect 65340 6870 65392 6876
rect 65444 6866 65472 8774
rect 65246 6831 65302 6840
rect 65432 6860 65484 6866
rect 65260 6225 65288 6831
rect 65432 6802 65484 6808
rect 65340 6792 65392 6798
rect 65340 6734 65392 6740
rect 65246 6216 65302 6225
rect 65246 6151 65302 6160
rect 65156 5160 65208 5166
rect 65156 5102 65208 5108
rect 65260 4842 65288 6151
rect 65168 4814 65288 4842
rect 65168 3913 65196 4814
rect 65248 4684 65300 4690
rect 65248 4626 65300 4632
rect 65154 3904 65210 3913
rect 65154 3839 65210 3848
rect 65260 3754 65288 4626
rect 65168 3726 65288 3754
rect 65168 2514 65196 3726
rect 65352 3618 65380 6734
rect 65260 3590 65380 3618
rect 65260 2582 65288 3590
rect 65340 2916 65392 2922
rect 65340 2858 65392 2864
rect 65248 2576 65300 2582
rect 65248 2518 65300 2524
rect 65156 2508 65208 2514
rect 65156 2450 65208 2456
rect 65168 800 65196 2450
rect 65352 800 65380 2858
rect 65444 800 65472 6802
rect 65536 3670 65564 8842
rect 65616 8356 65668 8362
rect 65616 8298 65668 8304
rect 65628 5710 65656 8298
rect 65616 5704 65668 5710
rect 65616 5646 65668 5652
rect 65616 5160 65668 5166
rect 65616 5102 65668 5108
rect 65524 3664 65576 3670
rect 65524 3606 65576 3612
rect 65522 3496 65578 3505
rect 65522 3431 65578 3440
rect 65536 2582 65564 3431
rect 65524 2576 65576 2582
rect 65524 2518 65576 2524
rect 65628 800 65656 5102
rect 65720 2990 65748 10406
rect 65812 9994 65840 17274
rect 65904 11082 65932 35158
rect 65996 11558 66024 52362
rect 66444 51332 66496 51338
rect 66444 51274 66496 51280
rect 66352 32292 66404 32298
rect 66352 32234 66404 32240
rect 66364 28558 66392 32234
rect 66352 28552 66404 28558
rect 66352 28494 66404 28500
rect 66166 28384 66222 28393
rect 66166 28319 66222 28328
rect 66180 27674 66208 28319
rect 66168 27668 66220 27674
rect 66168 27610 66220 27616
rect 66076 18692 66128 18698
rect 66076 18634 66128 18640
rect 66088 16574 66116 18634
rect 66088 16546 66208 16574
rect 65984 11552 66036 11558
rect 65984 11494 66036 11500
rect 65892 11076 65944 11082
rect 65892 11018 65944 11024
rect 66076 11076 66128 11082
rect 66076 11018 66128 11024
rect 65800 9988 65852 9994
rect 65800 9930 65852 9936
rect 65892 9920 65944 9926
rect 65892 9862 65944 9868
rect 65904 7834 65932 9862
rect 65984 9376 66036 9382
rect 65984 9318 66036 9324
rect 65812 7806 65932 7834
rect 65812 6905 65840 7806
rect 65892 7744 65944 7750
rect 65892 7686 65944 7692
rect 65798 6896 65854 6905
rect 65798 6831 65854 6840
rect 65800 6724 65852 6730
rect 65800 6666 65852 6672
rect 65812 3466 65840 6666
rect 65904 5166 65932 7686
rect 65996 7342 66024 9318
rect 65984 7336 66036 7342
rect 65984 7278 66036 7284
rect 65892 5160 65944 5166
rect 65892 5102 65944 5108
rect 65996 4978 66024 7278
rect 65904 4950 66024 4978
rect 65800 3460 65852 3466
rect 65800 3402 65852 3408
rect 65800 3120 65852 3126
rect 65800 3062 65852 3068
rect 65708 2984 65760 2990
rect 65708 2926 65760 2932
rect 65708 2848 65760 2854
rect 65708 2790 65760 2796
rect 65720 800 65748 2790
rect 65812 2582 65840 3062
rect 65800 2576 65852 2582
rect 65800 2518 65852 2524
rect 65904 800 65932 4950
rect 66088 4078 66116 11018
rect 66180 10538 66208 16546
rect 66456 14074 66484 51274
rect 66548 45082 66576 62206
rect 66824 60042 66852 64942
rect 66904 62824 66956 62830
rect 66904 62766 66956 62772
rect 66916 62490 66944 62766
rect 66904 62484 66956 62490
rect 66904 62426 66956 62432
rect 66812 60036 66864 60042
rect 66812 59978 66864 59984
rect 66720 59560 66772 59566
rect 66720 59502 66772 59508
rect 66628 59016 66680 59022
rect 66628 58958 66680 58964
rect 66536 45076 66588 45082
rect 66536 45018 66588 45024
rect 66640 17882 66668 58958
rect 66732 42770 66760 59502
rect 66996 58336 67048 58342
rect 66996 58278 67048 58284
rect 66904 54120 66956 54126
rect 66904 54062 66956 54068
rect 66812 48204 66864 48210
rect 66812 48146 66864 48152
rect 66720 42764 66772 42770
rect 66720 42706 66772 42712
rect 66824 34746 66852 48146
rect 66916 41818 66944 54062
rect 66904 41812 66956 41818
rect 66904 41754 66956 41760
rect 67008 39370 67036 58278
rect 67088 55276 67140 55282
rect 67088 55218 67140 55224
rect 66996 39364 67048 39370
rect 66996 39306 67048 39312
rect 66904 37732 66956 37738
rect 66904 37674 66956 37680
rect 66812 34740 66864 34746
rect 66812 34682 66864 34688
rect 66916 25498 66944 37674
rect 66996 36236 67048 36242
rect 66996 36178 67048 36184
rect 66904 25492 66956 25498
rect 66904 25434 66956 25440
rect 66720 23792 66772 23798
rect 66720 23734 66772 23740
rect 66628 17876 66680 17882
rect 66628 17818 66680 17824
rect 66444 14068 66496 14074
rect 66444 14010 66496 14016
rect 66732 12434 66760 23734
rect 67008 16046 67036 36178
rect 67100 21418 67128 55218
rect 67192 52154 67220 65078
rect 67652 64954 67680 65486
rect 67652 64926 67772 64954
rect 67640 64864 67692 64870
rect 67640 64806 67692 64812
rect 67652 64326 67680 64806
rect 67640 64320 67692 64326
rect 67640 64262 67692 64268
rect 67272 63776 67324 63782
rect 67272 63718 67324 63724
rect 67284 61878 67312 63718
rect 67272 61872 67324 61878
rect 67272 61814 67324 61820
rect 67272 61736 67324 61742
rect 67272 61678 67324 61684
rect 67284 57594 67312 61678
rect 67364 58404 67416 58410
rect 67364 58346 67416 58352
rect 67272 57588 67324 57594
rect 67272 57530 67324 57536
rect 67284 57390 67312 57530
rect 67272 57384 67324 57390
rect 67272 57326 67324 57332
rect 67180 52148 67232 52154
rect 67180 52090 67232 52096
rect 67180 46980 67232 46986
rect 67180 46922 67232 46928
rect 67192 33522 67220 46922
rect 67272 34672 67324 34678
rect 67272 34614 67324 34620
rect 67180 33516 67232 33522
rect 67180 33458 67232 33464
rect 67284 27130 67312 34614
rect 67272 27124 67324 27130
rect 67272 27066 67324 27072
rect 67284 26926 67312 27066
rect 67180 26920 67232 26926
rect 67180 26862 67232 26868
rect 67272 26920 67324 26926
rect 67272 26862 67324 26868
rect 67192 26234 67220 26862
rect 67192 26206 67312 26234
rect 67284 21690 67312 26206
rect 67376 23322 67404 58346
rect 67456 55344 67508 55350
rect 67456 55286 67508 55292
rect 67468 26042 67496 55286
rect 67548 43648 67600 43654
rect 67548 43590 67600 43596
rect 67560 30870 67588 43590
rect 67548 30864 67600 30870
rect 67548 30806 67600 30812
rect 67456 26036 67508 26042
rect 67456 25978 67508 25984
rect 67468 25838 67496 25978
rect 67456 25832 67508 25838
rect 67456 25774 67508 25780
rect 67364 23316 67416 23322
rect 67364 23258 67416 23264
rect 67272 21684 67324 21690
rect 67272 21626 67324 21632
rect 67284 21486 67312 21626
rect 67272 21480 67324 21486
rect 67272 21422 67324 21428
rect 67088 21412 67140 21418
rect 67088 21354 67140 21360
rect 67088 20392 67140 20398
rect 67088 20334 67140 20340
rect 66996 16040 67048 16046
rect 66996 15982 67048 15988
rect 66732 12406 66852 12434
rect 66352 11552 66404 11558
rect 66352 11494 66404 11500
rect 66628 11552 66680 11558
rect 66628 11494 66680 11500
rect 66168 10532 66220 10538
rect 66168 10474 66220 10480
rect 66168 7812 66220 7818
rect 66168 7754 66220 7760
rect 66180 5778 66208 7754
rect 66260 7336 66312 7342
rect 66260 7278 66312 7284
rect 66168 5772 66220 5778
rect 66168 5714 66220 5720
rect 66180 4146 66208 5714
rect 66168 4140 66220 4146
rect 66168 4082 66220 4088
rect 66076 4072 66128 4078
rect 66076 4014 66128 4020
rect 65984 3936 66036 3942
rect 66036 3884 66116 3890
rect 65984 3878 66116 3884
rect 65996 3862 66116 3878
rect 65984 3732 66036 3738
rect 65984 3674 66036 3680
rect 65996 800 66024 3674
rect 66088 3194 66116 3862
rect 66168 3392 66220 3398
rect 66168 3334 66220 3340
rect 66076 3188 66128 3194
rect 66076 3130 66128 3136
rect 2870 640 2926 649
rect 2870 575 2926 584
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 65982 0 66038 800
rect 66088 649 66116 3130
rect 66180 800 66208 3334
rect 66272 800 66300 7278
rect 66364 5098 66392 11494
rect 66536 11144 66588 11150
rect 66536 11086 66588 11092
rect 66444 8356 66496 8362
rect 66444 8298 66496 8304
rect 66456 6254 66484 8298
rect 66444 6248 66496 6254
rect 66444 6190 66496 6196
rect 66352 5092 66404 5098
rect 66352 5034 66404 5040
rect 66352 3460 66404 3466
rect 66352 3402 66404 3408
rect 66364 2650 66392 3402
rect 66352 2644 66404 2650
rect 66352 2586 66404 2592
rect 66456 800 66484 6190
rect 66548 5846 66576 11086
rect 66640 7886 66668 11494
rect 66824 11082 66852 12406
rect 67100 11558 67128 20334
rect 67744 15706 67772 64926
rect 67824 64932 67876 64938
rect 67824 64874 67876 64880
rect 67836 35018 67864 64874
rect 68098 64016 68154 64025
rect 68098 63951 68100 63960
rect 68152 63951 68154 63960
rect 68100 63922 68152 63928
rect 68100 63300 68152 63306
rect 68100 63242 68152 63248
rect 68112 62665 68140 63242
rect 68098 62656 68154 62665
rect 68098 62591 68154 62600
rect 68098 61296 68154 61305
rect 68098 61231 68100 61240
rect 68152 61231 68154 61240
rect 68100 61202 68152 61208
rect 68098 58712 68154 58721
rect 68098 58647 68154 58656
rect 68112 58614 68140 58647
rect 68100 58608 68152 58614
rect 68100 58550 68152 58556
rect 68098 57352 68154 57361
rect 68098 57287 68100 57296
rect 68152 57287 68154 57296
rect 68100 57258 68152 57264
rect 68100 56296 68152 56302
rect 68100 56238 68152 56244
rect 68112 56137 68140 56238
rect 68098 56128 68154 56137
rect 68098 56063 68154 56072
rect 68100 53508 68152 53514
rect 68100 53450 68152 53456
rect 68112 53417 68140 53450
rect 68098 53408 68154 53417
rect 68098 53343 68154 53352
rect 68098 52048 68154 52057
rect 68098 51983 68100 51992
rect 68152 51983 68154 51992
rect 68100 51954 68152 51960
rect 68100 50856 68152 50862
rect 68098 50824 68100 50833
rect 68152 50824 68154 50833
rect 68098 50759 68154 50768
rect 68098 48104 68154 48113
rect 68098 48039 68100 48048
rect 68152 48039 68154 48048
rect 68100 48010 68152 48016
rect 68100 46980 68152 46986
rect 68100 46922 68152 46928
rect 68112 46889 68140 46922
rect 68098 46880 68154 46889
rect 68098 46815 68154 46824
rect 68098 45520 68154 45529
rect 68098 45455 68154 45464
rect 68112 45422 68140 45455
rect 68100 45416 68152 45422
rect 68100 45358 68152 45364
rect 68098 42800 68154 42809
rect 68098 42735 68100 42744
rect 68152 42735 68154 42744
rect 68100 42706 68152 42712
rect 68098 41576 68154 41585
rect 68098 41511 68100 41520
rect 68152 41511 68154 41520
rect 68100 41482 68152 41488
rect 68098 40216 68154 40225
rect 68098 40151 68154 40160
rect 68112 39982 68140 40151
rect 68100 39976 68152 39982
rect 68100 39918 68152 39924
rect 68100 37732 68152 37738
rect 68100 37674 68152 37680
rect 68112 37641 68140 37674
rect 68098 37632 68154 37641
rect 68098 37567 68154 37576
rect 68098 36272 68154 36281
rect 68098 36207 68100 36216
rect 68152 36207 68154 36216
rect 68100 36178 68152 36184
rect 67916 35692 67968 35698
rect 67916 35634 67968 35640
rect 67928 35154 67956 35634
rect 67916 35148 67968 35154
rect 67916 35090 67968 35096
rect 67824 35012 67876 35018
rect 67824 34954 67876 34960
rect 68928 34944 68980 34950
rect 68926 34912 68928 34921
rect 68980 34912 68982 34921
rect 68926 34847 68982 34856
rect 68098 32328 68154 32337
rect 68098 32263 68100 32272
rect 68152 32263 68154 32272
rect 68100 32234 68152 32240
rect 68098 30968 68154 30977
rect 68098 30903 68154 30912
rect 68112 30870 68140 30903
rect 68100 30864 68152 30870
rect 68100 30806 68152 30812
rect 68100 29708 68152 29714
rect 68100 29650 68152 29656
rect 68112 29617 68140 29650
rect 68098 29608 68154 29617
rect 68098 29543 68154 29552
rect 68098 27024 68154 27033
rect 68098 26959 68100 26968
rect 68152 26959 68154 26968
rect 68100 26930 68152 26936
rect 68100 25764 68152 25770
rect 68100 25706 68152 25712
rect 68112 25673 68140 25706
rect 68098 25664 68154 25673
rect 68098 25599 68154 25608
rect 68100 24744 68152 24750
rect 68100 24686 68152 24692
rect 68112 24313 68140 24686
rect 68098 24304 68154 24313
rect 68098 24239 68154 24248
rect 68098 23080 68154 23089
rect 68098 23015 68100 23024
rect 68152 23015 68154 23024
rect 68100 22986 68152 22992
rect 68098 21720 68154 21729
rect 68098 21655 68154 21664
rect 68112 21622 68140 21655
rect 68100 21616 68152 21622
rect 68100 21558 68152 21564
rect 68100 20392 68152 20398
rect 68098 20360 68100 20369
rect 68152 20360 68154 20369
rect 68098 20295 68154 20304
rect 68100 19236 68152 19242
rect 68100 19178 68152 19184
rect 68112 19145 68140 19178
rect 68098 19136 68154 19145
rect 68098 19071 68154 19080
rect 68098 17776 68154 17785
rect 68098 17711 68100 17720
rect 68152 17711 68154 17720
rect 68100 17682 68152 17688
rect 68100 16652 68152 16658
rect 68100 16594 68152 16600
rect 68112 16425 68140 16594
rect 68098 16416 68154 16425
rect 68098 16351 68154 16360
rect 67732 15700 67784 15706
rect 67732 15642 67784 15648
rect 67744 14958 67772 15642
rect 68098 15056 68154 15065
rect 68098 14991 68100 15000
rect 68152 14991 68154 15000
rect 68100 14962 68152 14968
rect 67180 14952 67232 14958
rect 67180 14894 67232 14900
rect 67732 14952 67784 14958
rect 67732 14894 67784 14900
rect 67192 11694 67220 14894
rect 67272 14476 67324 14482
rect 67272 14418 67324 14424
rect 67180 11688 67232 11694
rect 67180 11630 67232 11636
rect 67088 11552 67140 11558
rect 67088 11494 67140 11500
rect 67284 11354 67312 14418
rect 67640 14272 67692 14278
rect 67640 14214 67692 14220
rect 67652 12434 67680 14214
rect 68100 13864 68152 13870
rect 68098 13832 68100 13841
rect 68152 13832 68154 13841
rect 68098 13767 68154 13776
rect 68098 12472 68154 12481
rect 67652 12406 67956 12434
rect 68098 12407 68154 12416
rect 67364 11552 67416 11558
rect 67364 11494 67416 11500
rect 67640 11552 67692 11558
rect 67640 11494 67692 11500
rect 67272 11348 67324 11354
rect 67272 11290 67324 11296
rect 66812 11076 66864 11082
rect 66812 11018 66864 11024
rect 66720 9376 66772 9382
rect 66720 9318 66772 9324
rect 66628 7880 66680 7886
rect 66628 7822 66680 7828
rect 66628 7744 66680 7750
rect 66628 7686 66680 7692
rect 66536 5840 66588 5846
rect 66536 5782 66588 5788
rect 66640 5166 66668 7686
rect 66732 7342 66760 9318
rect 66720 7336 66772 7342
rect 66720 7278 66772 7284
rect 66720 7200 66772 7206
rect 66720 7142 66772 7148
rect 66628 5160 66680 5166
rect 66548 5120 66628 5148
rect 66548 3738 66576 5120
rect 66628 5102 66680 5108
rect 66628 4004 66680 4010
rect 66628 3946 66680 3952
rect 66536 3732 66588 3738
rect 66536 3674 66588 3680
rect 66640 800 66668 3946
rect 66732 800 66760 7142
rect 66824 3670 66852 11018
rect 67180 10464 67232 10470
rect 67180 10406 67232 10412
rect 66904 9988 66956 9994
rect 66904 9930 66956 9936
rect 66916 7154 66944 9930
rect 66996 9920 67048 9926
rect 66996 9862 67048 9868
rect 67008 7274 67036 9862
rect 67088 8424 67140 8430
rect 67088 8366 67140 8372
rect 66996 7268 67048 7274
rect 66996 7210 67048 7216
rect 66916 7126 67036 7154
rect 66904 6248 66956 6254
rect 66904 6190 66956 6196
rect 66812 3664 66864 3670
rect 66812 3606 66864 3612
rect 66812 3528 66864 3534
rect 66812 3470 66864 3476
rect 66824 1426 66852 3470
rect 66812 1420 66864 1426
rect 66812 1362 66864 1368
rect 66916 800 66944 6190
rect 67008 5658 67036 7126
rect 67100 6254 67128 8366
rect 67192 7954 67220 10406
rect 67272 9376 67324 9382
rect 67272 9318 67324 9324
rect 67180 7948 67232 7954
rect 67180 7890 67232 7896
rect 67088 6248 67140 6254
rect 67088 6190 67140 6196
rect 67008 5630 67128 5658
rect 66996 5024 67048 5030
rect 66996 4966 67048 4972
rect 67008 4078 67036 4966
rect 66996 4072 67048 4078
rect 66996 4014 67048 4020
rect 66996 3460 67048 3466
rect 66996 3402 67048 3408
rect 67008 800 67036 3402
rect 67100 2922 67128 5630
rect 67088 2916 67140 2922
rect 67088 2858 67140 2864
rect 67192 800 67220 7890
rect 67284 6866 67312 9318
rect 67272 6860 67324 6866
rect 67272 6802 67324 6808
rect 67284 3534 67312 6802
rect 67376 3670 67404 11494
rect 67652 11218 67680 11494
rect 67640 11212 67692 11218
rect 67640 11154 67692 11160
rect 67456 10600 67508 10606
rect 67456 10542 67508 10548
rect 67468 8430 67496 10542
rect 67548 10532 67600 10538
rect 67548 10474 67600 10480
rect 67456 8424 67508 8430
rect 67456 8366 67508 8372
rect 67560 8242 67588 10474
rect 67652 10198 67680 11154
rect 67640 10192 67692 10198
rect 67640 10134 67692 10140
rect 67824 9172 67876 9178
rect 67824 9114 67876 9120
rect 67732 8900 67784 8906
rect 67732 8842 67784 8848
rect 67468 8214 67588 8242
rect 67468 4434 67496 8214
rect 67640 7948 67692 7954
rect 67640 7890 67692 7896
rect 67548 6656 67600 6662
rect 67548 6598 67600 6604
rect 67560 6254 67588 6598
rect 67548 6248 67600 6254
rect 67548 6190 67600 6196
rect 67560 4593 67588 6190
rect 67546 4584 67602 4593
rect 67546 4519 67602 4528
rect 67468 4406 67588 4434
rect 67456 4004 67508 4010
rect 67456 3946 67508 3952
rect 67364 3664 67416 3670
rect 67468 3641 67496 3946
rect 67364 3606 67416 3612
rect 67454 3632 67510 3641
rect 67454 3567 67510 3576
rect 67272 3528 67324 3534
rect 67560 3482 67588 4406
rect 67272 3470 67324 3476
rect 67376 3454 67588 3482
rect 67376 2582 67404 3454
rect 67454 3224 67510 3233
rect 67454 3159 67510 3168
rect 67364 2576 67416 2582
rect 67364 2518 67416 2524
rect 67272 1420 67324 1426
rect 67272 1362 67324 1368
rect 67284 800 67312 1362
rect 67468 800 67496 3159
rect 67652 2774 67680 7890
rect 67744 6866 67772 8842
rect 67836 7342 67864 9114
rect 67824 7336 67876 7342
rect 67824 7278 67876 7284
rect 67824 6996 67876 7002
rect 67824 6938 67876 6944
rect 67732 6860 67784 6866
rect 67732 6802 67784 6808
rect 67560 2746 67680 2774
rect 67560 800 67588 2746
rect 67744 800 67772 6802
rect 67836 5846 67864 6938
rect 67824 5840 67876 5846
rect 67824 5782 67876 5788
rect 67824 4548 67876 4554
rect 67824 4490 67876 4496
rect 67836 800 67864 4490
rect 67928 3058 67956 12406
rect 68112 12306 68140 12407
rect 68100 12300 68152 12306
rect 68100 12242 68152 12248
rect 68098 11112 68154 11121
rect 68098 11047 68100 11056
rect 68152 11047 68154 11056
rect 68100 11018 68152 11024
rect 68008 10464 68060 10470
rect 68008 10406 68060 10412
rect 68020 7954 68048 10406
rect 68100 9988 68152 9994
rect 68100 9930 68152 9936
rect 68112 9897 68140 9930
rect 68098 9888 68154 9897
rect 68098 9823 68154 9832
rect 68100 9444 68152 9450
rect 68100 9386 68152 9392
rect 68112 9042 68140 9386
rect 68100 9036 68152 9042
rect 68100 8978 68152 8984
rect 68836 9036 68888 9042
rect 68836 8978 68888 8984
rect 68100 8832 68152 8838
rect 68100 8774 68152 8780
rect 68112 8537 68140 8774
rect 68098 8528 68154 8537
rect 68098 8463 68154 8472
rect 68112 8430 68140 8463
rect 68100 8424 68152 8430
rect 68100 8366 68152 8372
rect 68192 8356 68244 8362
rect 68192 8298 68244 8304
rect 68008 7948 68060 7954
rect 68008 7890 68060 7896
rect 68204 7834 68232 8298
rect 68020 7806 68232 7834
rect 68284 7880 68336 7886
rect 68284 7822 68336 7828
rect 67916 3052 67968 3058
rect 67916 2994 67968 3000
rect 68020 800 68048 7806
rect 68100 7268 68152 7274
rect 68100 7210 68152 7216
rect 68112 7177 68140 7210
rect 68098 7168 68154 7177
rect 68098 7103 68154 7112
rect 68098 5808 68154 5817
rect 68098 5743 68100 5752
rect 68152 5743 68154 5752
rect 68100 5714 68152 5720
rect 68296 5137 68324 7822
rect 68468 6792 68520 6798
rect 68468 6734 68520 6740
rect 68282 5128 68338 5137
rect 68282 5063 68338 5072
rect 68192 4140 68244 4146
rect 68192 4082 68244 4088
rect 68098 3224 68154 3233
rect 68098 3159 68154 3168
rect 68112 3126 68140 3159
rect 68100 3120 68152 3126
rect 68100 3062 68152 3068
rect 68204 2774 68232 4082
rect 68296 4010 68324 5063
rect 68284 4004 68336 4010
rect 68284 3946 68336 3952
rect 68284 3528 68336 3534
rect 68284 3470 68336 3476
rect 68112 2746 68232 2774
rect 68112 800 68140 2746
rect 68192 2372 68244 2378
rect 68192 2314 68244 2320
rect 68204 1873 68232 2314
rect 68190 1864 68246 1873
rect 68190 1799 68246 1808
rect 68296 800 68324 3470
rect 68480 800 68508 6734
rect 68744 5092 68796 5098
rect 68744 5034 68796 5040
rect 68560 4072 68612 4078
rect 68560 4014 68612 4020
rect 68572 800 68600 4014
rect 68756 800 68784 5034
rect 68848 800 68876 8978
rect 69296 7404 69348 7410
rect 69296 7346 69348 7352
rect 69020 5704 69072 5710
rect 69020 5646 69072 5652
rect 69032 800 69060 5646
rect 69112 4480 69164 4486
rect 69112 4422 69164 4428
rect 69124 800 69152 4422
rect 69308 800 69336 7346
rect 69848 5636 69900 5642
rect 69848 5578 69900 5584
rect 69664 5024 69716 5030
rect 69664 4966 69716 4972
rect 69572 3936 69624 3942
rect 69572 3878 69624 3884
rect 69388 3188 69440 3194
rect 69388 3130 69440 3136
rect 69400 800 69428 3130
rect 69584 800 69612 3878
rect 69676 800 69704 4966
rect 69860 800 69888 5578
rect 66074 640 66130 649
rect 66074 575 66130 584
rect 66166 0 66222 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68098 0 68154 800
rect 68282 0 68338 800
rect 68466 0 68522 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69662 0 69718 800
rect 69846 0 69902 800
<< via2 >>
rect 67362 69264 67418 69320
rect 2778 67904 2834 67960
rect 1766 66716 1768 66736
rect 1768 66716 1820 66736
rect 1820 66716 1822 66736
rect 1766 66680 1822 66716
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4246 67482
rect 4246 67430 4276 67482
rect 4300 67430 4310 67482
rect 4310 67430 4356 67482
rect 4380 67430 4426 67482
rect 4426 67430 4436 67482
rect 4460 67430 4490 67482
rect 4490 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 14220 67482 14276 67484
rect 14300 67482 14356 67484
rect 14380 67482 14436 67484
rect 14460 67482 14516 67484
rect 14220 67430 14246 67482
rect 14246 67430 14276 67482
rect 14300 67430 14310 67482
rect 14310 67430 14356 67482
rect 14380 67430 14426 67482
rect 14426 67430 14436 67482
rect 14460 67430 14490 67482
rect 14490 67430 14516 67482
rect 14220 67428 14276 67430
rect 14300 67428 14356 67430
rect 14380 67428 14436 67430
rect 14460 67428 14516 67430
rect 24220 67482 24276 67484
rect 24300 67482 24356 67484
rect 24380 67482 24436 67484
rect 24460 67482 24516 67484
rect 24220 67430 24246 67482
rect 24246 67430 24276 67482
rect 24300 67430 24310 67482
rect 24310 67430 24356 67482
rect 24380 67430 24426 67482
rect 24426 67430 24436 67482
rect 24460 67430 24490 67482
rect 24490 67430 24516 67482
rect 24220 67428 24276 67430
rect 24300 67428 24356 67430
rect 24380 67428 24436 67430
rect 24460 67428 24516 67430
rect 34220 67482 34276 67484
rect 34300 67482 34356 67484
rect 34380 67482 34436 67484
rect 34460 67482 34516 67484
rect 34220 67430 34246 67482
rect 34246 67430 34276 67482
rect 34300 67430 34310 67482
rect 34310 67430 34356 67482
rect 34380 67430 34426 67482
rect 34426 67430 34436 67482
rect 34460 67430 34490 67482
rect 34490 67430 34516 67482
rect 34220 67428 34276 67430
rect 34300 67428 34356 67430
rect 34380 67428 34436 67430
rect 34460 67428 34516 67430
rect 44220 67482 44276 67484
rect 44300 67482 44356 67484
rect 44380 67482 44436 67484
rect 44460 67482 44516 67484
rect 44220 67430 44246 67482
rect 44246 67430 44276 67482
rect 44300 67430 44310 67482
rect 44310 67430 44356 67482
rect 44380 67430 44426 67482
rect 44426 67430 44436 67482
rect 44460 67430 44490 67482
rect 44490 67430 44516 67482
rect 44220 67428 44276 67430
rect 44300 67428 44356 67430
rect 44380 67428 44436 67430
rect 44460 67428 44516 67430
rect 54220 67482 54276 67484
rect 54300 67482 54356 67484
rect 54380 67482 54436 67484
rect 54460 67482 54516 67484
rect 54220 67430 54246 67482
rect 54246 67430 54276 67482
rect 54300 67430 54310 67482
rect 54310 67430 54356 67482
rect 54380 67430 54426 67482
rect 54426 67430 54436 67482
rect 54460 67430 54490 67482
rect 54490 67430 54516 67482
rect 54220 67428 54276 67430
rect 54300 67428 54356 67430
rect 54380 67428 54436 67430
rect 54460 67428 54516 67430
rect 64220 67482 64276 67484
rect 64300 67482 64356 67484
rect 64380 67482 64436 67484
rect 64460 67482 64516 67484
rect 64220 67430 64246 67482
rect 64246 67430 64276 67482
rect 64300 67430 64310 67482
rect 64310 67430 64356 67482
rect 64380 67430 64426 67482
rect 64426 67430 64436 67482
rect 64460 67430 64490 67482
rect 64490 67430 64516 67482
rect 64220 67428 64276 67430
rect 64300 67428 64356 67430
rect 64380 67428 64436 67430
rect 64460 67428 64516 67430
rect 67546 67904 67602 67960
rect 9220 66938 9276 66940
rect 9300 66938 9356 66940
rect 9380 66938 9436 66940
rect 9460 66938 9516 66940
rect 9220 66886 9246 66938
rect 9246 66886 9276 66938
rect 9300 66886 9310 66938
rect 9310 66886 9356 66938
rect 9380 66886 9426 66938
rect 9426 66886 9436 66938
rect 9460 66886 9490 66938
rect 9490 66886 9516 66938
rect 9220 66884 9276 66886
rect 9300 66884 9356 66886
rect 9380 66884 9436 66886
rect 9460 66884 9516 66886
rect 1858 65356 1860 65376
rect 1860 65356 1912 65376
rect 1912 65356 1914 65376
rect 1858 65320 1914 65356
rect 1582 62772 1584 62792
rect 1584 62772 1636 62792
rect 1636 62772 1638 62792
rect 1582 62736 1638 62772
rect 1858 61548 1860 61568
rect 1860 61548 1912 61568
rect 1912 61548 1914 61568
rect 1858 61512 1914 61548
rect 1766 60172 1822 60208
rect 1766 60152 1768 60172
rect 1768 60152 1820 60172
rect 1820 60152 1822 60172
rect 1582 57568 1638 57624
rect 1766 56364 1822 56400
rect 1766 56344 1768 56364
rect 1768 56344 1820 56364
rect 1820 56344 1822 56364
rect 1858 55020 1860 55040
rect 1860 55020 1912 55040
rect 1912 55020 1914 55040
rect 1858 54984 1914 55020
rect 1582 52400 1638 52456
rect 1858 51060 1914 51096
rect 1858 51040 1860 51060
rect 1860 51040 1912 51060
rect 1912 51040 1914 51060
rect 1766 49836 1822 49872
rect 1766 49816 1768 49836
rect 1768 49816 1820 49836
rect 1820 49816 1822 49836
rect 1858 47232 1914 47288
rect 1766 45908 1768 45928
rect 1768 45908 1820 45928
rect 1820 45908 1822 45928
rect 1766 45872 1822 45908
rect 1858 44684 1860 44704
rect 1860 44684 1912 44704
rect 1912 44684 1914 44704
rect 1858 44648 1914 44684
rect 1582 42100 1584 42120
rect 1584 42100 1636 42120
rect 1636 42100 1638 42120
rect 1582 42064 1638 42100
rect 1858 40724 1914 40760
rect 1858 40704 1860 40724
rect 1860 40704 1912 40724
rect 1912 40704 1914 40724
rect 1766 39500 1822 39536
rect 1766 39480 1768 39500
rect 1768 39480 1820 39500
rect 1820 39480 1822 39500
rect 1582 36896 1638 36952
rect 1766 35572 1768 35592
rect 1768 35572 1820 35592
rect 1820 35572 1822 35592
rect 1766 35536 1822 35572
rect 1858 34196 1914 34232
rect 1858 34176 1860 34196
rect 1860 34176 1912 34196
rect 1912 34176 1914 34196
rect 1582 31592 1638 31648
rect 1766 30368 1822 30424
rect 1766 29044 1768 29064
rect 1768 29044 1820 29064
rect 1820 29044 1822 29064
rect 1766 29008 1822 29044
rect 1582 26424 1638 26480
rect 1766 25220 1822 25256
rect 1766 25200 1768 25220
rect 1768 25200 1820 25220
rect 1820 25200 1822 25220
rect 1858 23860 1914 23896
rect 1858 23840 1860 23860
rect 1860 23840 1912 23860
rect 1912 23840 1914 23860
rect 1398 21256 1454 21312
rect 1858 20052 1914 20088
rect 1858 20032 1860 20052
rect 1860 20032 1912 20052
rect 1912 20032 1914 20052
rect 1766 18692 1822 18728
rect 1766 18672 1768 18692
rect 1768 18672 1820 18692
rect 1820 18672 1822 18692
rect 1582 16088 1638 16144
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4246 66394
rect 4246 66342 4276 66394
rect 4300 66342 4310 66394
rect 4310 66342 4356 66394
rect 4380 66342 4426 66394
rect 4426 66342 4436 66394
rect 4460 66342 4490 66394
rect 4490 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 9220 65850 9276 65852
rect 9300 65850 9356 65852
rect 9380 65850 9436 65852
rect 9460 65850 9516 65852
rect 9220 65798 9246 65850
rect 9246 65798 9276 65850
rect 9300 65798 9310 65850
rect 9310 65798 9356 65850
rect 9380 65798 9426 65850
rect 9426 65798 9436 65850
rect 9460 65798 9490 65850
rect 9490 65798 9516 65850
rect 9220 65796 9276 65798
rect 9300 65796 9356 65798
rect 9380 65796 9436 65798
rect 9460 65796 9516 65798
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4246 65306
rect 4246 65254 4276 65306
rect 4300 65254 4310 65306
rect 4310 65254 4356 65306
rect 4380 65254 4426 65306
rect 4426 65254 4436 65306
rect 4460 65254 4490 65306
rect 4490 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4246 64218
rect 4246 64166 4276 64218
rect 4300 64166 4310 64218
rect 4310 64166 4356 64218
rect 4380 64166 4426 64218
rect 4426 64166 4436 64218
rect 4460 64166 4490 64218
rect 4490 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4246 63130
rect 4246 63078 4276 63130
rect 4300 63078 4310 63130
rect 4310 63078 4356 63130
rect 4380 63078 4426 63130
rect 4426 63078 4436 63130
rect 4460 63078 4490 63130
rect 4490 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4246 62042
rect 4246 61990 4276 62042
rect 4300 61990 4310 62042
rect 4310 61990 4356 62042
rect 4380 61990 4426 62042
rect 4426 61990 4436 62042
rect 4460 61990 4490 62042
rect 4490 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4246 60954
rect 4246 60902 4276 60954
rect 4300 60902 4310 60954
rect 4310 60902 4356 60954
rect 4380 60902 4426 60954
rect 4426 60902 4436 60954
rect 4460 60902 4490 60954
rect 4490 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4246 59866
rect 4246 59814 4276 59866
rect 4300 59814 4310 59866
rect 4310 59814 4356 59866
rect 4380 59814 4426 59866
rect 4426 59814 4436 59866
rect 4460 59814 4490 59866
rect 4490 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4246 58778
rect 4246 58726 4276 58778
rect 4300 58726 4310 58778
rect 4310 58726 4356 58778
rect 4380 58726 4426 58778
rect 4426 58726 4436 58778
rect 4460 58726 4490 58778
rect 4490 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 1858 14764 1860 14784
rect 1860 14764 1912 14784
rect 1912 14764 1914 14784
rect 1858 14728 1914 14764
rect 1858 13524 1914 13560
rect 1858 13504 1860 13524
rect 1860 13504 1912 13524
rect 1912 13504 1914 13524
rect 1582 10920 1638 10976
rect 1766 9596 1768 9616
rect 1768 9596 1820 9616
rect 1820 9596 1822 9616
rect 1766 9560 1822 9596
rect 2686 11056 2742 11112
rect 1582 6976 1638 7032
rect 1766 8372 1768 8392
rect 1768 8372 1820 8392
rect 1820 8372 1822 8392
rect 1766 8336 1822 8372
rect 1766 5788 1768 5808
rect 1768 5788 1820 5808
rect 1820 5788 1822 5808
rect 1766 5752 1822 5788
rect 1582 3168 1638 3224
rect 1858 4428 1860 4448
rect 1860 4428 1912 4448
rect 1912 4428 1914 4448
rect 1858 4392 1914 4428
rect 1858 1808 1914 1864
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 9220 64762 9276 64764
rect 9300 64762 9356 64764
rect 9380 64762 9436 64764
rect 9460 64762 9516 64764
rect 9220 64710 9246 64762
rect 9246 64710 9276 64762
rect 9300 64710 9310 64762
rect 9310 64710 9356 64762
rect 9380 64710 9426 64762
rect 9426 64710 9436 64762
rect 9460 64710 9490 64762
rect 9490 64710 9516 64762
rect 9220 64708 9276 64710
rect 9300 64708 9356 64710
rect 9380 64708 9436 64710
rect 9460 64708 9516 64710
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 3974 5208 4030 5264
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 4526 1944 4582 2000
rect 5262 2760 5318 2816
rect 5446 5108 5448 5128
rect 5448 5108 5500 5128
rect 5500 5108 5502 5128
rect 5446 5072 5502 5108
rect 5722 7148 5724 7168
rect 5724 7148 5776 7168
rect 5776 7148 5778 7168
rect 5722 7112 5778 7148
rect 9220 63674 9276 63676
rect 9300 63674 9356 63676
rect 9380 63674 9436 63676
rect 9460 63674 9516 63676
rect 9220 63622 9246 63674
rect 9246 63622 9276 63674
rect 9300 63622 9310 63674
rect 9310 63622 9356 63674
rect 9380 63622 9426 63674
rect 9426 63622 9436 63674
rect 9460 63622 9490 63674
rect 9490 63622 9516 63674
rect 9220 63620 9276 63622
rect 9300 63620 9356 63622
rect 9380 63620 9436 63622
rect 9460 63620 9516 63622
rect 9220 62586 9276 62588
rect 9300 62586 9356 62588
rect 9380 62586 9436 62588
rect 9460 62586 9516 62588
rect 9220 62534 9246 62586
rect 9246 62534 9276 62586
rect 9300 62534 9310 62586
rect 9310 62534 9356 62586
rect 9380 62534 9426 62586
rect 9426 62534 9436 62586
rect 9460 62534 9490 62586
rect 9490 62534 9516 62586
rect 9220 62532 9276 62534
rect 9300 62532 9356 62534
rect 9380 62532 9436 62534
rect 9460 62532 9516 62534
rect 9220 61498 9276 61500
rect 9300 61498 9356 61500
rect 9380 61498 9436 61500
rect 9460 61498 9516 61500
rect 9220 61446 9246 61498
rect 9246 61446 9276 61498
rect 9300 61446 9310 61498
rect 9310 61446 9356 61498
rect 9380 61446 9426 61498
rect 9426 61446 9436 61498
rect 9460 61446 9490 61498
rect 9490 61446 9516 61498
rect 9220 61444 9276 61446
rect 9300 61444 9356 61446
rect 9380 61444 9436 61446
rect 9460 61444 9516 61446
rect 9220 60410 9276 60412
rect 9300 60410 9356 60412
rect 9380 60410 9436 60412
rect 9460 60410 9516 60412
rect 9220 60358 9246 60410
rect 9246 60358 9276 60410
rect 9300 60358 9310 60410
rect 9310 60358 9356 60410
rect 9380 60358 9426 60410
rect 9426 60358 9436 60410
rect 9460 60358 9490 60410
rect 9490 60358 9516 60410
rect 9220 60356 9276 60358
rect 9300 60356 9356 60358
rect 9380 60356 9436 60358
rect 9460 60356 9516 60358
rect 9220 59322 9276 59324
rect 9300 59322 9356 59324
rect 9380 59322 9436 59324
rect 9460 59322 9516 59324
rect 9220 59270 9246 59322
rect 9246 59270 9276 59322
rect 9300 59270 9310 59322
rect 9310 59270 9356 59322
rect 9380 59270 9426 59322
rect 9426 59270 9436 59322
rect 9460 59270 9490 59322
rect 9490 59270 9516 59322
rect 9220 59268 9276 59270
rect 9300 59268 9356 59270
rect 9380 59268 9436 59270
rect 9460 59268 9516 59270
rect 9220 58234 9276 58236
rect 9300 58234 9356 58236
rect 9380 58234 9436 58236
rect 9460 58234 9516 58236
rect 9220 58182 9246 58234
rect 9246 58182 9276 58234
rect 9300 58182 9310 58234
rect 9310 58182 9356 58234
rect 9380 58182 9426 58234
rect 9426 58182 9436 58234
rect 9460 58182 9490 58234
rect 9490 58182 9516 58234
rect 9220 58180 9276 58182
rect 9300 58180 9356 58182
rect 9380 58180 9436 58182
rect 9460 58180 9516 58182
rect 5998 2760 6054 2816
rect 7194 32408 7250 32464
rect 6826 4156 6828 4176
rect 6828 4156 6880 4176
rect 6880 4156 6882 4176
rect 6826 4120 6882 4156
rect 7378 21392 7434 21448
rect 9220 57146 9276 57148
rect 9300 57146 9356 57148
rect 9380 57146 9436 57148
rect 9460 57146 9516 57148
rect 9220 57094 9246 57146
rect 9246 57094 9276 57146
rect 9300 57094 9310 57146
rect 9310 57094 9356 57146
rect 9380 57094 9426 57146
rect 9426 57094 9436 57146
rect 9460 57094 9490 57146
rect 9490 57094 9516 57146
rect 9220 57092 9276 57094
rect 9300 57092 9356 57094
rect 9380 57092 9436 57094
rect 9460 57092 9516 57094
rect 9220 56058 9276 56060
rect 9300 56058 9356 56060
rect 9380 56058 9436 56060
rect 9460 56058 9516 56060
rect 9220 56006 9246 56058
rect 9246 56006 9276 56058
rect 9300 56006 9310 56058
rect 9310 56006 9356 56058
rect 9380 56006 9426 56058
rect 9426 56006 9436 56058
rect 9460 56006 9490 56058
rect 9490 56006 9516 56058
rect 9220 56004 9276 56006
rect 9300 56004 9356 56006
rect 9380 56004 9436 56006
rect 9460 56004 9516 56006
rect 9220 54970 9276 54972
rect 9300 54970 9356 54972
rect 9380 54970 9436 54972
rect 9460 54970 9516 54972
rect 9220 54918 9246 54970
rect 9246 54918 9276 54970
rect 9300 54918 9310 54970
rect 9310 54918 9356 54970
rect 9380 54918 9426 54970
rect 9426 54918 9436 54970
rect 9460 54918 9490 54970
rect 9490 54918 9516 54970
rect 9220 54916 9276 54918
rect 9300 54916 9356 54918
rect 9380 54916 9436 54918
rect 9460 54916 9516 54918
rect 9220 53882 9276 53884
rect 9300 53882 9356 53884
rect 9380 53882 9436 53884
rect 9460 53882 9516 53884
rect 9220 53830 9246 53882
rect 9246 53830 9276 53882
rect 9300 53830 9310 53882
rect 9310 53830 9356 53882
rect 9380 53830 9426 53882
rect 9426 53830 9436 53882
rect 9460 53830 9490 53882
rect 9490 53830 9516 53882
rect 9220 53828 9276 53830
rect 9300 53828 9356 53830
rect 9380 53828 9436 53830
rect 9460 53828 9516 53830
rect 9220 52794 9276 52796
rect 9300 52794 9356 52796
rect 9380 52794 9436 52796
rect 9460 52794 9516 52796
rect 9220 52742 9246 52794
rect 9246 52742 9276 52794
rect 9300 52742 9310 52794
rect 9310 52742 9356 52794
rect 9380 52742 9426 52794
rect 9426 52742 9436 52794
rect 9460 52742 9490 52794
rect 9490 52742 9516 52794
rect 9220 52740 9276 52742
rect 9300 52740 9356 52742
rect 9380 52740 9436 52742
rect 9460 52740 9516 52742
rect 9220 51706 9276 51708
rect 9300 51706 9356 51708
rect 9380 51706 9436 51708
rect 9460 51706 9516 51708
rect 9220 51654 9246 51706
rect 9246 51654 9276 51706
rect 9300 51654 9310 51706
rect 9310 51654 9356 51706
rect 9380 51654 9426 51706
rect 9426 51654 9436 51706
rect 9460 51654 9490 51706
rect 9490 51654 9516 51706
rect 9220 51652 9276 51654
rect 9300 51652 9356 51654
rect 9380 51652 9436 51654
rect 9460 51652 9516 51654
rect 9220 50618 9276 50620
rect 9300 50618 9356 50620
rect 9380 50618 9436 50620
rect 9460 50618 9516 50620
rect 9220 50566 9246 50618
rect 9246 50566 9276 50618
rect 9300 50566 9310 50618
rect 9310 50566 9356 50618
rect 9380 50566 9426 50618
rect 9426 50566 9436 50618
rect 9460 50566 9490 50618
rect 9490 50566 9516 50618
rect 9220 50564 9276 50566
rect 9300 50564 9356 50566
rect 9380 50564 9436 50566
rect 9460 50564 9516 50566
rect 9220 49530 9276 49532
rect 9300 49530 9356 49532
rect 9380 49530 9436 49532
rect 9460 49530 9516 49532
rect 9220 49478 9246 49530
rect 9246 49478 9276 49530
rect 9300 49478 9310 49530
rect 9310 49478 9356 49530
rect 9380 49478 9426 49530
rect 9426 49478 9436 49530
rect 9460 49478 9490 49530
rect 9490 49478 9516 49530
rect 9220 49476 9276 49478
rect 9300 49476 9356 49478
rect 9380 49476 9436 49478
rect 9460 49476 9516 49478
rect 9220 48442 9276 48444
rect 9300 48442 9356 48444
rect 9380 48442 9436 48444
rect 9460 48442 9516 48444
rect 9220 48390 9246 48442
rect 9246 48390 9276 48442
rect 9300 48390 9310 48442
rect 9310 48390 9356 48442
rect 9380 48390 9426 48442
rect 9426 48390 9436 48442
rect 9460 48390 9490 48442
rect 9490 48390 9516 48442
rect 9220 48388 9276 48390
rect 9300 48388 9356 48390
rect 9380 48388 9436 48390
rect 9460 48388 9516 48390
rect 9220 47354 9276 47356
rect 9300 47354 9356 47356
rect 9380 47354 9436 47356
rect 9460 47354 9516 47356
rect 9220 47302 9246 47354
rect 9246 47302 9276 47354
rect 9300 47302 9310 47354
rect 9310 47302 9356 47354
rect 9380 47302 9426 47354
rect 9426 47302 9436 47354
rect 9460 47302 9490 47354
rect 9490 47302 9516 47354
rect 9220 47300 9276 47302
rect 9300 47300 9356 47302
rect 9380 47300 9436 47302
rect 9460 47300 9516 47302
rect 9220 46266 9276 46268
rect 9300 46266 9356 46268
rect 9380 46266 9436 46268
rect 9460 46266 9516 46268
rect 9220 46214 9246 46266
rect 9246 46214 9276 46266
rect 9300 46214 9310 46266
rect 9310 46214 9356 46266
rect 9380 46214 9426 46266
rect 9426 46214 9436 46266
rect 9460 46214 9490 46266
rect 9490 46214 9516 46266
rect 9220 46212 9276 46214
rect 9300 46212 9356 46214
rect 9380 46212 9436 46214
rect 9460 46212 9516 46214
rect 9220 45178 9276 45180
rect 9300 45178 9356 45180
rect 9380 45178 9436 45180
rect 9460 45178 9516 45180
rect 9220 45126 9246 45178
rect 9246 45126 9276 45178
rect 9300 45126 9310 45178
rect 9310 45126 9356 45178
rect 9380 45126 9426 45178
rect 9426 45126 9436 45178
rect 9460 45126 9490 45178
rect 9490 45126 9516 45178
rect 9220 45124 9276 45126
rect 9300 45124 9356 45126
rect 9380 45124 9436 45126
rect 9460 45124 9516 45126
rect 9220 44090 9276 44092
rect 9300 44090 9356 44092
rect 9380 44090 9436 44092
rect 9460 44090 9516 44092
rect 9220 44038 9246 44090
rect 9246 44038 9276 44090
rect 9300 44038 9310 44090
rect 9310 44038 9356 44090
rect 9380 44038 9426 44090
rect 9426 44038 9436 44090
rect 9460 44038 9490 44090
rect 9490 44038 9516 44090
rect 9220 44036 9276 44038
rect 9300 44036 9356 44038
rect 9380 44036 9436 44038
rect 9460 44036 9516 44038
rect 9220 43002 9276 43004
rect 9300 43002 9356 43004
rect 9380 43002 9436 43004
rect 9460 43002 9516 43004
rect 9220 42950 9246 43002
rect 9246 42950 9276 43002
rect 9300 42950 9310 43002
rect 9310 42950 9356 43002
rect 9380 42950 9426 43002
rect 9426 42950 9436 43002
rect 9460 42950 9490 43002
rect 9490 42950 9516 43002
rect 9220 42948 9276 42950
rect 9300 42948 9356 42950
rect 9380 42948 9436 42950
rect 9460 42948 9516 42950
rect 9220 41914 9276 41916
rect 9300 41914 9356 41916
rect 9380 41914 9436 41916
rect 9460 41914 9516 41916
rect 9220 41862 9246 41914
rect 9246 41862 9276 41914
rect 9300 41862 9310 41914
rect 9310 41862 9356 41914
rect 9380 41862 9426 41914
rect 9426 41862 9436 41914
rect 9460 41862 9490 41914
rect 9490 41862 9516 41914
rect 9220 41860 9276 41862
rect 9300 41860 9356 41862
rect 9380 41860 9436 41862
rect 9460 41860 9516 41862
rect 9220 40826 9276 40828
rect 9300 40826 9356 40828
rect 9380 40826 9436 40828
rect 9460 40826 9516 40828
rect 9220 40774 9246 40826
rect 9246 40774 9276 40826
rect 9300 40774 9310 40826
rect 9310 40774 9356 40826
rect 9380 40774 9426 40826
rect 9426 40774 9436 40826
rect 9460 40774 9490 40826
rect 9490 40774 9516 40826
rect 9220 40772 9276 40774
rect 9300 40772 9356 40774
rect 9380 40772 9436 40774
rect 9460 40772 9516 40774
rect 9220 39738 9276 39740
rect 9300 39738 9356 39740
rect 9380 39738 9436 39740
rect 9460 39738 9516 39740
rect 9220 39686 9246 39738
rect 9246 39686 9276 39738
rect 9300 39686 9310 39738
rect 9310 39686 9356 39738
rect 9380 39686 9426 39738
rect 9426 39686 9436 39738
rect 9460 39686 9490 39738
rect 9490 39686 9516 39738
rect 9220 39684 9276 39686
rect 9300 39684 9356 39686
rect 9380 39684 9436 39686
rect 9460 39684 9516 39686
rect 9220 38650 9276 38652
rect 9300 38650 9356 38652
rect 9380 38650 9436 38652
rect 9460 38650 9516 38652
rect 9220 38598 9246 38650
rect 9246 38598 9276 38650
rect 9300 38598 9310 38650
rect 9310 38598 9356 38650
rect 9380 38598 9426 38650
rect 9426 38598 9436 38650
rect 9460 38598 9490 38650
rect 9490 38598 9516 38650
rect 9220 38596 9276 38598
rect 9300 38596 9356 38598
rect 9380 38596 9436 38598
rect 9460 38596 9516 38598
rect 9220 37562 9276 37564
rect 9300 37562 9356 37564
rect 9380 37562 9436 37564
rect 9460 37562 9516 37564
rect 9220 37510 9246 37562
rect 9246 37510 9276 37562
rect 9300 37510 9310 37562
rect 9310 37510 9356 37562
rect 9380 37510 9426 37562
rect 9426 37510 9436 37562
rect 9460 37510 9490 37562
rect 9490 37510 9516 37562
rect 9220 37508 9276 37510
rect 9300 37508 9356 37510
rect 9380 37508 9436 37510
rect 9460 37508 9516 37510
rect 9220 36474 9276 36476
rect 9300 36474 9356 36476
rect 9380 36474 9436 36476
rect 9460 36474 9516 36476
rect 9220 36422 9246 36474
rect 9246 36422 9276 36474
rect 9300 36422 9310 36474
rect 9310 36422 9356 36474
rect 9380 36422 9426 36474
rect 9426 36422 9436 36474
rect 9460 36422 9490 36474
rect 9490 36422 9516 36474
rect 9220 36420 9276 36422
rect 9300 36420 9356 36422
rect 9380 36420 9436 36422
rect 9460 36420 9516 36422
rect 9220 35386 9276 35388
rect 9300 35386 9356 35388
rect 9380 35386 9436 35388
rect 9460 35386 9516 35388
rect 9220 35334 9246 35386
rect 9246 35334 9276 35386
rect 9300 35334 9310 35386
rect 9310 35334 9356 35386
rect 9380 35334 9426 35386
rect 9426 35334 9436 35386
rect 9460 35334 9490 35386
rect 9490 35334 9516 35386
rect 9220 35332 9276 35334
rect 9300 35332 9356 35334
rect 9380 35332 9436 35334
rect 9460 35332 9516 35334
rect 9220 34298 9276 34300
rect 9300 34298 9356 34300
rect 9380 34298 9436 34300
rect 9460 34298 9516 34300
rect 9220 34246 9246 34298
rect 9246 34246 9276 34298
rect 9300 34246 9310 34298
rect 9310 34246 9356 34298
rect 9380 34246 9426 34298
rect 9426 34246 9436 34298
rect 9460 34246 9490 34298
rect 9490 34246 9516 34298
rect 9220 34244 9276 34246
rect 9300 34244 9356 34246
rect 9380 34244 9436 34246
rect 9460 34244 9516 34246
rect 9220 33210 9276 33212
rect 9300 33210 9356 33212
rect 9380 33210 9436 33212
rect 9460 33210 9516 33212
rect 9220 33158 9246 33210
rect 9246 33158 9276 33210
rect 9300 33158 9310 33210
rect 9310 33158 9356 33210
rect 9380 33158 9426 33210
rect 9426 33158 9436 33210
rect 9460 33158 9490 33210
rect 9490 33158 9516 33210
rect 9220 33156 9276 33158
rect 9300 33156 9356 33158
rect 9380 33156 9436 33158
rect 9460 33156 9516 33158
rect 9220 32122 9276 32124
rect 9300 32122 9356 32124
rect 9380 32122 9436 32124
rect 9460 32122 9516 32124
rect 9220 32070 9246 32122
rect 9246 32070 9276 32122
rect 9300 32070 9310 32122
rect 9310 32070 9356 32122
rect 9380 32070 9426 32122
rect 9426 32070 9436 32122
rect 9460 32070 9490 32122
rect 9490 32070 9516 32122
rect 9220 32068 9276 32070
rect 9300 32068 9356 32070
rect 9380 32068 9436 32070
rect 9460 32068 9516 32070
rect 9220 31034 9276 31036
rect 9300 31034 9356 31036
rect 9380 31034 9436 31036
rect 9460 31034 9516 31036
rect 9220 30982 9246 31034
rect 9246 30982 9276 31034
rect 9300 30982 9310 31034
rect 9310 30982 9356 31034
rect 9380 30982 9426 31034
rect 9426 30982 9436 31034
rect 9460 30982 9490 31034
rect 9490 30982 9516 31034
rect 9220 30980 9276 30982
rect 9300 30980 9356 30982
rect 9380 30980 9436 30982
rect 9460 30980 9516 30982
rect 9220 29946 9276 29948
rect 9300 29946 9356 29948
rect 9380 29946 9436 29948
rect 9460 29946 9516 29948
rect 9220 29894 9246 29946
rect 9246 29894 9276 29946
rect 9300 29894 9310 29946
rect 9310 29894 9356 29946
rect 9380 29894 9426 29946
rect 9426 29894 9436 29946
rect 9460 29894 9490 29946
rect 9490 29894 9516 29946
rect 9220 29892 9276 29894
rect 9300 29892 9356 29894
rect 9380 29892 9436 29894
rect 9460 29892 9516 29894
rect 9220 28858 9276 28860
rect 9300 28858 9356 28860
rect 9380 28858 9436 28860
rect 9460 28858 9516 28860
rect 9220 28806 9246 28858
rect 9246 28806 9276 28858
rect 9300 28806 9310 28858
rect 9310 28806 9356 28858
rect 9380 28806 9426 28858
rect 9426 28806 9436 28858
rect 9460 28806 9490 28858
rect 9490 28806 9516 28858
rect 9220 28804 9276 28806
rect 9300 28804 9356 28806
rect 9380 28804 9436 28806
rect 9460 28804 9516 28806
rect 9220 27770 9276 27772
rect 9300 27770 9356 27772
rect 9380 27770 9436 27772
rect 9460 27770 9516 27772
rect 9220 27718 9246 27770
rect 9246 27718 9276 27770
rect 9300 27718 9310 27770
rect 9310 27718 9356 27770
rect 9380 27718 9426 27770
rect 9426 27718 9436 27770
rect 9460 27718 9490 27770
rect 9490 27718 9516 27770
rect 9220 27716 9276 27718
rect 9300 27716 9356 27718
rect 9380 27716 9436 27718
rect 9460 27716 9516 27718
rect 9220 26682 9276 26684
rect 9300 26682 9356 26684
rect 9380 26682 9436 26684
rect 9460 26682 9516 26684
rect 9220 26630 9246 26682
rect 9246 26630 9276 26682
rect 9300 26630 9310 26682
rect 9310 26630 9356 26682
rect 9380 26630 9426 26682
rect 9426 26630 9436 26682
rect 9460 26630 9490 26682
rect 9490 26630 9516 26682
rect 9220 26628 9276 26630
rect 9300 26628 9356 26630
rect 9380 26628 9436 26630
rect 9460 26628 9516 26630
rect 9220 25594 9276 25596
rect 9300 25594 9356 25596
rect 9380 25594 9436 25596
rect 9460 25594 9516 25596
rect 9220 25542 9246 25594
rect 9246 25542 9276 25594
rect 9300 25542 9310 25594
rect 9310 25542 9356 25594
rect 9380 25542 9426 25594
rect 9426 25542 9436 25594
rect 9460 25542 9490 25594
rect 9490 25542 9516 25594
rect 9220 25540 9276 25542
rect 9300 25540 9356 25542
rect 9380 25540 9436 25542
rect 9460 25540 9516 25542
rect 9220 24506 9276 24508
rect 9300 24506 9356 24508
rect 9380 24506 9436 24508
rect 9460 24506 9516 24508
rect 9220 24454 9246 24506
rect 9246 24454 9276 24506
rect 9300 24454 9310 24506
rect 9310 24454 9356 24506
rect 9380 24454 9426 24506
rect 9426 24454 9436 24506
rect 9460 24454 9490 24506
rect 9490 24454 9516 24506
rect 9220 24452 9276 24454
rect 9300 24452 9356 24454
rect 9380 24452 9436 24454
rect 9460 24452 9516 24454
rect 9220 23418 9276 23420
rect 9300 23418 9356 23420
rect 9380 23418 9436 23420
rect 9460 23418 9516 23420
rect 9220 23366 9246 23418
rect 9246 23366 9276 23418
rect 9300 23366 9310 23418
rect 9310 23366 9356 23418
rect 9380 23366 9426 23418
rect 9426 23366 9436 23418
rect 9460 23366 9490 23418
rect 9490 23366 9516 23418
rect 9220 23364 9276 23366
rect 9300 23364 9356 23366
rect 9380 23364 9436 23366
rect 9460 23364 9516 23366
rect 9220 22330 9276 22332
rect 9300 22330 9356 22332
rect 9380 22330 9436 22332
rect 9460 22330 9516 22332
rect 9220 22278 9246 22330
rect 9246 22278 9276 22330
rect 9300 22278 9310 22330
rect 9310 22278 9356 22330
rect 9380 22278 9426 22330
rect 9426 22278 9436 22330
rect 9460 22278 9490 22330
rect 9490 22278 9516 22330
rect 9220 22276 9276 22278
rect 9300 22276 9356 22278
rect 9380 22276 9436 22278
rect 9460 22276 9516 22278
rect 9220 21242 9276 21244
rect 9300 21242 9356 21244
rect 9380 21242 9436 21244
rect 9460 21242 9516 21244
rect 9220 21190 9246 21242
rect 9246 21190 9276 21242
rect 9300 21190 9310 21242
rect 9310 21190 9356 21242
rect 9380 21190 9426 21242
rect 9426 21190 9436 21242
rect 9460 21190 9490 21242
rect 9490 21190 9516 21242
rect 9220 21188 9276 21190
rect 9300 21188 9356 21190
rect 9380 21188 9436 21190
rect 9460 21188 9516 21190
rect 9220 20154 9276 20156
rect 9300 20154 9356 20156
rect 9380 20154 9436 20156
rect 9460 20154 9516 20156
rect 9220 20102 9246 20154
rect 9246 20102 9276 20154
rect 9300 20102 9310 20154
rect 9310 20102 9356 20154
rect 9380 20102 9426 20154
rect 9426 20102 9436 20154
rect 9460 20102 9490 20154
rect 9490 20102 9516 20154
rect 9220 20100 9276 20102
rect 9300 20100 9356 20102
rect 9380 20100 9436 20102
rect 9460 20100 9516 20102
rect 9220 19066 9276 19068
rect 9300 19066 9356 19068
rect 9380 19066 9436 19068
rect 9460 19066 9516 19068
rect 9220 19014 9246 19066
rect 9246 19014 9276 19066
rect 9300 19014 9310 19066
rect 9310 19014 9356 19066
rect 9380 19014 9426 19066
rect 9426 19014 9436 19066
rect 9460 19014 9490 19066
rect 9490 19014 9516 19066
rect 9220 19012 9276 19014
rect 9300 19012 9356 19014
rect 9380 19012 9436 19014
rect 9460 19012 9516 19014
rect 9220 17978 9276 17980
rect 9300 17978 9356 17980
rect 9380 17978 9436 17980
rect 9460 17978 9516 17980
rect 9220 17926 9246 17978
rect 9246 17926 9276 17978
rect 9300 17926 9310 17978
rect 9310 17926 9356 17978
rect 9380 17926 9426 17978
rect 9426 17926 9436 17978
rect 9460 17926 9490 17978
rect 9490 17926 9516 17978
rect 9220 17924 9276 17926
rect 9300 17924 9356 17926
rect 9380 17924 9436 17926
rect 9460 17924 9516 17926
rect 9220 16890 9276 16892
rect 9300 16890 9356 16892
rect 9380 16890 9436 16892
rect 9460 16890 9516 16892
rect 9220 16838 9246 16890
rect 9246 16838 9276 16890
rect 9300 16838 9310 16890
rect 9310 16838 9356 16890
rect 9380 16838 9426 16890
rect 9426 16838 9436 16890
rect 9460 16838 9490 16890
rect 9490 16838 9516 16890
rect 9220 16836 9276 16838
rect 9300 16836 9356 16838
rect 9380 16836 9436 16838
rect 9460 16836 9516 16838
rect 9220 15802 9276 15804
rect 9300 15802 9356 15804
rect 9380 15802 9436 15804
rect 9460 15802 9516 15804
rect 9220 15750 9246 15802
rect 9246 15750 9276 15802
rect 9300 15750 9310 15802
rect 9310 15750 9356 15802
rect 9380 15750 9426 15802
rect 9426 15750 9436 15802
rect 9460 15750 9490 15802
rect 9490 15750 9516 15802
rect 9220 15748 9276 15750
rect 9300 15748 9356 15750
rect 9380 15748 9436 15750
rect 9460 15748 9516 15750
rect 9220 14714 9276 14716
rect 9300 14714 9356 14716
rect 9380 14714 9436 14716
rect 9460 14714 9516 14716
rect 9220 14662 9246 14714
rect 9246 14662 9276 14714
rect 9300 14662 9310 14714
rect 9310 14662 9356 14714
rect 9380 14662 9426 14714
rect 9426 14662 9436 14714
rect 9460 14662 9490 14714
rect 9490 14662 9516 14714
rect 9220 14660 9276 14662
rect 9300 14660 9356 14662
rect 9380 14660 9436 14662
rect 9460 14660 9516 14662
rect 9220 13626 9276 13628
rect 9300 13626 9356 13628
rect 9380 13626 9436 13628
rect 9460 13626 9516 13628
rect 9220 13574 9246 13626
rect 9246 13574 9276 13626
rect 9300 13574 9310 13626
rect 9310 13574 9356 13626
rect 9380 13574 9426 13626
rect 9426 13574 9436 13626
rect 9460 13574 9490 13626
rect 9490 13574 9516 13626
rect 9220 13572 9276 13574
rect 9300 13572 9356 13574
rect 9380 13572 9436 13574
rect 9460 13572 9516 13574
rect 9220 12538 9276 12540
rect 9300 12538 9356 12540
rect 9380 12538 9436 12540
rect 9460 12538 9516 12540
rect 9220 12486 9246 12538
rect 9246 12486 9276 12538
rect 9300 12486 9310 12538
rect 9310 12486 9356 12538
rect 9380 12486 9426 12538
rect 9426 12486 9436 12538
rect 9460 12486 9490 12538
rect 9490 12486 9516 12538
rect 9220 12484 9276 12486
rect 9300 12484 9356 12486
rect 9380 12484 9436 12486
rect 9460 12484 9516 12486
rect 9220 11450 9276 11452
rect 9300 11450 9356 11452
rect 9380 11450 9436 11452
rect 9460 11450 9516 11452
rect 9220 11398 9246 11450
rect 9246 11398 9276 11450
rect 9300 11398 9310 11450
rect 9310 11398 9356 11450
rect 9380 11398 9426 11450
rect 9426 11398 9436 11450
rect 9460 11398 9490 11450
rect 9490 11398 9516 11450
rect 9220 11396 9276 11398
rect 9300 11396 9356 11398
rect 9380 11396 9436 11398
rect 9460 11396 9516 11398
rect 9678 11212 9734 11248
rect 9678 11192 9680 11212
rect 9680 11192 9732 11212
rect 9732 11192 9734 11212
rect 9954 10648 10010 10704
rect 9220 10362 9276 10364
rect 9300 10362 9356 10364
rect 9380 10362 9436 10364
rect 9460 10362 9516 10364
rect 9220 10310 9246 10362
rect 9246 10310 9276 10362
rect 9300 10310 9310 10362
rect 9310 10310 9356 10362
rect 9380 10310 9426 10362
rect 9426 10310 9436 10362
rect 9460 10310 9490 10362
rect 9490 10310 9516 10362
rect 9220 10308 9276 10310
rect 9300 10308 9356 10310
rect 9380 10308 9436 10310
rect 9460 10308 9516 10310
rect 9220 9274 9276 9276
rect 9300 9274 9356 9276
rect 9380 9274 9436 9276
rect 9460 9274 9516 9276
rect 9220 9222 9246 9274
rect 9246 9222 9276 9274
rect 9300 9222 9310 9274
rect 9310 9222 9356 9274
rect 9380 9222 9426 9274
rect 9426 9222 9436 9274
rect 9460 9222 9490 9274
rect 9490 9222 9516 9274
rect 9220 9220 9276 9222
rect 9300 9220 9356 9222
rect 9380 9220 9436 9222
rect 9460 9220 9516 9222
rect 9220 8186 9276 8188
rect 9300 8186 9356 8188
rect 9380 8186 9436 8188
rect 9460 8186 9516 8188
rect 9220 8134 9246 8186
rect 9246 8134 9276 8186
rect 9300 8134 9310 8186
rect 9310 8134 9356 8186
rect 9380 8134 9426 8186
rect 9426 8134 9436 8186
rect 9460 8134 9490 8186
rect 9490 8134 9516 8186
rect 9220 8132 9276 8134
rect 9300 8132 9356 8134
rect 9380 8132 9436 8134
rect 9460 8132 9516 8134
rect 9220 7098 9276 7100
rect 9300 7098 9356 7100
rect 9380 7098 9436 7100
rect 9460 7098 9516 7100
rect 9220 7046 9246 7098
rect 9246 7046 9276 7098
rect 9300 7046 9310 7098
rect 9310 7046 9356 7098
rect 9380 7046 9426 7098
rect 9426 7046 9436 7098
rect 9460 7046 9490 7098
rect 9490 7046 9516 7098
rect 9220 7044 9276 7046
rect 9300 7044 9356 7046
rect 9380 7044 9436 7046
rect 9460 7044 9516 7046
rect 8942 3848 8998 3904
rect 9220 6010 9276 6012
rect 9300 6010 9356 6012
rect 9380 6010 9436 6012
rect 9460 6010 9516 6012
rect 9220 5958 9246 6010
rect 9246 5958 9276 6010
rect 9300 5958 9310 6010
rect 9310 5958 9356 6010
rect 9380 5958 9426 6010
rect 9426 5958 9436 6010
rect 9460 5958 9490 6010
rect 9490 5958 9516 6010
rect 9220 5956 9276 5958
rect 9300 5956 9356 5958
rect 9380 5956 9436 5958
rect 9460 5956 9516 5958
rect 9220 4922 9276 4924
rect 9300 4922 9356 4924
rect 9380 4922 9436 4924
rect 9460 4922 9516 4924
rect 9220 4870 9246 4922
rect 9246 4870 9276 4922
rect 9300 4870 9310 4922
rect 9310 4870 9356 4922
rect 9380 4870 9426 4922
rect 9426 4870 9436 4922
rect 9460 4870 9490 4922
rect 9490 4870 9516 4922
rect 9220 4868 9276 4870
rect 9300 4868 9356 4870
rect 9380 4868 9436 4870
rect 9460 4868 9516 4870
rect 9218 3984 9274 4040
rect 9220 3834 9276 3836
rect 9300 3834 9356 3836
rect 9380 3834 9436 3836
rect 9460 3834 9516 3836
rect 9220 3782 9246 3834
rect 9246 3782 9276 3834
rect 9300 3782 9310 3834
rect 9310 3782 9356 3834
rect 9380 3782 9426 3834
rect 9426 3782 9436 3834
rect 9460 3782 9490 3834
rect 9490 3782 9516 3834
rect 9220 3780 9276 3782
rect 9300 3780 9356 3782
rect 9380 3780 9436 3782
rect 9460 3780 9516 3782
rect 9220 2746 9276 2748
rect 9300 2746 9356 2748
rect 9380 2746 9436 2748
rect 9460 2746 9516 2748
rect 9220 2694 9246 2746
rect 9246 2694 9276 2746
rect 9300 2694 9310 2746
rect 9310 2694 9356 2746
rect 9380 2694 9426 2746
rect 9426 2694 9436 2746
rect 9460 2694 9490 2746
rect 9490 2694 9516 2746
rect 9220 2692 9276 2694
rect 9300 2692 9356 2694
rect 9380 2692 9436 2694
rect 9460 2692 9516 2694
rect 9770 3712 9826 3768
rect 9862 3440 9918 3496
rect 9770 2760 9826 2816
rect 10046 3576 10102 3632
rect 10506 3576 10562 3632
rect 11058 3848 11114 3904
rect 11610 10004 11612 10024
rect 11612 10004 11664 10024
rect 11664 10004 11666 10024
rect 11610 9968 11666 10004
rect 11426 7384 11482 7440
rect 11518 3712 11574 3768
rect 13358 12588 13360 12608
rect 13360 12588 13412 12608
rect 13412 12588 13414 12608
rect 13358 12552 13414 12588
rect 14220 66394 14276 66396
rect 14300 66394 14356 66396
rect 14380 66394 14436 66396
rect 14460 66394 14516 66396
rect 14220 66342 14246 66394
rect 14246 66342 14276 66394
rect 14300 66342 14310 66394
rect 14310 66342 14356 66394
rect 14380 66342 14426 66394
rect 14426 66342 14436 66394
rect 14460 66342 14490 66394
rect 14490 66342 14516 66394
rect 14220 66340 14276 66342
rect 14300 66340 14356 66342
rect 14380 66340 14436 66342
rect 14460 66340 14516 66342
rect 14220 65306 14276 65308
rect 14300 65306 14356 65308
rect 14380 65306 14436 65308
rect 14460 65306 14516 65308
rect 14220 65254 14246 65306
rect 14246 65254 14276 65306
rect 14300 65254 14310 65306
rect 14310 65254 14356 65306
rect 14380 65254 14426 65306
rect 14426 65254 14436 65306
rect 14460 65254 14490 65306
rect 14490 65254 14516 65306
rect 14220 65252 14276 65254
rect 14300 65252 14356 65254
rect 14380 65252 14436 65254
rect 14460 65252 14516 65254
rect 14220 64218 14276 64220
rect 14300 64218 14356 64220
rect 14380 64218 14436 64220
rect 14460 64218 14516 64220
rect 14220 64166 14246 64218
rect 14246 64166 14276 64218
rect 14300 64166 14310 64218
rect 14310 64166 14356 64218
rect 14380 64166 14426 64218
rect 14426 64166 14436 64218
rect 14460 64166 14490 64218
rect 14490 64166 14516 64218
rect 14220 64164 14276 64166
rect 14300 64164 14356 64166
rect 14380 64164 14436 64166
rect 14460 64164 14516 64166
rect 13542 13132 13544 13152
rect 13544 13132 13596 13152
rect 13596 13132 13598 13152
rect 13542 13096 13598 13132
rect 12254 8472 12310 8528
rect 12162 6840 12218 6896
rect 12070 3712 12126 3768
rect 12254 4004 12310 4040
rect 12254 3984 12256 4004
rect 12256 3984 12308 4004
rect 12308 3984 12310 4004
rect 12438 3712 12494 3768
rect 14220 63130 14276 63132
rect 14300 63130 14356 63132
rect 14380 63130 14436 63132
rect 14460 63130 14516 63132
rect 14220 63078 14246 63130
rect 14246 63078 14276 63130
rect 14300 63078 14310 63130
rect 14310 63078 14356 63130
rect 14380 63078 14426 63130
rect 14426 63078 14436 63130
rect 14460 63078 14490 63130
rect 14490 63078 14516 63130
rect 14220 63076 14276 63078
rect 14300 63076 14356 63078
rect 14380 63076 14436 63078
rect 14460 63076 14516 63078
rect 14220 62042 14276 62044
rect 14300 62042 14356 62044
rect 14380 62042 14436 62044
rect 14460 62042 14516 62044
rect 14220 61990 14246 62042
rect 14246 61990 14276 62042
rect 14300 61990 14310 62042
rect 14310 61990 14356 62042
rect 14380 61990 14426 62042
rect 14426 61990 14436 62042
rect 14460 61990 14490 62042
rect 14490 61990 14516 62042
rect 14220 61988 14276 61990
rect 14300 61988 14356 61990
rect 14380 61988 14436 61990
rect 14460 61988 14516 61990
rect 14220 60954 14276 60956
rect 14300 60954 14356 60956
rect 14380 60954 14436 60956
rect 14460 60954 14516 60956
rect 14220 60902 14246 60954
rect 14246 60902 14276 60954
rect 14300 60902 14310 60954
rect 14310 60902 14356 60954
rect 14380 60902 14426 60954
rect 14426 60902 14436 60954
rect 14460 60902 14490 60954
rect 14490 60902 14516 60954
rect 14220 60900 14276 60902
rect 14300 60900 14356 60902
rect 14380 60900 14436 60902
rect 14460 60900 14516 60902
rect 14220 59866 14276 59868
rect 14300 59866 14356 59868
rect 14380 59866 14436 59868
rect 14460 59866 14516 59868
rect 14220 59814 14246 59866
rect 14246 59814 14276 59866
rect 14300 59814 14310 59866
rect 14310 59814 14356 59866
rect 14380 59814 14426 59866
rect 14426 59814 14436 59866
rect 14460 59814 14490 59866
rect 14490 59814 14516 59866
rect 14220 59812 14276 59814
rect 14300 59812 14356 59814
rect 14380 59812 14436 59814
rect 14460 59812 14516 59814
rect 14220 58778 14276 58780
rect 14300 58778 14356 58780
rect 14380 58778 14436 58780
rect 14460 58778 14516 58780
rect 14220 58726 14246 58778
rect 14246 58726 14276 58778
rect 14300 58726 14310 58778
rect 14310 58726 14356 58778
rect 14380 58726 14426 58778
rect 14426 58726 14436 58778
rect 14460 58726 14490 58778
rect 14490 58726 14516 58778
rect 14220 58724 14276 58726
rect 14300 58724 14356 58726
rect 14380 58724 14436 58726
rect 14460 58724 14516 58726
rect 14220 57690 14276 57692
rect 14300 57690 14356 57692
rect 14380 57690 14436 57692
rect 14460 57690 14516 57692
rect 14220 57638 14246 57690
rect 14246 57638 14276 57690
rect 14300 57638 14310 57690
rect 14310 57638 14356 57690
rect 14380 57638 14426 57690
rect 14426 57638 14436 57690
rect 14460 57638 14490 57690
rect 14490 57638 14516 57690
rect 14220 57636 14276 57638
rect 14300 57636 14356 57638
rect 14380 57636 14436 57638
rect 14460 57636 14516 57638
rect 14220 56602 14276 56604
rect 14300 56602 14356 56604
rect 14380 56602 14436 56604
rect 14460 56602 14516 56604
rect 14220 56550 14246 56602
rect 14246 56550 14276 56602
rect 14300 56550 14310 56602
rect 14310 56550 14356 56602
rect 14380 56550 14426 56602
rect 14426 56550 14436 56602
rect 14460 56550 14490 56602
rect 14490 56550 14516 56602
rect 14220 56548 14276 56550
rect 14300 56548 14356 56550
rect 14380 56548 14436 56550
rect 14460 56548 14516 56550
rect 14220 55514 14276 55516
rect 14300 55514 14356 55516
rect 14380 55514 14436 55516
rect 14460 55514 14516 55516
rect 14220 55462 14246 55514
rect 14246 55462 14276 55514
rect 14300 55462 14310 55514
rect 14310 55462 14356 55514
rect 14380 55462 14426 55514
rect 14426 55462 14436 55514
rect 14460 55462 14490 55514
rect 14490 55462 14516 55514
rect 14220 55460 14276 55462
rect 14300 55460 14356 55462
rect 14380 55460 14436 55462
rect 14460 55460 14516 55462
rect 14220 54426 14276 54428
rect 14300 54426 14356 54428
rect 14380 54426 14436 54428
rect 14460 54426 14516 54428
rect 14220 54374 14246 54426
rect 14246 54374 14276 54426
rect 14300 54374 14310 54426
rect 14310 54374 14356 54426
rect 14380 54374 14426 54426
rect 14426 54374 14436 54426
rect 14460 54374 14490 54426
rect 14490 54374 14516 54426
rect 14220 54372 14276 54374
rect 14300 54372 14356 54374
rect 14380 54372 14436 54374
rect 14460 54372 14516 54374
rect 14220 53338 14276 53340
rect 14300 53338 14356 53340
rect 14380 53338 14436 53340
rect 14460 53338 14516 53340
rect 14220 53286 14246 53338
rect 14246 53286 14276 53338
rect 14300 53286 14310 53338
rect 14310 53286 14356 53338
rect 14380 53286 14426 53338
rect 14426 53286 14436 53338
rect 14460 53286 14490 53338
rect 14490 53286 14516 53338
rect 14220 53284 14276 53286
rect 14300 53284 14356 53286
rect 14380 53284 14436 53286
rect 14460 53284 14516 53286
rect 14220 52250 14276 52252
rect 14300 52250 14356 52252
rect 14380 52250 14436 52252
rect 14460 52250 14516 52252
rect 14220 52198 14246 52250
rect 14246 52198 14276 52250
rect 14300 52198 14310 52250
rect 14310 52198 14356 52250
rect 14380 52198 14426 52250
rect 14426 52198 14436 52250
rect 14460 52198 14490 52250
rect 14490 52198 14516 52250
rect 14220 52196 14276 52198
rect 14300 52196 14356 52198
rect 14380 52196 14436 52198
rect 14460 52196 14516 52198
rect 14220 51162 14276 51164
rect 14300 51162 14356 51164
rect 14380 51162 14436 51164
rect 14460 51162 14516 51164
rect 14220 51110 14246 51162
rect 14246 51110 14276 51162
rect 14300 51110 14310 51162
rect 14310 51110 14356 51162
rect 14380 51110 14426 51162
rect 14426 51110 14436 51162
rect 14460 51110 14490 51162
rect 14490 51110 14516 51162
rect 14220 51108 14276 51110
rect 14300 51108 14356 51110
rect 14380 51108 14436 51110
rect 14460 51108 14516 51110
rect 14220 50074 14276 50076
rect 14300 50074 14356 50076
rect 14380 50074 14436 50076
rect 14460 50074 14516 50076
rect 14220 50022 14246 50074
rect 14246 50022 14276 50074
rect 14300 50022 14310 50074
rect 14310 50022 14356 50074
rect 14380 50022 14426 50074
rect 14426 50022 14436 50074
rect 14460 50022 14490 50074
rect 14490 50022 14516 50074
rect 14220 50020 14276 50022
rect 14300 50020 14356 50022
rect 14380 50020 14436 50022
rect 14460 50020 14516 50022
rect 14220 48986 14276 48988
rect 14300 48986 14356 48988
rect 14380 48986 14436 48988
rect 14460 48986 14516 48988
rect 14220 48934 14246 48986
rect 14246 48934 14276 48986
rect 14300 48934 14310 48986
rect 14310 48934 14356 48986
rect 14380 48934 14426 48986
rect 14426 48934 14436 48986
rect 14460 48934 14490 48986
rect 14490 48934 14516 48986
rect 14220 48932 14276 48934
rect 14300 48932 14356 48934
rect 14380 48932 14436 48934
rect 14460 48932 14516 48934
rect 14220 47898 14276 47900
rect 14300 47898 14356 47900
rect 14380 47898 14436 47900
rect 14460 47898 14516 47900
rect 14220 47846 14246 47898
rect 14246 47846 14276 47898
rect 14300 47846 14310 47898
rect 14310 47846 14356 47898
rect 14380 47846 14426 47898
rect 14426 47846 14436 47898
rect 14460 47846 14490 47898
rect 14490 47846 14516 47898
rect 14220 47844 14276 47846
rect 14300 47844 14356 47846
rect 14380 47844 14436 47846
rect 14460 47844 14516 47846
rect 14220 46810 14276 46812
rect 14300 46810 14356 46812
rect 14380 46810 14436 46812
rect 14460 46810 14516 46812
rect 14220 46758 14246 46810
rect 14246 46758 14276 46810
rect 14300 46758 14310 46810
rect 14310 46758 14356 46810
rect 14380 46758 14426 46810
rect 14426 46758 14436 46810
rect 14460 46758 14490 46810
rect 14490 46758 14516 46810
rect 14220 46756 14276 46758
rect 14300 46756 14356 46758
rect 14380 46756 14436 46758
rect 14460 46756 14516 46758
rect 14220 45722 14276 45724
rect 14300 45722 14356 45724
rect 14380 45722 14436 45724
rect 14460 45722 14516 45724
rect 14220 45670 14246 45722
rect 14246 45670 14276 45722
rect 14300 45670 14310 45722
rect 14310 45670 14356 45722
rect 14380 45670 14426 45722
rect 14426 45670 14436 45722
rect 14460 45670 14490 45722
rect 14490 45670 14516 45722
rect 14220 45668 14276 45670
rect 14300 45668 14356 45670
rect 14380 45668 14436 45670
rect 14460 45668 14516 45670
rect 14220 44634 14276 44636
rect 14300 44634 14356 44636
rect 14380 44634 14436 44636
rect 14460 44634 14516 44636
rect 14220 44582 14246 44634
rect 14246 44582 14276 44634
rect 14300 44582 14310 44634
rect 14310 44582 14356 44634
rect 14380 44582 14426 44634
rect 14426 44582 14436 44634
rect 14460 44582 14490 44634
rect 14490 44582 14516 44634
rect 14220 44580 14276 44582
rect 14300 44580 14356 44582
rect 14380 44580 14436 44582
rect 14460 44580 14516 44582
rect 14220 43546 14276 43548
rect 14300 43546 14356 43548
rect 14380 43546 14436 43548
rect 14460 43546 14516 43548
rect 14220 43494 14246 43546
rect 14246 43494 14276 43546
rect 14300 43494 14310 43546
rect 14310 43494 14356 43546
rect 14380 43494 14426 43546
rect 14426 43494 14436 43546
rect 14460 43494 14490 43546
rect 14490 43494 14516 43546
rect 14220 43492 14276 43494
rect 14300 43492 14356 43494
rect 14380 43492 14436 43494
rect 14460 43492 14516 43494
rect 14220 42458 14276 42460
rect 14300 42458 14356 42460
rect 14380 42458 14436 42460
rect 14460 42458 14516 42460
rect 14220 42406 14246 42458
rect 14246 42406 14276 42458
rect 14300 42406 14310 42458
rect 14310 42406 14356 42458
rect 14380 42406 14426 42458
rect 14426 42406 14436 42458
rect 14460 42406 14490 42458
rect 14490 42406 14516 42458
rect 14220 42404 14276 42406
rect 14300 42404 14356 42406
rect 14380 42404 14436 42406
rect 14460 42404 14516 42406
rect 14220 41370 14276 41372
rect 14300 41370 14356 41372
rect 14380 41370 14436 41372
rect 14460 41370 14516 41372
rect 14220 41318 14246 41370
rect 14246 41318 14276 41370
rect 14300 41318 14310 41370
rect 14310 41318 14356 41370
rect 14380 41318 14426 41370
rect 14426 41318 14436 41370
rect 14460 41318 14490 41370
rect 14490 41318 14516 41370
rect 14220 41316 14276 41318
rect 14300 41316 14356 41318
rect 14380 41316 14436 41318
rect 14460 41316 14516 41318
rect 14220 40282 14276 40284
rect 14300 40282 14356 40284
rect 14380 40282 14436 40284
rect 14460 40282 14516 40284
rect 14220 40230 14246 40282
rect 14246 40230 14276 40282
rect 14300 40230 14310 40282
rect 14310 40230 14356 40282
rect 14380 40230 14426 40282
rect 14426 40230 14436 40282
rect 14460 40230 14490 40282
rect 14490 40230 14516 40282
rect 14220 40228 14276 40230
rect 14300 40228 14356 40230
rect 14380 40228 14436 40230
rect 14460 40228 14516 40230
rect 14220 39194 14276 39196
rect 14300 39194 14356 39196
rect 14380 39194 14436 39196
rect 14460 39194 14516 39196
rect 14220 39142 14246 39194
rect 14246 39142 14276 39194
rect 14300 39142 14310 39194
rect 14310 39142 14356 39194
rect 14380 39142 14426 39194
rect 14426 39142 14436 39194
rect 14460 39142 14490 39194
rect 14490 39142 14516 39194
rect 14220 39140 14276 39142
rect 14300 39140 14356 39142
rect 14380 39140 14436 39142
rect 14460 39140 14516 39142
rect 14220 38106 14276 38108
rect 14300 38106 14356 38108
rect 14380 38106 14436 38108
rect 14460 38106 14516 38108
rect 14220 38054 14246 38106
rect 14246 38054 14276 38106
rect 14300 38054 14310 38106
rect 14310 38054 14356 38106
rect 14380 38054 14426 38106
rect 14426 38054 14436 38106
rect 14460 38054 14490 38106
rect 14490 38054 14516 38106
rect 14220 38052 14276 38054
rect 14300 38052 14356 38054
rect 14380 38052 14436 38054
rect 14460 38052 14516 38054
rect 14220 37018 14276 37020
rect 14300 37018 14356 37020
rect 14380 37018 14436 37020
rect 14460 37018 14516 37020
rect 14220 36966 14246 37018
rect 14246 36966 14276 37018
rect 14300 36966 14310 37018
rect 14310 36966 14356 37018
rect 14380 36966 14426 37018
rect 14426 36966 14436 37018
rect 14460 36966 14490 37018
rect 14490 36966 14516 37018
rect 14220 36964 14276 36966
rect 14300 36964 14356 36966
rect 14380 36964 14436 36966
rect 14460 36964 14516 36966
rect 14220 35930 14276 35932
rect 14300 35930 14356 35932
rect 14380 35930 14436 35932
rect 14460 35930 14516 35932
rect 14220 35878 14246 35930
rect 14246 35878 14276 35930
rect 14300 35878 14310 35930
rect 14310 35878 14356 35930
rect 14380 35878 14426 35930
rect 14426 35878 14436 35930
rect 14460 35878 14490 35930
rect 14490 35878 14516 35930
rect 14220 35876 14276 35878
rect 14300 35876 14356 35878
rect 14380 35876 14436 35878
rect 14460 35876 14516 35878
rect 14220 34842 14276 34844
rect 14300 34842 14356 34844
rect 14380 34842 14436 34844
rect 14460 34842 14516 34844
rect 14220 34790 14246 34842
rect 14246 34790 14276 34842
rect 14300 34790 14310 34842
rect 14310 34790 14356 34842
rect 14380 34790 14426 34842
rect 14426 34790 14436 34842
rect 14460 34790 14490 34842
rect 14490 34790 14516 34842
rect 14220 34788 14276 34790
rect 14300 34788 14356 34790
rect 14380 34788 14436 34790
rect 14460 34788 14516 34790
rect 14220 33754 14276 33756
rect 14300 33754 14356 33756
rect 14380 33754 14436 33756
rect 14460 33754 14516 33756
rect 14220 33702 14246 33754
rect 14246 33702 14276 33754
rect 14300 33702 14310 33754
rect 14310 33702 14356 33754
rect 14380 33702 14426 33754
rect 14426 33702 14436 33754
rect 14460 33702 14490 33754
rect 14490 33702 14516 33754
rect 14220 33700 14276 33702
rect 14300 33700 14356 33702
rect 14380 33700 14436 33702
rect 14460 33700 14516 33702
rect 14220 32666 14276 32668
rect 14300 32666 14356 32668
rect 14380 32666 14436 32668
rect 14460 32666 14516 32668
rect 14220 32614 14246 32666
rect 14246 32614 14276 32666
rect 14300 32614 14310 32666
rect 14310 32614 14356 32666
rect 14380 32614 14426 32666
rect 14426 32614 14436 32666
rect 14460 32614 14490 32666
rect 14490 32614 14516 32666
rect 14220 32612 14276 32614
rect 14300 32612 14356 32614
rect 14380 32612 14436 32614
rect 14460 32612 14516 32614
rect 14220 31578 14276 31580
rect 14300 31578 14356 31580
rect 14380 31578 14436 31580
rect 14460 31578 14516 31580
rect 14220 31526 14246 31578
rect 14246 31526 14276 31578
rect 14300 31526 14310 31578
rect 14310 31526 14356 31578
rect 14380 31526 14426 31578
rect 14426 31526 14436 31578
rect 14460 31526 14490 31578
rect 14490 31526 14516 31578
rect 14220 31524 14276 31526
rect 14300 31524 14356 31526
rect 14380 31524 14436 31526
rect 14460 31524 14516 31526
rect 14220 30490 14276 30492
rect 14300 30490 14356 30492
rect 14380 30490 14436 30492
rect 14460 30490 14516 30492
rect 14220 30438 14246 30490
rect 14246 30438 14276 30490
rect 14300 30438 14310 30490
rect 14310 30438 14356 30490
rect 14380 30438 14426 30490
rect 14426 30438 14436 30490
rect 14460 30438 14490 30490
rect 14490 30438 14516 30490
rect 14220 30436 14276 30438
rect 14300 30436 14356 30438
rect 14380 30436 14436 30438
rect 14460 30436 14516 30438
rect 14220 29402 14276 29404
rect 14300 29402 14356 29404
rect 14380 29402 14436 29404
rect 14460 29402 14516 29404
rect 14220 29350 14246 29402
rect 14246 29350 14276 29402
rect 14300 29350 14310 29402
rect 14310 29350 14356 29402
rect 14380 29350 14426 29402
rect 14426 29350 14436 29402
rect 14460 29350 14490 29402
rect 14490 29350 14516 29402
rect 14220 29348 14276 29350
rect 14300 29348 14356 29350
rect 14380 29348 14436 29350
rect 14460 29348 14516 29350
rect 14220 28314 14276 28316
rect 14300 28314 14356 28316
rect 14380 28314 14436 28316
rect 14460 28314 14516 28316
rect 14220 28262 14246 28314
rect 14246 28262 14276 28314
rect 14300 28262 14310 28314
rect 14310 28262 14356 28314
rect 14380 28262 14426 28314
rect 14426 28262 14436 28314
rect 14460 28262 14490 28314
rect 14490 28262 14516 28314
rect 14220 28260 14276 28262
rect 14300 28260 14356 28262
rect 14380 28260 14436 28262
rect 14460 28260 14516 28262
rect 14220 27226 14276 27228
rect 14300 27226 14356 27228
rect 14380 27226 14436 27228
rect 14460 27226 14516 27228
rect 14220 27174 14246 27226
rect 14246 27174 14276 27226
rect 14300 27174 14310 27226
rect 14310 27174 14356 27226
rect 14380 27174 14426 27226
rect 14426 27174 14436 27226
rect 14460 27174 14490 27226
rect 14490 27174 14516 27226
rect 14220 27172 14276 27174
rect 14300 27172 14356 27174
rect 14380 27172 14436 27174
rect 14460 27172 14516 27174
rect 14220 26138 14276 26140
rect 14300 26138 14356 26140
rect 14380 26138 14436 26140
rect 14460 26138 14516 26140
rect 14220 26086 14246 26138
rect 14246 26086 14276 26138
rect 14300 26086 14310 26138
rect 14310 26086 14356 26138
rect 14380 26086 14426 26138
rect 14426 26086 14436 26138
rect 14460 26086 14490 26138
rect 14490 26086 14516 26138
rect 14220 26084 14276 26086
rect 14300 26084 14356 26086
rect 14380 26084 14436 26086
rect 14460 26084 14516 26086
rect 14220 25050 14276 25052
rect 14300 25050 14356 25052
rect 14380 25050 14436 25052
rect 14460 25050 14516 25052
rect 14220 24998 14246 25050
rect 14246 24998 14276 25050
rect 14300 24998 14310 25050
rect 14310 24998 14356 25050
rect 14380 24998 14426 25050
rect 14426 24998 14436 25050
rect 14460 24998 14490 25050
rect 14490 24998 14516 25050
rect 14220 24996 14276 24998
rect 14300 24996 14356 24998
rect 14380 24996 14436 24998
rect 14460 24996 14516 24998
rect 14220 23962 14276 23964
rect 14300 23962 14356 23964
rect 14380 23962 14436 23964
rect 14460 23962 14516 23964
rect 14220 23910 14246 23962
rect 14246 23910 14276 23962
rect 14300 23910 14310 23962
rect 14310 23910 14356 23962
rect 14380 23910 14426 23962
rect 14426 23910 14436 23962
rect 14460 23910 14490 23962
rect 14490 23910 14516 23962
rect 14220 23908 14276 23910
rect 14300 23908 14356 23910
rect 14380 23908 14436 23910
rect 14460 23908 14516 23910
rect 14220 22874 14276 22876
rect 14300 22874 14356 22876
rect 14380 22874 14436 22876
rect 14460 22874 14516 22876
rect 14220 22822 14246 22874
rect 14246 22822 14276 22874
rect 14300 22822 14310 22874
rect 14310 22822 14356 22874
rect 14380 22822 14426 22874
rect 14426 22822 14436 22874
rect 14460 22822 14490 22874
rect 14490 22822 14516 22874
rect 14220 22820 14276 22822
rect 14300 22820 14356 22822
rect 14380 22820 14436 22822
rect 14460 22820 14516 22822
rect 14220 21786 14276 21788
rect 14300 21786 14356 21788
rect 14380 21786 14436 21788
rect 14460 21786 14516 21788
rect 14220 21734 14246 21786
rect 14246 21734 14276 21786
rect 14300 21734 14310 21786
rect 14310 21734 14356 21786
rect 14380 21734 14426 21786
rect 14426 21734 14436 21786
rect 14460 21734 14490 21786
rect 14490 21734 14516 21786
rect 14220 21732 14276 21734
rect 14300 21732 14356 21734
rect 14380 21732 14436 21734
rect 14460 21732 14516 21734
rect 14220 20698 14276 20700
rect 14300 20698 14356 20700
rect 14380 20698 14436 20700
rect 14460 20698 14516 20700
rect 14220 20646 14246 20698
rect 14246 20646 14276 20698
rect 14300 20646 14310 20698
rect 14310 20646 14356 20698
rect 14380 20646 14426 20698
rect 14426 20646 14436 20698
rect 14460 20646 14490 20698
rect 14490 20646 14516 20698
rect 14220 20644 14276 20646
rect 14300 20644 14356 20646
rect 14380 20644 14436 20646
rect 14460 20644 14516 20646
rect 14220 19610 14276 19612
rect 14300 19610 14356 19612
rect 14380 19610 14436 19612
rect 14460 19610 14516 19612
rect 14220 19558 14246 19610
rect 14246 19558 14276 19610
rect 14300 19558 14310 19610
rect 14310 19558 14356 19610
rect 14380 19558 14426 19610
rect 14426 19558 14436 19610
rect 14460 19558 14490 19610
rect 14490 19558 14516 19610
rect 14220 19556 14276 19558
rect 14300 19556 14356 19558
rect 14380 19556 14436 19558
rect 14460 19556 14516 19558
rect 14220 18522 14276 18524
rect 14300 18522 14356 18524
rect 14380 18522 14436 18524
rect 14460 18522 14516 18524
rect 14220 18470 14246 18522
rect 14246 18470 14276 18522
rect 14300 18470 14310 18522
rect 14310 18470 14356 18522
rect 14380 18470 14426 18522
rect 14426 18470 14436 18522
rect 14460 18470 14490 18522
rect 14490 18470 14516 18522
rect 14220 18468 14276 18470
rect 14300 18468 14356 18470
rect 14380 18468 14436 18470
rect 14460 18468 14516 18470
rect 14220 17434 14276 17436
rect 14300 17434 14356 17436
rect 14380 17434 14436 17436
rect 14460 17434 14516 17436
rect 14220 17382 14246 17434
rect 14246 17382 14276 17434
rect 14300 17382 14310 17434
rect 14310 17382 14356 17434
rect 14380 17382 14426 17434
rect 14426 17382 14436 17434
rect 14460 17382 14490 17434
rect 14490 17382 14516 17434
rect 14220 17380 14276 17382
rect 14300 17380 14356 17382
rect 14380 17380 14436 17382
rect 14460 17380 14516 17382
rect 14220 16346 14276 16348
rect 14300 16346 14356 16348
rect 14380 16346 14436 16348
rect 14460 16346 14516 16348
rect 14220 16294 14246 16346
rect 14246 16294 14276 16346
rect 14300 16294 14310 16346
rect 14310 16294 14356 16346
rect 14380 16294 14426 16346
rect 14426 16294 14436 16346
rect 14460 16294 14490 16346
rect 14490 16294 14516 16346
rect 14220 16292 14276 16294
rect 14300 16292 14356 16294
rect 14380 16292 14436 16294
rect 14460 16292 14516 16294
rect 14220 15258 14276 15260
rect 14300 15258 14356 15260
rect 14380 15258 14436 15260
rect 14460 15258 14516 15260
rect 14220 15206 14246 15258
rect 14246 15206 14276 15258
rect 14300 15206 14310 15258
rect 14310 15206 14356 15258
rect 14380 15206 14426 15258
rect 14426 15206 14436 15258
rect 14460 15206 14490 15258
rect 14490 15206 14516 15258
rect 14220 15204 14276 15206
rect 14300 15204 14356 15206
rect 14380 15204 14436 15206
rect 14460 15204 14516 15206
rect 14220 14170 14276 14172
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14220 14118 14246 14170
rect 14246 14118 14276 14170
rect 14300 14118 14310 14170
rect 14310 14118 14356 14170
rect 14380 14118 14426 14170
rect 14426 14118 14436 14170
rect 14460 14118 14490 14170
rect 14490 14118 14516 14170
rect 14220 14116 14276 14118
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14220 13082 14276 13084
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14220 13030 14246 13082
rect 14246 13030 14276 13082
rect 14300 13030 14310 13082
rect 14310 13030 14356 13082
rect 14380 13030 14426 13082
rect 14426 13030 14436 13082
rect 14460 13030 14490 13082
rect 14490 13030 14516 13082
rect 14220 13028 14276 13030
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 13174 5888 13230 5944
rect 13082 2624 13138 2680
rect 13910 12144 13966 12200
rect 13818 11328 13874 11384
rect 13358 3712 13414 3768
rect 13634 7656 13690 7712
rect 13634 5752 13690 5808
rect 13542 3848 13598 3904
rect 13726 2896 13782 2952
rect 14220 11994 14276 11996
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14220 11942 14246 11994
rect 14246 11942 14276 11994
rect 14300 11942 14310 11994
rect 14310 11942 14356 11994
rect 14380 11942 14426 11994
rect 14426 11942 14436 11994
rect 14460 11942 14490 11994
rect 14490 11942 14516 11994
rect 14220 11940 14276 11942
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14220 10906 14276 10908
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14220 10854 14246 10906
rect 14246 10854 14276 10906
rect 14300 10854 14310 10906
rect 14310 10854 14356 10906
rect 14380 10854 14426 10906
rect 14426 10854 14436 10906
rect 14460 10854 14490 10906
rect 14490 10854 14516 10906
rect 14220 10852 14276 10854
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14462 10512 14518 10568
rect 14554 9968 14610 10024
rect 14220 9818 14276 9820
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14220 9766 14246 9818
rect 14246 9766 14276 9818
rect 14300 9766 14310 9818
rect 14310 9766 14356 9818
rect 14380 9766 14426 9818
rect 14426 9766 14436 9818
rect 14460 9766 14490 9818
rect 14490 9766 14516 9818
rect 14220 9764 14276 9766
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14370 9632 14426 9688
rect 14094 9016 14150 9072
rect 14370 8880 14426 8936
rect 14220 8730 14276 8732
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14220 8678 14246 8730
rect 14246 8678 14276 8730
rect 14300 8678 14310 8730
rect 14310 8678 14356 8730
rect 14380 8678 14426 8730
rect 14426 8678 14436 8730
rect 14460 8678 14490 8730
rect 14490 8678 14516 8730
rect 14220 8676 14276 8678
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14220 7642 14276 7644
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14220 7590 14246 7642
rect 14246 7590 14276 7642
rect 14300 7590 14310 7642
rect 14310 7590 14356 7642
rect 14380 7590 14426 7642
rect 14426 7590 14436 7642
rect 14460 7590 14490 7642
rect 14490 7590 14516 7642
rect 14220 7588 14276 7590
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14220 6554 14276 6556
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14220 6502 14246 6554
rect 14246 6502 14276 6554
rect 14300 6502 14310 6554
rect 14310 6502 14356 6554
rect 14380 6502 14426 6554
rect 14426 6502 14436 6554
rect 14460 6502 14490 6554
rect 14490 6502 14516 6554
rect 14220 6500 14276 6502
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14462 6296 14518 6352
rect 14220 5466 14276 5468
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14220 5414 14246 5466
rect 14246 5414 14276 5466
rect 14300 5414 14310 5466
rect 14310 5414 14356 5466
rect 14380 5414 14426 5466
rect 14426 5414 14436 5466
rect 14460 5414 14490 5466
rect 14490 5414 14516 5466
rect 14220 5412 14276 5414
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14830 11600 14886 11656
rect 14830 10240 14886 10296
rect 14738 10104 14794 10160
rect 14738 9632 14794 9688
rect 14002 3848 14058 3904
rect 13818 2624 13874 2680
rect 14220 4378 14276 4380
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14220 4326 14246 4378
rect 14246 4326 14276 4378
rect 14300 4326 14310 4378
rect 14310 4326 14356 4378
rect 14380 4326 14426 4378
rect 14426 4326 14436 4378
rect 14460 4326 14490 4378
rect 14490 4326 14516 4378
rect 14220 4324 14276 4326
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14462 4004 14518 4040
rect 14462 3984 14464 4004
rect 14464 3984 14516 4004
rect 14516 3984 14518 4004
rect 14370 3848 14426 3904
rect 14220 3290 14276 3292
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14220 3238 14246 3290
rect 14246 3238 14276 3290
rect 14300 3238 14310 3290
rect 14310 3238 14356 3290
rect 14380 3238 14426 3290
rect 14426 3238 14436 3290
rect 14460 3238 14490 3290
rect 14490 3238 14516 3290
rect 14220 3236 14276 3238
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14220 2202 14276 2204
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14220 2150 14246 2202
rect 14246 2150 14276 2202
rect 14300 2150 14310 2202
rect 14310 2150 14356 2202
rect 14380 2150 14426 2202
rect 14426 2150 14436 2202
rect 14460 2150 14490 2202
rect 14490 2150 14516 2202
rect 14220 2148 14276 2150
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14922 9288 14978 9344
rect 15842 13812 15844 13832
rect 15844 13812 15896 13832
rect 15896 13812 15898 13832
rect 15842 13776 15898 13812
rect 15198 9968 15254 10024
rect 15290 6024 15346 6080
rect 15474 6024 15530 6080
rect 14922 2760 14978 2816
rect 15474 3712 15530 3768
rect 15842 6976 15898 7032
rect 15198 2624 15254 2680
rect 16302 13812 16304 13832
rect 16304 13812 16356 13832
rect 16356 13812 16358 13832
rect 16302 13776 16358 13812
rect 16118 12008 16174 12064
rect 16210 9424 16266 9480
rect 16118 6704 16174 6760
rect 16302 8336 16358 8392
rect 15934 3032 15990 3088
rect 16210 4800 16266 4856
rect 16210 3984 16266 4040
rect 16578 5652 16580 5672
rect 16580 5652 16632 5672
rect 16632 5652 16634 5672
rect 16578 5616 16634 5652
rect 16486 4120 16542 4176
rect 16210 2760 16266 2816
rect 16578 3576 16634 3632
rect 17222 9016 17278 9072
rect 17222 5208 17278 5264
rect 19220 66938 19276 66940
rect 19300 66938 19356 66940
rect 19380 66938 19436 66940
rect 19460 66938 19516 66940
rect 19220 66886 19246 66938
rect 19246 66886 19276 66938
rect 19300 66886 19310 66938
rect 19310 66886 19356 66938
rect 19380 66886 19426 66938
rect 19426 66886 19436 66938
rect 19460 66886 19490 66938
rect 19490 66886 19516 66938
rect 19220 66884 19276 66886
rect 19300 66884 19356 66886
rect 19380 66884 19436 66886
rect 19460 66884 19516 66886
rect 24220 66394 24276 66396
rect 24300 66394 24356 66396
rect 24380 66394 24436 66396
rect 24460 66394 24516 66396
rect 24220 66342 24246 66394
rect 24246 66342 24276 66394
rect 24300 66342 24310 66394
rect 24310 66342 24356 66394
rect 24380 66342 24426 66394
rect 24426 66342 24436 66394
rect 24460 66342 24490 66394
rect 24490 66342 24516 66394
rect 24220 66340 24276 66342
rect 24300 66340 24356 66342
rect 24380 66340 24436 66342
rect 24460 66340 24516 66342
rect 19220 65850 19276 65852
rect 19300 65850 19356 65852
rect 19380 65850 19436 65852
rect 19460 65850 19516 65852
rect 19220 65798 19246 65850
rect 19246 65798 19276 65850
rect 19300 65798 19310 65850
rect 19310 65798 19356 65850
rect 19380 65798 19426 65850
rect 19426 65798 19436 65850
rect 19460 65798 19490 65850
rect 19490 65798 19516 65850
rect 19220 65796 19276 65798
rect 19300 65796 19356 65798
rect 19380 65796 19436 65798
rect 19460 65796 19516 65798
rect 24220 65306 24276 65308
rect 24300 65306 24356 65308
rect 24380 65306 24436 65308
rect 24460 65306 24516 65308
rect 24220 65254 24246 65306
rect 24246 65254 24276 65306
rect 24300 65254 24310 65306
rect 24310 65254 24356 65306
rect 24380 65254 24426 65306
rect 24426 65254 24436 65306
rect 24460 65254 24490 65306
rect 24490 65254 24516 65306
rect 24220 65252 24276 65254
rect 24300 65252 24356 65254
rect 24380 65252 24436 65254
rect 24460 65252 24516 65254
rect 19220 64762 19276 64764
rect 19300 64762 19356 64764
rect 19380 64762 19436 64764
rect 19460 64762 19516 64764
rect 19220 64710 19246 64762
rect 19246 64710 19276 64762
rect 19300 64710 19310 64762
rect 19310 64710 19356 64762
rect 19380 64710 19426 64762
rect 19426 64710 19436 64762
rect 19460 64710 19490 64762
rect 19490 64710 19516 64762
rect 19220 64708 19276 64710
rect 19300 64708 19356 64710
rect 19380 64708 19436 64710
rect 19460 64708 19516 64710
rect 24220 64218 24276 64220
rect 24300 64218 24356 64220
rect 24380 64218 24436 64220
rect 24460 64218 24516 64220
rect 24220 64166 24246 64218
rect 24246 64166 24276 64218
rect 24300 64166 24310 64218
rect 24310 64166 24356 64218
rect 24380 64166 24426 64218
rect 24426 64166 24436 64218
rect 24460 64166 24490 64218
rect 24490 64166 24516 64218
rect 24220 64164 24276 64166
rect 24300 64164 24356 64166
rect 24380 64164 24436 64166
rect 24460 64164 24516 64166
rect 19220 63674 19276 63676
rect 19300 63674 19356 63676
rect 19380 63674 19436 63676
rect 19460 63674 19516 63676
rect 19220 63622 19246 63674
rect 19246 63622 19276 63674
rect 19300 63622 19310 63674
rect 19310 63622 19356 63674
rect 19380 63622 19426 63674
rect 19426 63622 19436 63674
rect 19460 63622 19490 63674
rect 19490 63622 19516 63674
rect 19220 63620 19276 63622
rect 19300 63620 19356 63622
rect 19380 63620 19436 63622
rect 19460 63620 19516 63622
rect 24220 63130 24276 63132
rect 24300 63130 24356 63132
rect 24380 63130 24436 63132
rect 24460 63130 24516 63132
rect 24220 63078 24246 63130
rect 24246 63078 24276 63130
rect 24300 63078 24310 63130
rect 24310 63078 24356 63130
rect 24380 63078 24426 63130
rect 24426 63078 24436 63130
rect 24460 63078 24490 63130
rect 24490 63078 24516 63130
rect 24220 63076 24276 63078
rect 24300 63076 24356 63078
rect 24380 63076 24436 63078
rect 24460 63076 24516 63078
rect 19220 62586 19276 62588
rect 19300 62586 19356 62588
rect 19380 62586 19436 62588
rect 19460 62586 19516 62588
rect 19220 62534 19246 62586
rect 19246 62534 19276 62586
rect 19300 62534 19310 62586
rect 19310 62534 19356 62586
rect 19380 62534 19426 62586
rect 19426 62534 19436 62586
rect 19460 62534 19490 62586
rect 19490 62534 19516 62586
rect 19220 62532 19276 62534
rect 19300 62532 19356 62534
rect 19380 62532 19436 62534
rect 19460 62532 19516 62534
rect 19220 61498 19276 61500
rect 19300 61498 19356 61500
rect 19380 61498 19436 61500
rect 19460 61498 19516 61500
rect 19220 61446 19246 61498
rect 19246 61446 19276 61498
rect 19300 61446 19310 61498
rect 19310 61446 19356 61498
rect 19380 61446 19426 61498
rect 19426 61446 19436 61498
rect 19460 61446 19490 61498
rect 19490 61446 19516 61498
rect 19220 61444 19276 61446
rect 19300 61444 19356 61446
rect 19380 61444 19436 61446
rect 19460 61444 19516 61446
rect 19220 60410 19276 60412
rect 19300 60410 19356 60412
rect 19380 60410 19436 60412
rect 19460 60410 19516 60412
rect 19220 60358 19246 60410
rect 19246 60358 19276 60410
rect 19300 60358 19310 60410
rect 19310 60358 19356 60410
rect 19380 60358 19426 60410
rect 19426 60358 19436 60410
rect 19460 60358 19490 60410
rect 19490 60358 19516 60410
rect 19220 60356 19276 60358
rect 19300 60356 19356 60358
rect 19380 60356 19436 60358
rect 19460 60356 19516 60358
rect 19220 59322 19276 59324
rect 19300 59322 19356 59324
rect 19380 59322 19436 59324
rect 19460 59322 19516 59324
rect 19220 59270 19246 59322
rect 19246 59270 19276 59322
rect 19300 59270 19310 59322
rect 19310 59270 19356 59322
rect 19380 59270 19426 59322
rect 19426 59270 19436 59322
rect 19460 59270 19490 59322
rect 19490 59270 19516 59322
rect 19220 59268 19276 59270
rect 19300 59268 19356 59270
rect 19380 59268 19436 59270
rect 19460 59268 19516 59270
rect 19220 58234 19276 58236
rect 19300 58234 19356 58236
rect 19380 58234 19436 58236
rect 19460 58234 19516 58236
rect 19220 58182 19246 58234
rect 19246 58182 19276 58234
rect 19300 58182 19310 58234
rect 19310 58182 19356 58234
rect 19380 58182 19426 58234
rect 19426 58182 19436 58234
rect 19460 58182 19490 58234
rect 19490 58182 19516 58234
rect 19220 58180 19276 58182
rect 19300 58180 19356 58182
rect 19380 58180 19436 58182
rect 19460 58180 19516 58182
rect 19220 57146 19276 57148
rect 19300 57146 19356 57148
rect 19380 57146 19436 57148
rect 19460 57146 19516 57148
rect 19220 57094 19246 57146
rect 19246 57094 19276 57146
rect 19300 57094 19310 57146
rect 19310 57094 19356 57146
rect 19380 57094 19426 57146
rect 19426 57094 19436 57146
rect 19460 57094 19490 57146
rect 19490 57094 19516 57146
rect 19220 57092 19276 57094
rect 19300 57092 19356 57094
rect 19380 57092 19436 57094
rect 19460 57092 19516 57094
rect 19220 56058 19276 56060
rect 19300 56058 19356 56060
rect 19380 56058 19436 56060
rect 19460 56058 19516 56060
rect 19220 56006 19246 56058
rect 19246 56006 19276 56058
rect 19300 56006 19310 56058
rect 19310 56006 19356 56058
rect 19380 56006 19426 56058
rect 19426 56006 19436 56058
rect 19460 56006 19490 56058
rect 19490 56006 19516 56058
rect 19220 56004 19276 56006
rect 19300 56004 19356 56006
rect 19380 56004 19436 56006
rect 19460 56004 19516 56006
rect 19220 54970 19276 54972
rect 19300 54970 19356 54972
rect 19380 54970 19436 54972
rect 19460 54970 19516 54972
rect 19220 54918 19246 54970
rect 19246 54918 19276 54970
rect 19300 54918 19310 54970
rect 19310 54918 19356 54970
rect 19380 54918 19426 54970
rect 19426 54918 19436 54970
rect 19460 54918 19490 54970
rect 19490 54918 19516 54970
rect 19220 54916 19276 54918
rect 19300 54916 19356 54918
rect 19380 54916 19436 54918
rect 19460 54916 19516 54918
rect 19220 53882 19276 53884
rect 19300 53882 19356 53884
rect 19380 53882 19436 53884
rect 19460 53882 19516 53884
rect 19220 53830 19246 53882
rect 19246 53830 19276 53882
rect 19300 53830 19310 53882
rect 19310 53830 19356 53882
rect 19380 53830 19426 53882
rect 19426 53830 19436 53882
rect 19460 53830 19490 53882
rect 19490 53830 19516 53882
rect 19220 53828 19276 53830
rect 19300 53828 19356 53830
rect 19380 53828 19436 53830
rect 19460 53828 19516 53830
rect 24220 62042 24276 62044
rect 24300 62042 24356 62044
rect 24380 62042 24436 62044
rect 24460 62042 24516 62044
rect 24220 61990 24246 62042
rect 24246 61990 24276 62042
rect 24300 61990 24310 62042
rect 24310 61990 24356 62042
rect 24380 61990 24426 62042
rect 24426 61990 24436 62042
rect 24460 61990 24490 62042
rect 24490 61990 24516 62042
rect 24220 61988 24276 61990
rect 24300 61988 24356 61990
rect 24380 61988 24436 61990
rect 24460 61988 24516 61990
rect 24220 60954 24276 60956
rect 24300 60954 24356 60956
rect 24380 60954 24436 60956
rect 24460 60954 24516 60956
rect 24220 60902 24246 60954
rect 24246 60902 24276 60954
rect 24300 60902 24310 60954
rect 24310 60902 24356 60954
rect 24380 60902 24426 60954
rect 24426 60902 24436 60954
rect 24460 60902 24490 60954
rect 24490 60902 24516 60954
rect 24220 60900 24276 60902
rect 24300 60900 24356 60902
rect 24380 60900 24436 60902
rect 24460 60900 24516 60902
rect 24220 59866 24276 59868
rect 24300 59866 24356 59868
rect 24380 59866 24436 59868
rect 24460 59866 24516 59868
rect 24220 59814 24246 59866
rect 24246 59814 24276 59866
rect 24300 59814 24310 59866
rect 24310 59814 24356 59866
rect 24380 59814 24426 59866
rect 24426 59814 24436 59866
rect 24460 59814 24490 59866
rect 24490 59814 24516 59866
rect 24220 59812 24276 59814
rect 24300 59812 24356 59814
rect 24380 59812 24436 59814
rect 24460 59812 24516 59814
rect 24220 58778 24276 58780
rect 24300 58778 24356 58780
rect 24380 58778 24436 58780
rect 24460 58778 24516 58780
rect 24220 58726 24246 58778
rect 24246 58726 24276 58778
rect 24300 58726 24310 58778
rect 24310 58726 24356 58778
rect 24380 58726 24426 58778
rect 24426 58726 24436 58778
rect 24460 58726 24490 58778
rect 24490 58726 24516 58778
rect 24220 58724 24276 58726
rect 24300 58724 24356 58726
rect 24380 58724 24436 58726
rect 24460 58724 24516 58726
rect 24220 57690 24276 57692
rect 24300 57690 24356 57692
rect 24380 57690 24436 57692
rect 24460 57690 24516 57692
rect 24220 57638 24246 57690
rect 24246 57638 24276 57690
rect 24300 57638 24310 57690
rect 24310 57638 24356 57690
rect 24380 57638 24426 57690
rect 24426 57638 24436 57690
rect 24460 57638 24490 57690
rect 24490 57638 24516 57690
rect 24220 57636 24276 57638
rect 24300 57636 24356 57638
rect 24380 57636 24436 57638
rect 24460 57636 24516 57638
rect 24220 56602 24276 56604
rect 24300 56602 24356 56604
rect 24380 56602 24436 56604
rect 24460 56602 24516 56604
rect 24220 56550 24246 56602
rect 24246 56550 24276 56602
rect 24300 56550 24310 56602
rect 24310 56550 24356 56602
rect 24380 56550 24426 56602
rect 24426 56550 24436 56602
rect 24460 56550 24490 56602
rect 24490 56550 24516 56602
rect 24220 56548 24276 56550
rect 24300 56548 24356 56550
rect 24380 56548 24436 56550
rect 24460 56548 24516 56550
rect 24220 55514 24276 55516
rect 24300 55514 24356 55516
rect 24380 55514 24436 55516
rect 24460 55514 24516 55516
rect 24220 55462 24246 55514
rect 24246 55462 24276 55514
rect 24300 55462 24310 55514
rect 24310 55462 24356 55514
rect 24380 55462 24426 55514
rect 24426 55462 24436 55514
rect 24460 55462 24490 55514
rect 24490 55462 24516 55514
rect 24220 55460 24276 55462
rect 24300 55460 24356 55462
rect 24380 55460 24436 55462
rect 24460 55460 24516 55462
rect 24220 54426 24276 54428
rect 24300 54426 24356 54428
rect 24380 54426 24436 54428
rect 24460 54426 24516 54428
rect 24220 54374 24246 54426
rect 24246 54374 24276 54426
rect 24300 54374 24310 54426
rect 24310 54374 24356 54426
rect 24380 54374 24426 54426
rect 24426 54374 24436 54426
rect 24460 54374 24490 54426
rect 24490 54374 24516 54426
rect 24220 54372 24276 54374
rect 24300 54372 24356 54374
rect 24380 54372 24436 54374
rect 24460 54372 24516 54374
rect 19220 52794 19276 52796
rect 19300 52794 19356 52796
rect 19380 52794 19436 52796
rect 19460 52794 19516 52796
rect 19220 52742 19246 52794
rect 19246 52742 19276 52794
rect 19300 52742 19310 52794
rect 19310 52742 19356 52794
rect 19380 52742 19426 52794
rect 19426 52742 19436 52794
rect 19460 52742 19490 52794
rect 19490 52742 19516 52794
rect 19220 52740 19276 52742
rect 19300 52740 19356 52742
rect 19380 52740 19436 52742
rect 19460 52740 19516 52742
rect 24220 53338 24276 53340
rect 24300 53338 24356 53340
rect 24380 53338 24436 53340
rect 24460 53338 24516 53340
rect 24220 53286 24246 53338
rect 24246 53286 24276 53338
rect 24300 53286 24310 53338
rect 24310 53286 24356 53338
rect 24380 53286 24426 53338
rect 24426 53286 24436 53338
rect 24460 53286 24490 53338
rect 24490 53286 24516 53338
rect 24220 53284 24276 53286
rect 24300 53284 24356 53286
rect 24380 53284 24436 53286
rect 24460 53284 24516 53286
rect 19220 51706 19276 51708
rect 19300 51706 19356 51708
rect 19380 51706 19436 51708
rect 19460 51706 19516 51708
rect 19220 51654 19246 51706
rect 19246 51654 19276 51706
rect 19300 51654 19310 51706
rect 19310 51654 19356 51706
rect 19380 51654 19426 51706
rect 19426 51654 19436 51706
rect 19460 51654 19490 51706
rect 19490 51654 19516 51706
rect 19220 51652 19276 51654
rect 19300 51652 19356 51654
rect 19380 51652 19436 51654
rect 19460 51652 19516 51654
rect 19220 50618 19276 50620
rect 19300 50618 19356 50620
rect 19380 50618 19436 50620
rect 19460 50618 19516 50620
rect 19220 50566 19246 50618
rect 19246 50566 19276 50618
rect 19300 50566 19310 50618
rect 19310 50566 19356 50618
rect 19380 50566 19426 50618
rect 19426 50566 19436 50618
rect 19460 50566 19490 50618
rect 19490 50566 19516 50618
rect 19220 50564 19276 50566
rect 19300 50564 19356 50566
rect 19380 50564 19436 50566
rect 19460 50564 19516 50566
rect 19220 49530 19276 49532
rect 19300 49530 19356 49532
rect 19380 49530 19436 49532
rect 19460 49530 19516 49532
rect 19220 49478 19246 49530
rect 19246 49478 19276 49530
rect 19300 49478 19310 49530
rect 19310 49478 19356 49530
rect 19380 49478 19426 49530
rect 19426 49478 19436 49530
rect 19460 49478 19490 49530
rect 19490 49478 19516 49530
rect 19220 49476 19276 49478
rect 19300 49476 19356 49478
rect 19380 49476 19436 49478
rect 19460 49476 19516 49478
rect 19220 48442 19276 48444
rect 19300 48442 19356 48444
rect 19380 48442 19436 48444
rect 19460 48442 19516 48444
rect 19220 48390 19246 48442
rect 19246 48390 19276 48442
rect 19300 48390 19310 48442
rect 19310 48390 19356 48442
rect 19380 48390 19426 48442
rect 19426 48390 19436 48442
rect 19460 48390 19490 48442
rect 19490 48390 19516 48442
rect 19220 48388 19276 48390
rect 19300 48388 19356 48390
rect 19380 48388 19436 48390
rect 19460 48388 19516 48390
rect 19220 47354 19276 47356
rect 19300 47354 19356 47356
rect 19380 47354 19436 47356
rect 19460 47354 19516 47356
rect 19220 47302 19246 47354
rect 19246 47302 19276 47354
rect 19300 47302 19310 47354
rect 19310 47302 19356 47354
rect 19380 47302 19426 47354
rect 19426 47302 19436 47354
rect 19460 47302 19490 47354
rect 19490 47302 19516 47354
rect 19220 47300 19276 47302
rect 19300 47300 19356 47302
rect 19380 47300 19436 47302
rect 19460 47300 19516 47302
rect 19220 46266 19276 46268
rect 19300 46266 19356 46268
rect 19380 46266 19436 46268
rect 19460 46266 19516 46268
rect 19220 46214 19246 46266
rect 19246 46214 19276 46266
rect 19300 46214 19310 46266
rect 19310 46214 19356 46266
rect 19380 46214 19426 46266
rect 19426 46214 19436 46266
rect 19460 46214 19490 46266
rect 19490 46214 19516 46266
rect 19220 46212 19276 46214
rect 19300 46212 19356 46214
rect 19380 46212 19436 46214
rect 19460 46212 19516 46214
rect 19220 45178 19276 45180
rect 19300 45178 19356 45180
rect 19380 45178 19436 45180
rect 19460 45178 19516 45180
rect 19220 45126 19246 45178
rect 19246 45126 19276 45178
rect 19300 45126 19310 45178
rect 19310 45126 19356 45178
rect 19380 45126 19426 45178
rect 19426 45126 19436 45178
rect 19460 45126 19490 45178
rect 19490 45126 19516 45178
rect 19220 45124 19276 45126
rect 19300 45124 19356 45126
rect 19380 45124 19436 45126
rect 19460 45124 19516 45126
rect 19220 44090 19276 44092
rect 19300 44090 19356 44092
rect 19380 44090 19436 44092
rect 19460 44090 19516 44092
rect 19220 44038 19246 44090
rect 19246 44038 19276 44090
rect 19300 44038 19310 44090
rect 19310 44038 19356 44090
rect 19380 44038 19426 44090
rect 19426 44038 19436 44090
rect 19460 44038 19490 44090
rect 19490 44038 19516 44090
rect 19220 44036 19276 44038
rect 19300 44036 19356 44038
rect 19380 44036 19436 44038
rect 19460 44036 19516 44038
rect 19220 43002 19276 43004
rect 19300 43002 19356 43004
rect 19380 43002 19436 43004
rect 19460 43002 19516 43004
rect 19220 42950 19246 43002
rect 19246 42950 19276 43002
rect 19300 42950 19310 43002
rect 19310 42950 19356 43002
rect 19380 42950 19426 43002
rect 19426 42950 19436 43002
rect 19460 42950 19490 43002
rect 19490 42950 19516 43002
rect 19220 42948 19276 42950
rect 19300 42948 19356 42950
rect 19380 42948 19436 42950
rect 19460 42948 19516 42950
rect 19220 41914 19276 41916
rect 19300 41914 19356 41916
rect 19380 41914 19436 41916
rect 19460 41914 19516 41916
rect 19220 41862 19246 41914
rect 19246 41862 19276 41914
rect 19300 41862 19310 41914
rect 19310 41862 19356 41914
rect 19380 41862 19426 41914
rect 19426 41862 19436 41914
rect 19460 41862 19490 41914
rect 19490 41862 19516 41914
rect 19220 41860 19276 41862
rect 19300 41860 19356 41862
rect 19380 41860 19436 41862
rect 19460 41860 19516 41862
rect 19220 40826 19276 40828
rect 19300 40826 19356 40828
rect 19380 40826 19436 40828
rect 19460 40826 19516 40828
rect 19220 40774 19246 40826
rect 19246 40774 19276 40826
rect 19300 40774 19310 40826
rect 19310 40774 19356 40826
rect 19380 40774 19426 40826
rect 19426 40774 19436 40826
rect 19460 40774 19490 40826
rect 19490 40774 19516 40826
rect 19220 40772 19276 40774
rect 19300 40772 19356 40774
rect 19380 40772 19436 40774
rect 19460 40772 19516 40774
rect 19220 39738 19276 39740
rect 19300 39738 19356 39740
rect 19380 39738 19436 39740
rect 19460 39738 19516 39740
rect 19220 39686 19246 39738
rect 19246 39686 19276 39738
rect 19300 39686 19310 39738
rect 19310 39686 19356 39738
rect 19380 39686 19426 39738
rect 19426 39686 19436 39738
rect 19460 39686 19490 39738
rect 19490 39686 19516 39738
rect 19220 39684 19276 39686
rect 19300 39684 19356 39686
rect 19380 39684 19436 39686
rect 19460 39684 19516 39686
rect 19220 38650 19276 38652
rect 19300 38650 19356 38652
rect 19380 38650 19436 38652
rect 19460 38650 19516 38652
rect 19220 38598 19246 38650
rect 19246 38598 19276 38650
rect 19300 38598 19310 38650
rect 19310 38598 19356 38650
rect 19380 38598 19426 38650
rect 19426 38598 19436 38650
rect 19460 38598 19490 38650
rect 19490 38598 19516 38650
rect 19220 38596 19276 38598
rect 19300 38596 19356 38598
rect 19380 38596 19436 38598
rect 19460 38596 19516 38598
rect 19220 37562 19276 37564
rect 19300 37562 19356 37564
rect 19380 37562 19436 37564
rect 19460 37562 19516 37564
rect 19220 37510 19246 37562
rect 19246 37510 19276 37562
rect 19300 37510 19310 37562
rect 19310 37510 19356 37562
rect 19380 37510 19426 37562
rect 19426 37510 19436 37562
rect 19460 37510 19490 37562
rect 19490 37510 19516 37562
rect 19220 37508 19276 37510
rect 19300 37508 19356 37510
rect 19380 37508 19436 37510
rect 19460 37508 19516 37510
rect 19220 36474 19276 36476
rect 19300 36474 19356 36476
rect 19380 36474 19436 36476
rect 19460 36474 19516 36476
rect 19220 36422 19246 36474
rect 19246 36422 19276 36474
rect 19300 36422 19310 36474
rect 19310 36422 19356 36474
rect 19380 36422 19426 36474
rect 19426 36422 19436 36474
rect 19460 36422 19490 36474
rect 19490 36422 19516 36474
rect 19220 36420 19276 36422
rect 19300 36420 19356 36422
rect 19380 36420 19436 36422
rect 19460 36420 19516 36422
rect 19220 35386 19276 35388
rect 19300 35386 19356 35388
rect 19380 35386 19436 35388
rect 19460 35386 19516 35388
rect 19220 35334 19246 35386
rect 19246 35334 19276 35386
rect 19300 35334 19310 35386
rect 19310 35334 19356 35386
rect 19380 35334 19426 35386
rect 19426 35334 19436 35386
rect 19460 35334 19490 35386
rect 19490 35334 19516 35386
rect 19220 35332 19276 35334
rect 19300 35332 19356 35334
rect 19380 35332 19436 35334
rect 19460 35332 19516 35334
rect 19220 34298 19276 34300
rect 19300 34298 19356 34300
rect 19380 34298 19436 34300
rect 19460 34298 19516 34300
rect 19220 34246 19246 34298
rect 19246 34246 19276 34298
rect 19300 34246 19310 34298
rect 19310 34246 19356 34298
rect 19380 34246 19426 34298
rect 19426 34246 19436 34298
rect 19460 34246 19490 34298
rect 19490 34246 19516 34298
rect 19220 34244 19276 34246
rect 19300 34244 19356 34246
rect 19380 34244 19436 34246
rect 19460 34244 19516 34246
rect 19220 33210 19276 33212
rect 19300 33210 19356 33212
rect 19380 33210 19436 33212
rect 19460 33210 19516 33212
rect 19220 33158 19246 33210
rect 19246 33158 19276 33210
rect 19300 33158 19310 33210
rect 19310 33158 19356 33210
rect 19380 33158 19426 33210
rect 19426 33158 19436 33210
rect 19460 33158 19490 33210
rect 19490 33158 19516 33210
rect 19220 33156 19276 33158
rect 19300 33156 19356 33158
rect 19380 33156 19436 33158
rect 19460 33156 19516 33158
rect 19220 32122 19276 32124
rect 19300 32122 19356 32124
rect 19380 32122 19436 32124
rect 19460 32122 19516 32124
rect 19220 32070 19246 32122
rect 19246 32070 19276 32122
rect 19300 32070 19310 32122
rect 19310 32070 19356 32122
rect 19380 32070 19426 32122
rect 19426 32070 19436 32122
rect 19460 32070 19490 32122
rect 19490 32070 19516 32122
rect 19220 32068 19276 32070
rect 19300 32068 19356 32070
rect 19380 32068 19436 32070
rect 19460 32068 19516 32070
rect 19220 31034 19276 31036
rect 19300 31034 19356 31036
rect 19380 31034 19436 31036
rect 19460 31034 19516 31036
rect 19220 30982 19246 31034
rect 19246 30982 19276 31034
rect 19300 30982 19310 31034
rect 19310 30982 19356 31034
rect 19380 30982 19426 31034
rect 19426 30982 19436 31034
rect 19460 30982 19490 31034
rect 19490 30982 19516 31034
rect 19220 30980 19276 30982
rect 19300 30980 19356 30982
rect 19380 30980 19436 30982
rect 19460 30980 19516 30982
rect 19220 29946 19276 29948
rect 19300 29946 19356 29948
rect 19380 29946 19436 29948
rect 19460 29946 19516 29948
rect 19220 29894 19246 29946
rect 19246 29894 19276 29946
rect 19300 29894 19310 29946
rect 19310 29894 19356 29946
rect 19380 29894 19426 29946
rect 19426 29894 19436 29946
rect 19460 29894 19490 29946
rect 19490 29894 19516 29946
rect 19220 29892 19276 29894
rect 19300 29892 19356 29894
rect 19380 29892 19436 29894
rect 19460 29892 19516 29894
rect 19220 28858 19276 28860
rect 19300 28858 19356 28860
rect 19380 28858 19436 28860
rect 19460 28858 19516 28860
rect 19220 28806 19246 28858
rect 19246 28806 19276 28858
rect 19300 28806 19310 28858
rect 19310 28806 19356 28858
rect 19380 28806 19426 28858
rect 19426 28806 19436 28858
rect 19460 28806 19490 28858
rect 19490 28806 19516 28858
rect 19220 28804 19276 28806
rect 19300 28804 19356 28806
rect 19380 28804 19436 28806
rect 19460 28804 19516 28806
rect 19220 27770 19276 27772
rect 19300 27770 19356 27772
rect 19380 27770 19436 27772
rect 19460 27770 19516 27772
rect 19220 27718 19246 27770
rect 19246 27718 19276 27770
rect 19300 27718 19310 27770
rect 19310 27718 19356 27770
rect 19380 27718 19426 27770
rect 19426 27718 19436 27770
rect 19460 27718 19490 27770
rect 19490 27718 19516 27770
rect 19220 27716 19276 27718
rect 19300 27716 19356 27718
rect 19380 27716 19436 27718
rect 19460 27716 19516 27718
rect 17498 12280 17554 12336
rect 17498 8744 17554 8800
rect 17498 3440 17554 3496
rect 19220 26682 19276 26684
rect 19300 26682 19356 26684
rect 19380 26682 19436 26684
rect 19460 26682 19516 26684
rect 19220 26630 19246 26682
rect 19246 26630 19276 26682
rect 19300 26630 19310 26682
rect 19310 26630 19356 26682
rect 19380 26630 19426 26682
rect 19426 26630 19436 26682
rect 19460 26630 19490 26682
rect 19490 26630 19516 26682
rect 19220 26628 19276 26630
rect 19300 26628 19356 26630
rect 19380 26628 19436 26630
rect 19460 26628 19516 26630
rect 19220 25594 19276 25596
rect 19300 25594 19356 25596
rect 19380 25594 19436 25596
rect 19460 25594 19516 25596
rect 19220 25542 19246 25594
rect 19246 25542 19276 25594
rect 19300 25542 19310 25594
rect 19310 25542 19356 25594
rect 19380 25542 19426 25594
rect 19426 25542 19436 25594
rect 19460 25542 19490 25594
rect 19490 25542 19516 25594
rect 19220 25540 19276 25542
rect 19300 25540 19356 25542
rect 19380 25540 19436 25542
rect 19460 25540 19516 25542
rect 19220 24506 19276 24508
rect 19300 24506 19356 24508
rect 19380 24506 19436 24508
rect 19460 24506 19516 24508
rect 19220 24454 19246 24506
rect 19246 24454 19276 24506
rect 19300 24454 19310 24506
rect 19310 24454 19356 24506
rect 19380 24454 19426 24506
rect 19426 24454 19436 24506
rect 19460 24454 19490 24506
rect 19490 24454 19516 24506
rect 19220 24452 19276 24454
rect 19300 24452 19356 24454
rect 19380 24452 19436 24454
rect 19460 24452 19516 24454
rect 24220 52250 24276 52252
rect 24300 52250 24356 52252
rect 24380 52250 24436 52252
rect 24460 52250 24516 52252
rect 24220 52198 24246 52250
rect 24246 52198 24276 52250
rect 24300 52198 24310 52250
rect 24310 52198 24356 52250
rect 24380 52198 24426 52250
rect 24426 52198 24436 52250
rect 24460 52198 24490 52250
rect 24490 52198 24516 52250
rect 24220 52196 24276 52198
rect 24300 52196 24356 52198
rect 24380 52196 24436 52198
rect 24460 52196 24516 52198
rect 24220 51162 24276 51164
rect 24300 51162 24356 51164
rect 24380 51162 24436 51164
rect 24460 51162 24516 51164
rect 24220 51110 24246 51162
rect 24246 51110 24276 51162
rect 24300 51110 24310 51162
rect 24310 51110 24356 51162
rect 24380 51110 24426 51162
rect 24426 51110 24436 51162
rect 24460 51110 24490 51162
rect 24490 51110 24516 51162
rect 24220 51108 24276 51110
rect 24300 51108 24356 51110
rect 24380 51108 24436 51110
rect 24460 51108 24516 51110
rect 24220 50074 24276 50076
rect 24300 50074 24356 50076
rect 24380 50074 24436 50076
rect 24460 50074 24516 50076
rect 24220 50022 24246 50074
rect 24246 50022 24276 50074
rect 24300 50022 24310 50074
rect 24310 50022 24356 50074
rect 24380 50022 24426 50074
rect 24426 50022 24436 50074
rect 24460 50022 24490 50074
rect 24490 50022 24516 50074
rect 24220 50020 24276 50022
rect 24300 50020 24356 50022
rect 24380 50020 24436 50022
rect 24460 50020 24516 50022
rect 24220 48986 24276 48988
rect 24300 48986 24356 48988
rect 24380 48986 24436 48988
rect 24460 48986 24516 48988
rect 24220 48934 24246 48986
rect 24246 48934 24276 48986
rect 24300 48934 24310 48986
rect 24310 48934 24356 48986
rect 24380 48934 24426 48986
rect 24426 48934 24436 48986
rect 24460 48934 24490 48986
rect 24490 48934 24516 48986
rect 24220 48932 24276 48934
rect 24300 48932 24356 48934
rect 24380 48932 24436 48934
rect 24460 48932 24516 48934
rect 24220 47898 24276 47900
rect 24300 47898 24356 47900
rect 24380 47898 24436 47900
rect 24460 47898 24516 47900
rect 24220 47846 24246 47898
rect 24246 47846 24276 47898
rect 24300 47846 24310 47898
rect 24310 47846 24356 47898
rect 24380 47846 24426 47898
rect 24426 47846 24436 47898
rect 24460 47846 24490 47898
rect 24490 47846 24516 47898
rect 24220 47844 24276 47846
rect 24300 47844 24356 47846
rect 24380 47844 24436 47846
rect 24460 47844 24516 47846
rect 24220 46810 24276 46812
rect 24300 46810 24356 46812
rect 24380 46810 24436 46812
rect 24460 46810 24516 46812
rect 24220 46758 24246 46810
rect 24246 46758 24276 46810
rect 24300 46758 24310 46810
rect 24310 46758 24356 46810
rect 24380 46758 24426 46810
rect 24426 46758 24436 46810
rect 24460 46758 24490 46810
rect 24490 46758 24516 46810
rect 24220 46756 24276 46758
rect 24300 46756 24356 46758
rect 24380 46756 24436 46758
rect 24460 46756 24516 46758
rect 24220 45722 24276 45724
rect 24300 45722 24356 45724
rect 24380 45722 24436 45724
rect 24460 45722 24516 45724
rect 24220 45670 24246 45722
rect 24246 45670 24276 45722
rect 24300 45670 24310 45722
rect 24310 45670 24356 45722
rect 24380 45670 24426 45722
rect 24426 45670 24436 45722
rect 24460 45670 24490 45722
rect 24490 45670 24516 45722
rect 24220 45668 24276 45670
rect 24300 45668 24356 45670
rect 24380 45668 24436 45670
rect 24460 45668 24516 45670
rect 24220 44634 24276 44636
rect 24300 44634 24356 44636
rect 24380 44634 24436 44636
rect 24460 44634 24516 44636
rect 24220 44582 24246 44634
rect 24246 44582 24276 44634
rect 24300 44582 24310 44634
rect 24310 44582 24356 44634
rect 24380 44582 24426 44634
rect 24426 44582 24436 44634
rect 24460 44582 24490 44634
rect 24490 44582 24516 44634
rect 24220 44580 24276 44582
rect 24300 44580 24356 44582
rect 24380 44580 24436 44582
rect 24460 44580 24516 44582
rect 24220 43546 24276 43548
rect 24300 43546 24356 43548
rect 24380 43546 24436 43548
rect 24460 43546 24516 43548
rect 24220 43494 24246 43546
rect 24246 43494 24276 43546
rect 24300 43494 24310 43546
rect 24310 43494 24356 43546
rect 24380 43494 24426 43546
rect 24426 43494 24436 43546
rect 24460 43494 24490 43546
rect 24490 43494 24516 43546
rect 24220 43492 24276 43494
rect 24300 43492 24356 43494
rect 24380 43492 24436 43494
rect 24460 43492 24516 43494
rect 24220 42458 24276 42460
rect 24300 42458 24356 42460
rect 24380 42458 24436 42460
rect 24460 42458 24516 42460
rect 24220 42406 24246 42458
rect 24246 42406 24276 42458
rect 24300 42406 24310 42458
rect 24310 42406 24356 42458
rect 24380 42406 24426 42458
rect 24426 42406 24436 42458
rect 24460 42406 24490 42458
rect 24490 42406 24516 42458
rect 24220 42404 24276 42406
rect 24300 42404 24356 42406
rect 24380 42404 24436 42406
rect 24460 42404 24516 42406
rect 24220 41370 24276 41372
rect 24300 41370 24356 41372
rect 24380 41370 24436 41372
rect 24460 41370 24516 41372
rect 24220 41318 24246 41370
rect 24246 41318 24276 41370
rect 24300 41318 24310 41370
rect 24310 41318 24356 41370
rect 24380 41318 24426 41370
rect 24426 41318 24436 41370
rect 24460 41318 24490 41370
rect 24490 41318 24516 41370
rect 24220 41316 24276 41318
rect 24300 41316 24356 41318
rect 24380 41316 24436 41318
rect 24460 41316 24516 41318
rect 19220 23418 19276 23420
rect 19300 23418 19356 23420
rect 19380 23418 19436 23420
rect 19460 23418 19516 23420
rect 19220 23366 19246 23418
rect 19246 23366 19276 23418
rect 19300 23366 19310 23418
rect 19310 23366 19356 23418
rect 19380 23366 19426 23418
rect 19426 23366 19436 23418
rect 19460 23366 19490 23418
rect 19490 23366 19516 23418
rect 19220 23364 19276 23366
rect 19300 23364 19356 23366
rect 19380 23364 19436 23366
rect 19460 23364 19516 23366
rect 19220 22330 19276 22332
rect 19300 22330 19356 22332
rect 19380 22330 19436 22332
rect 19460 22330 19516 22332
rect 19220 22278 19246 22330
rect 19246 22278 19276 22330
rect 19300 22278 19310 22330
rect 19310 22278 19356 22330
rect 19380 22278 19426 22330
rect 19426 22278 19436 22330
rect 19460 22278 19490 22330
rect 19490 22278 19516 22330
rect 19220 22276 19276 22278
rect 19300 22276 19356 22278
rect 19380 22276 19436 22278
rect 19460 22276 19516 22278
rect 18326 11192 18382 11248
rect 18234 10804 18290 10840
rect 18234 10784 18236 10804
rect 18236 10784 18288 10804
rect 18288 10784 18290 10804
rect 18326 2760 18382 2816
rect 18326 2624 18382 2680
rect 19220 21242 19276 21244
rect 19300 21242 19356 21244
rect 19380 21242 19436 21244
rect 19460 21242 19516 21244
rect 19220 21190 19246 21242
rect 19246 21190 19276 21242
rect 19300 21190 19310 21242
rect 19310 21190 19356 21242
rect 19380 21190 19426 21242
rect 19426 21190 19436 21242
rect 19460 21190 19490 21242
rect 19490 21190 19516 21242
rect 19220 21188 19276 21190
rect 19300 21188 19356 21190
rect 19380 21188 19436 21190
rect 19460 21188 19516 21190
rect 19220 20154 19276 20156
rect 19300 20154 19356 20156
rect 19380 20154 19436 20156
rect 19460 20154 19516 20156
rect 19220 20102 19246 20154
rect 19246 20102 19276 20154
rect 19300 20102 19310 20154
rect 19310 20102 19356 20154
rect 19380 20102 19426 20154
rect 19426 20102 19436 20154
rect 19460 20102 19490 20154
rect 19490 20102 19516 20154
rect 19220 20100 19276 20102
rect 19300 20100 19356 20102
rect 19380 20100 19436 20102
rect 19460 20100 19516 20102
rect 24220 40282 24276 40284
rect 24300 40282 24356 40284
rect 24380 40282 24436 40284
rect 24460 40282 24516 40284
rect 24220 40230 24246 40282
rect 24246 40230 24276 40282
rect 24300 40230 24310 40282
rect 24310 40230 24356 40282
rect 24380 40230 24426 40282
rect 24426 40230 24436 40282
rect 24460 40230 24490 40282
rect 24490 40230 24516 40282
rect 24220 40228 24276 40230
rect 24300 40228 24356 40230
rect 24380 40228 24436 40230
rect 24460 40228 24516 40230
rect 24220 39194 24276 39196
rect 24300 39194 24356 39196
rect 24380 39194 24436 39196
rect 24460 39194 24516 39196
rect 24220 39142 24246 39194
rect 24246 39142 24276 39194
rect 24300 39142 24310 39194
rect 24310 39142 24356 39194
rect 24380 39142 24426 39194
rect 24426 39142 24436 39194
rect 24460 39142 24490 39194
rect 24490 39142 24516 39194
rect 24220 39140 24276 39142
rect 24300 39140 24356 39142
rect 24380 39140 24436 39142
rect 24460 39140 24516 39142
rect 24220 38106 24276 38108
rect 24300 38106 24356 38108
rect 24380 38106 24436 38108
rect 24460 38106 24516 38108
rect 24220 38054 24246 38106
rect 24246 38054 24276 38106
rect 24300 38054 24310 38106
rect 24310 38054 24356 38106
rect 24380 38054 24426 38106
rect 24426 38054 24436 38106
rect 24460 38054 24490 38106
rect 24490 38054 24516 38106
rect 24220 38052 24276 38054
rect 24300 38052 24356 38054
rect 24380 38052 24436 38054
rect 24460 38052 24516 38054
rect 24220 37018 24276 37020
rect 24300 37018 24356 37020
rect 24380 37018 24436 37020
rect 24460 37018 24516 37020
rect 24220 36966 24246 37018
rect 24246 36966 24276 37018
rect 24300 36966 24310 37018
rect 24310 36966 24356 37018
rect 24380 36966 24426 37018
rect 24426 36966 24436 37018
rect 24460 36966 24490 37018
rect 24490 36966 24516 37018
rect 24220 36964 24276 36966
rect 24300 36964 24356 36966
rect 24380 36964 24436 36966
rect 24460 36964 24516 36966
rect 24220 35930 24276 35932
rect 24300 35930 24356 35932
rect 24380 35930 24436 35932
rect 24460 35930 24516 35932
rect 24220 35878 24246 35930
rect 24246 35878 24276 35930
rect 24300 35878 24310 35930
rect 24310 35878 24356 35930
rect 24380 35878 24426 35930
rect 24426 35878 24436 35930
rect 24460 35878 24490 35930
rect 24490 35878 24516 35930
rect 24220 35876 24276 35878
rect 24300 35876 24356 35878
rect 24380 35876 24436 35878
rect 24460 35876 24516 35878
rect 24220 34842 24276 34844
rect 24300 34842 24356 34844
rect 24380 34842 24436 34844
rect 24460 34842 24516 34844
rect 24220 34790 24246 34842
rect 24246 34790 24276 34842
rect 24300 34790 24310 34842
rect 24310 34790 24356 34842
rect 24380 34790 24426 34842
rect 24426 34790 24436 34842
rect 24460 34790 24490 34842
rect 24490 34790 24516 34842
rect 24220 34788 24276 34790
rect 24300 34788 24356 34790
rect 24380 34788 24436 34790
rect 24460 34788 24516 34790
rect 24220 33754 24276 33756
rect 24300 33754 24356 33756
rect 24380 33754 24436 33756
rect 24460 33754 24516 33756
rect 24220 33702 24246 33754
rect 24246 33702 24276 33754
rect 24300 33702 24310 33754
rect 24310 33702 24356 33754
rect 24380 33702 24426 33754
rect 24426 33702 24436 33754
rect 24460 33702 24490 33754
rect 24490 33702 24516 33754
rect 24220 33700 24276 33702
rect 24300 33700 24356 33702
rect 24380 33700 24436 33702
rect 24460 33700 24516 33702
rect 24220 32666 24276 32668
rect 24300 32666 24356 32668
rect 24380 32666 24436 32668
rect 24460 32666 24516 32668
rect 24220 32614 24246 32666
rect 24246 32614 24276 32666
rect 24300 32614 24310 32666
rect 24310 32614 24356 32666
rect 24380 32614 24426 32666
rect 24426 32614 24436 32666
rect 24460 32614 24490 32666
rect 24490 32614 24516 32666
rect 24220 32612 24276 32614
rect 24300 32612 24356 32614
rect 24380 32612 24436 32614
rect 24460 32612 24516 32614
rect 24220 31578 24276 31580
rect 24300 31578 24356 31580
rect 24380 31578 24436 31580
rect 24460 31578 24516 31580
rect 24220 31526 24246 31578
rect 24246 31526 24276 31578
rect 24300 31526 24310 31578
rect 24310 31526 24356 31578
rect 24380 31526 24426 31578
rect 24426 31526 24436 31578
rect 24460 31526 24490 31578
rect 24490 31526 24516 31578
rect 24220 31524 24276 31526
rect 24300 31524 24356 31526
rect 24380 31524 24436 31526
rect 24460 31524 24516 31526
rect 24220 30490 24276 30492
rect 24300 30490 24356 30492
rect 24380 30490 24436 30492
rect 24460 30490 24516 30492
rect 24220 30438 24246 30490
rect 24246 30438 24276 30490
rect 24300 30438 24310 30490
rect 24310 30438 24356 30490
rect 24380 30438 24426 30490
rect 24426 30438 24436 30490
rect 24460 30438 24490 30490
rect 24490 30438 24516 30490
rect 24220 30436 24276 30438
rect 24300 30436 24356 30438
rect 24380 30436 24436 30438
rect 24460 30436 24516 30438
rect 24220 29402 24276 29404
rect 24300 29402 24356 29404
rect 24380 29402 24436 29404
rect 24460 29402 24516 29404
rect 24220 29350 24246 29402
rect 24246 29350 24276 29402
rect 24300 29350 24310 29402
rect 24310 29350 24356 29402
rect 24380 29350 24426 29402
rect 24426 29350 24436 29402
rect 24460 29350 24490 29402
rect 24490 29350 24516 29402
rect 24220 29348 24276 29350
rect 24300 29348 24356 29350
rect 24380 29348 24436 29350
rect 24460 29348 24516 29350
rect 24220 28314 24276 28316
rect 24300 28314 24356 28316
rect 24380 28314 24436 28316
rect 24460 28314 24516 28316
rect 24220 28262 24246 28314
rect 24246 28262 24276 28314
rect 24300 28262 24310 28314
rect 24310 28262 24356 28314
rect 24380 28262 24426 28314
rect 24426 28262 24436 28314
rect 24460 28262 24490 28314
rect 24490 28262 24516 28314
rect 24220 28260 24276 28262
rect 24300 28260 24356 28262
rect 24380 28260 24436 28262
rect 24460 28260 24516 28262
rect 24220 27226 24276 27228
rect 24300 27226 24356 27228
rect 24380 27226 24436 27228
rect 24460 27226 24516 27228
rect 24220 27174 24246 27226
rect 24246 27174 24276 27226
rect 24300 27174 24310 27226
rect 24310 27174 24356 27226
rect 24380 27174 24426 27226
rect 24426 27174 24436 27226
rect 24460 27174 24490 27226
rect 24490 27174 24516 27226
rect 24220 27172 24276 27174
rect 24300 27172 24356 27174
rect 24380 27172 24436 27174
rect 24460 27172 24516 27174
rect 24220 26138 24276 26140
rect 24300 26138 24356 26140
rect 24380 26138 24436 26140
rect 24460 26138 24516 26140
rect 24220 26086 24246 26138
rect 24246 26086 24276 26138
rect 24300 26086 24310 26138
rect 24310 26086 24356 26138
rect 24380 26086 24426 26138
rect 24426 26086 24436 26138
rect 24460 26086 24490 26138
rect 24490 26086 24516 26138
rect 24220 26084 24276 26086
rect 24300 26084 24356 26086
rect 24380 26084 24436 26086
rect 24460 26084 24516 26086
rect 24220 25050 24276 25052
rect 24300 25050 24356 25052
rect 24380 25050 24436 25052
rect 24460 25050 24516 25052
rect 24220 24998 24246 25050
rect 24246 24998 24276 25050
rect 24300 24998 24310 25050
rect 24310 24998 24356 25050
rect 24380 24998 24426 25050
rect 24426 24998 24436 25050
rect 24460 24998 24490 25050
rect 24490 24998 24516 25050
rect 24220 24996 24276 24998
rect 24300 24996 24356 24998
rect 24380 24996 24436 24998
rect 24460 24996 24516 24998
rect 24220 23962 24276 23964
rect 24300 23962 24356 23964
rect 24380 23962 24436 23964
rect 24460 23962 24516 23964
rect 24220 23910 24246 23962
rect 24246 23910 24276 23962
rect 24300 23910 24310 23962
rect 24310 23910 24356 23962
rect 24380 23910 24426 23962
rect 24426 23910 24436 23962
rect 24460 23910 24490 23962
rect 24490 23910 24516 23962
rect 24220 23908 24276 23910
rect 24300 23908 24356 23910
rect 24380 23908 24436 23910
rect 24460 23908 24516 23910
rect 24220 22874 24276 22876
rect 24300 22874 24356 22876
rect 24380 22874 24436 22876
rect 24460 22874 24516 22876
rect 24220 22822 24246 22874
rect 24246 22822 24276 22874
rect 24300 22822 24310 22874
rect 24310 22822 24356 22874
rect 24380 22822 24426 22874
rect 24426 22822 24436 22874
rect 24460 22822 24490 22874
rect 24490 22822 24516 22874
rect 24220 22820 24276 22822
rect 24300 22820 24356 22822
rect 24380 22820 24436 22822
rect 24460 22820 24516 22822
rect 22098 17176 22154 17232
rect 24220 21786 24276 21788
rect 24300 21786 24356 21788
rect 24380 21786 24436 21788
rect 24460 21786 24516 21788
rect 24220 21734 24246 21786
rect 24246 21734 24276 21786
rect 24300 21734 24310 21786
rect 24310 21734 24356 21786
rect 24380 21734 24426 21786
rect 24426 21734 24436 21786
rect 24460 21734 24490 21786
rect 24490 21734 24516 21786
rect 24220 21732 24276 21734
rect 24300 21732 24356 21734
rect 24380 21732 24436 21734
rect 24460 21732 24516 21734
rect 29220 66938 29276 66940
rect 29300 66938 29356 66940
rect 29380 66938 29436 66940
rect 29460 66938 29516 66940
rect 29220 66886 29246 66938
rect 29246 66886 29276 66938
rect 29300 66886 29310 66938
rect 29310 66886 29356 66938
rect 29380 66886 29426 66938
rect 29426 66886 29436 66938
rect 29460 66886 29490 66938
rect 29490 66886 29516 66938
rect 29220 66884 29276 66886
rect 29300 66884 29356 66886
rect 29380 66884 29436 66886
rect 29460 66884 29516 66886
rect 29220 65850 29276 65852
rect 29300 65850 29356 65852
rect 29380 65850 29436 65852
rect 29460 65850 29516 65852
rect 29220 65798 29246 65850
rect 29246 65798 29276 65850
rect 29300 65798 29310 65850
rect 29310 65798 29356 65850
rect 29380 65798 29426 65850
rect 29426 65798 29436 65850
rect 29460 65798 29490 65850
rect 29490 65798 29516 65850
rect 29220 65796 29276 65798
rect 29300 65796 29356 65798
rect 29380 65796 29436 65798
rect 29460 65796 29516 65798
rect 29220 64762 29276 64764
rect 29300 64762 29356 64764
rect 29380 64762 29436 64764
rect 29460 64762 29516 64764
rect 29220 64710 29246 64762
rect 29246 64710 29276 64762
rect 29300 64710 29310 64762
rect 29310 64710 29356 64762
rect 29380 64710 29426 64762
rect 29426 64710 29436 64762
rect 29460 64710 29490 64762
rect 29490 64710 29516 64762
rect 29220 64708 29276 64710
rect 29300 64708 29356 64710
rect 29380 64708 29436 64710
rect 29460 64708 29516 64710
rect 29220 63674 29276 63676
rect 29300 63674 29356 63676
rect 29380 63674 29436 63676
rect 29460 63674 29516 63676
rect 29220 63622 29246 63674
rect 29246 63622 29276 63674
rect 29300 63622 29310 63674
rect 29310 63622 29356 63674
rect 29380 63622 29426 63674
rect 29426 63622 29436 63674
rect 29460 63622 29490 63674
rect 29490 63622 29516 63674
rect 29220 63620 29276 63622
rect 29300 63620 29356 63622
rect 29380 63620 29436 63622
rect 29460 63620 29516 63622
rect 29220 62586 29276 62588
rect 29300 62586 29356 62588
rect 29380 62586 29436 62588
rect 29460 62586 29516 62588
rect 29220 62534 29246 62586
rect 29246 62534 29276 62586
rect 29300 62534 29310 62586
rect 29310 62534 29356 62586
rect 29380 62534 29426 62586
rect 29426 62534 29436 62586
rect 29460 62534 29490 62586
rect 29490 62534 29516 62586
rect 29220 62532 29276 62534
rect 29300 62532 29356 62534
rect 29380 62532 29436 62534
rect 29460 62532 29516 62534
rect 29220 61498 29276 61500
rect 29300 61498 29356 61500
rect 29380 61498 29436 61500
rect 29460 61498 29516 61500
rect 29220 61446 29246 61498
rect 29246 61446 29276 61498
rect 29300 61446 29310 61498
rect 29310 61446 29356 61498
rect 29380 61446 29426 61498
rect 29426 61446 29436 61498
rect 29460 61446 29490 61498
rect 29490 61446 29516 61498
rect 29220 61444 29276 61446
rect 29300 61444 29356 61446
rect 29380 61444 29436 61446
rect 29460 61444 29516 61446
rect 29220 60410 29276 60412
rect 29300 60410 29356 60412
rect 29380 60410 29436 60412
rect 29460 60410 29516 60412
rect 29220 60358 29246 60410
rect 29246 60358 29276 60410
rect 29300 60358 29310 60410
rect 29310 60358 29356 60410
rect 29380 60358 29426 60410
rect 29426 60358 29436 60410
rect 29460 60358 29490 60410
rect 29490 60358 29516 60410
rect 29220 60356 29276 60358
rect 29300 60356 29356 60358
rect 29380 60356 29436 60358
rect 29460 60356 29516 60358
rect 29220 59322 29276 59324
rect 29300 59322 29356 59324
rect 29380 59322 29436 59324
rect 29460 59322 29516 59324
rect 29220 59270 29246 59322
rect 29246 59270 29276 59322
rect 29300 59270 29310 59322
rect 29310 59270 29356 59322
rect 29380 59270 29426 59322
rect 29426 59270 29436 59322
rect 29460 59270 29490 59322
rect 29490 59270 29516 59322
rect 29220 59268 29276 59270
rect 29300 59268 29356 59270
rect 29380 59268 29436 59270
rect 29460 59268 29516 59270
rect 24220 20698 24276 20700
rect 24300 20698 24356 20700
rect 24380 20698 24436 20700
rect 24460 20698 24516 20700
rect 24220 20646 24246 20698
rect 24246 20646 24276 20698
rect 24300 20646 24310 20698
rect 24310 20646 24356 20698
rect 24380 20646 24426 20698
rect 24426 20646 24436 20698
rect 24460 20646 24490 20698
rect 24490 20646 24516 20698
rect 24220 20644 24276 20646
rect 24300 20644 24356 20646
rect 24380 20644 24436 20646
rect 24460 20644 24516 20646
rect 24220 19610 24276 19612
rect 24300 19610 24356 19612
rect 24380 19610 24436 19612
rect 24460 19610 24516 19612
rect 24220 19558 24246 19610
rect 24246 19558 24276 19610
rect 24300 19558 24310 19610
rect 24310 19558 24356 19610
rect 24380 19558 24426 19610
rect 24426 19558 24436 19610
rect 24460 19558 24490 19610
rect 24490 19558 24516 19610
rect 24220 19556 24276 19558
rect 24300 19556 24356 19558
rect 24380 19556 24436 19558
rect 24460 19556 24516 19558
rect 29220 58234 29276 58236
rect 29300 58234 29356 58236
rect 29380 58234 29436 58236
rect 29460 58234 29516 58236
rect 29220 58182 29246 58234
rect 29246 58182 29276 58234
rect 29300 58182 29310 58234
rect 29310 58182 29356 58234
rect 29380 58182 29426 58234
rect 29426 58182 29436 58234
rect 29460 58182 29490 58234
rect 29490 58182 29516 58234
rect 29220 58180 29276 58182
rect 29300 58180 29356 58182
rect 29380 58180 29436 58182
rect 29460 58180 29516 58182
rect 29220 57146 29276 57148
rect 29300 57146 29356 57148
rect 29380 57146 29436 57148
rect 29460 57146 29516 57148
rect 29220 57094 29246 57146
rect 29246 57094 29276 57146
rect 29300 57094 29310 57146
rect 29310 57094 29356 57146
rect 29380 57094 29426 57146
rect 29426 57094 29436 57146
rect 29460 57094 29490 57146
rect 29490 57094 29516 57146
rect 29220 57092 29276 57094
rect 29300 57092 29356 57094
rect 29380 57092 29436 57094
rect 29460 57092 29516 57094
rect 29220 56058 29276 56060
rect 29300 56058 29356 56060
rect 29380 56058 29436 56060
rect 29460 56058 29516 56060
rect 29220 56006 29246 56058
rect 29246 56006 29276 56058
rect 29300 56006 29310 56058
rect 29310 56006 29356 56058
rect 29380 56006 29426 56058
rect 29426 56006 29436 56058
rect 29460 56006 29490 56058
rect 29490 56006 29516 56058
rect 29220 56004 29276 56006
rect 29300 56004 29356 56006
rect 29380 56004 29436 56006
rect 29460 56004 29516 56006
rect 29220 54970 29276 54972
rect 29300 54970 29356 54972
rect 29380 54970 29436 54972
rect 29460 54970 29516 54972
rect 29220 54918 29246 54970
rect 29246 54918 29276 54970
rect 29300 54918 29310 54970
rect 29310 54918 29356 54970
rect 29380 54918 29426 54970
rect 29426 54918 29436 54970
rect 29460 54918 29490 54970
rect 29490 54918 29516 54970
rect 29220 54916 29276 54918
rect 29300 54916 29356 54918
rect 29380 54916 29436 54918
rect 29460 54916 29516 54918
rect 29220 53882 29276 53884
rect 29300 53882 29356 53884
rect 29380 53882 29436 53884
rect 29460 53882 29516 53884
rect 29220 53830 29246 53882
rect 29246 53830 29276 53882
rect 29300 53830 29310 53882
rect 29310 53830 29356 53882
rect 29380 53830 29426 53882
rect 29426 53830 29436 53882
rect 29460 53830 29490 53882
rect 29490 53830 29516 53882
rect 29220 53828 29276 53830
rect 29300 53828 29356 53830
rect 29380 53828 29436 53830
rect 29460 53828 29516 53830
rect 29220 52794 29276 52796
rect 29300 52794 29356 52796
rect 29380 52794 29436 52796
rect 29460 52794 29516 52796
rect 29220 52742 29246 52794
rect 29246 52742 29276 52794
rect 29300 52742 29310 52794
rect 29310 52742 29356 52794
rect 29380 52742 29426 52794
rect 29426 52742 29436 52794
rect 29460 52742 29490 52794
rect 29490 52742 29516 52794
rect 29220 52740 29276 52742
rect 29300 52740 29356 52742
rect 29380 52740 29436 52742
rect 29460 52740 29516 52742
rect 29220 51706 29276 51708
rect 29300 51706 29356 51708
rect 29380 51706 29436 51708
rect 29460 51706 29516 51708
rect 29220 51654 29246 51706
rect 29246 51654 29276 51706
rect 29300 51654 29310 51706
rect 29310 51654 29356 51706
rect 29380 51654 29426 51706
rect 29426 51654 29436 51706
rect 29460 51654 29490 51706
rect 29490 51654 29516 51706
rect 29220 51652 29276 51654
rect 29300 51652 29356 51654
rect 29380 51652 29436 51654
rect 29460 51652 29516 51654
rect 29220 50618 29276 50620
rect 29300 50618 29356 50620
rect 29380 50618 29436 50620
rect 29460 50618 29516 50620
rect 29220 50566 29246 50618
rect 29246 50566 29276 50618
rect 29300 50566 29310 50618
rect 29310 50566 29356 50618
rect 29380 50566 29426 50618
rect 29426 50566 29436 50618
rect 29460 50566 29490 50618
rect 29490 50566 29516 50618
rect 29220 50564 29276 50566
rect 29300 50564 29356 50566
rect 29380 50564 29436 50566
rect 29460 50564 29516 50566
rect 29220 49530 29276 49532
rect 29300 49530 29356 49532
rect 29380 49530 29436 49532
rect 29460 49530 29516 49532
rect 29220 49478 29246 49530
rect 29246 49478 29276 49530
rect 29300 49478 29310 49530
rect 29310 49478 29356 49530
rect 29380 49478 29426 49530
rect 29426 49478 29436 49530
rect 29460 49478 29490 49530
rect 29490 49478 29516 49530
rect 29220 49476 29276 49478
rect 29300 49476 29356 49478
rect 29380 49476 29436 49478
rect 29460 49476 29516 49478
rect 29220 48442 29276 48444
rect 29300 48442 29356 48444
rect 29380 48442 29436 48444
rect 29460 48442 29516 48444
rect 29220 48390 29246 48442
rect 29246 48390 29276 48442
rect 29300 48390 29310 48442
rect 29310 48390 29356 48442
rect 29380 48390 29426 48442
rect 29426 48390 29436 48442
rect 29460 48390 29490 48442
rect 29490 48390 29516 48442
rect 29220 48388 29276 48390
rect 29300 48388 29356 48390
rect 29380 48388 29436 48390
rect 29460 48388 29516 48390
rect 29220 47354 29276 47356
rect 29300 47354 29356 47356
rect 29380 47354 29436 47356
rect 29460 47354 29516 47356
rect 29220 47302 29246 47354
rect 29246 47302 29276 47354
rect 29300 47302 29310 47354
rect 29310 47302 29356 47354
rect 29380 47302 29426 47354
rect 29426 47302 29436 47354
rect 29460 47302 29490 47354
rect 29490 47302 29516 47354
rect 29220 47300 29276 47302
rect 29300 47300 29356 47302
rect 29380 47300 29436 47302
rect 29460 47300 29516 47302
rect 29220 46266 29276 46268
rect 29300 46266 29356 46268
rect 29380 46266 29436 46268
rect 29460 46266 29516 46268
rect 29220 46214 29246 46266
rect 29246 46214 29276 46266
rect 29300 46214 29310 46266
rect 29310 46214 29356 46266
rect 29380 46214 29426 46266
rect 29426 46214 29436 46266
rect 29460 46214 29490 46266
rect 29490 46214 29516 46266
rect 29220 46212 29276 46214
rect 29300 46212 29356 46214
rect 29380 46212 29436 46214
rect 29460 46212 29516 46214
rect 29220 45178 29276 45180
rect 29300 45178 29356 45180
rect 29380 45178 29436 45180
rect 29460 45178 29516 45180
rect 29220 45126 29246 45178
rect 29246 45126 29276 45178
rect 29300 45126 29310 45178
rect 29310 45126 29356 45178
rect 29380 45126 29426 45178
rect 29426 45126 29436 45178
rect 29460 45126 29490 45178
rect 29490 45126 29516 45178
rect 29220 45124 29276 45126
rect 29300 45124 29356 45126
rect 29380 45124 29436 45126
rect 29460 45124 29516 45126
rect 29220 44090 29276 44092
rect 29300 44090 29356 44092
rect 29380 44090 29436 44092
rect 29460 44090 29516 44092
rect 29220 44038 29246 44090
rect 29246 44038 29276 44090
rect 29300 44038 29310 44090
rect 29310 44038 29356 44090
rect 29380 44038 29426 44090
rect 29426 44038 29436 44090
rect 29460 44038 29490 44090
rect 29490 44038 29516 44090
rect 29220 44036 29276 44038
rect 29300 44036 29356 44038
rect 29380 44036 29436 44038
rect 29460 44036 29516 44038
rect 29220 43002 29276 43004
rect 29300 43002 29356 43004
rect 29380 43002 29436 43004
rect 29460 43002 29516 43004
rect 29220 42950 29246 43002
rect 29246 42950 29276 43002
rect 29300 42950 29310 43002
rect 29310 42950 29356 43002
rect 29380 42950 29426 43002
rect 29426 42950 29436 43002
rect 29460 42950 29490 43002
rect 29490 42950 29516 43002
rect 29220 42948 29276 42950
rect 29300 42948 29356 42950
rect 29380 42948 29436 42950
rect 29460 42948 29516 42950
rect 29220 41914 29276 41916
rect 29300 41914 29356 41916
rect 29380 41914 29436 41916
rect 29460 41914 29516 41916
rect 29220 41862 29246 41914
rect 29246 41862 29276 41914
rect 29300 41862 29310 41914
rect 29310 41862 29356 41914
rect 29380 41862 29426 41914
rect 29426 41862 29436 41914
rect 29460 41862 29490 41914
rect 29490 41862 29516 41914
rect 29220 41860 29276 41862
rect 29300 41860 29356 41862
rect 29380 41860 29436 41862
rect 29460 41860 29516 41862
rect 29220 40826 29276 40828
rect 29300 40826 29356 40828
rect 29380 40826 29436 40828
rect 29460 40826 29516 40828
rect 29220 40774 29246 40826
rect 29246 40774 29276 40826
rect 29300 40774 29310 40826
rect 29310 40774 29356 40826
rect 29380 40774 29426 40826
rect 29426 40774 29436 40826
rect 29460 40774 29490 40826
rect 29490 40774 29516 40826
rect 29220 40772 29276 40774
rect 29300 40772 29356 40774
rect 29380 40772 29436 40774
rect 29460 40772 29516 40774
rect 29220 39738 29276 39740
rect 29300 39738 29356 39740
rect 29380 39738 29436 39740
rect 29460 39738 29516 39740
rect 29220 39686 29246 39738
rect 29246 39686 29276 39738
rect 29300 39686 29310 39738
rect 29310 39686 29356 39738
rect 29380 39686 29426 39738
rect 29426 39686 29436 39738
rect 29460 39686 29490 39738
rect 29490 39686 29516 39738
rect 29220 39684 29276 39686
rect 29300 39684 29356 39686
rect 29380 39684 29436 39686
rect 29460 39684 29516 39686
rect 29220 38650 29276 38652
rect 29300 38650 29356 38652
rect 29380 38650 29436 38652
rect 29460 38650 29516 38652
rect 29220 38598 29246 38650
rect 29246 38598 29276 38650
rect 29300 38598 29310 38650
rect 29310 38598 29356 38650
rect 29380 38598 29426 38650
rect 29426 38598 29436 38650
rect 29460 38598 29490 38650
rect 29490 38598 29516 38650
rect 29220 38596 29276 38598
rect 29300 38596 29356 38598
rect 29380 38596 29436 38598
rect 29460 38596 29516 38598
rect 29220 37562 29276 37564
rect 29300 37562 29356 37564
rect 29380 37562 29436 37564
rect 29460 37562 29516 37564
rect 29220 37510 29246 37562
rect 29246 37510 29276 37562
rect 29300 37510 29310 37562
rect 29310 37510 29356 37562
rect 29380 37510 29426 37562
rect 29426 37510 29436 37562
rect 29460 37510 29490 37562
rect 29490 37510 29516 37562
rect 29220 37508 29276 37510
rect 29300 37508 29356 37510
rect 29380 37508 29436 37510
rect 29460 37508 29516 37510
rect 29220 36474 29276 36476
rect 29300 36474 29356 36476
rect 29380 36474 29436 36476
rect 29460 36474 29516 36476
rect 29220 36422 29246 36474
rect 29246 36422 29276 36474
rect 29300 36422 29310 36474
rect 29310 36422 29356 36474
rect 29380 36422 29426 36474
rect 29426 36422 29436 36474
rect 29460 36422 29490 36474
rect 29490 36422 29516 36474
rect 29220 36420 29276 36422
rect 29300 36420 29356 36422
rect 29380 36420 29436 36422
rect 29460 36420 29516 36422
rect 29220 35386 29276 35388
rect 29300 35386 29356 35388
rect 29380 35386 29436 35388
rect 29460 35386 29516 35388
rect 29220 35334 29246 35386
rect 29246 35334 29276 35386
rect 29300 35334 29310 35386
rect 29310 35334 29356 35386
rect 29380 35334 29426 35386
rect 29426 35334 29436 35386
rect 29460 35334 29490 35386
rect 29490 35334 29516 35386
rect 29220 35332 29276 35334
rect 29300 35332 29356 35334
rect 29380 35332 29436 35334
rect 29460 35332 29516 35334
rect 29220 34298 29276 34300
rect 29300 34298 29356 34300
rect 29380 34298 29436 34300
rect 29460 34298 29516 34300
rect 29220 34246 29246 34298
rect 29246 34246 29276 34298
rect 29300 34246 29310 34298
rect 29310 34246 29356 34298
rect 29380 34246 29426 34298
rect 29426 34246 29436 34298
rect 29460 34246 29490 34298
rect 29490 34246 29516 34298
rect 29220 34244 29276 34246
rect 29300 34244 29356 34246
rect 29380 34244 29436 34246
rect 29460 34244 29516 34246
rect 29220 33210 29276 33212
rect 29300 33210 29356 33212
rect 29380 33210 29436 33212
rect 29460 33210 29516 33212
rect 29220 33158 29246 33210
rect 29246 33158 29276 33210
rect 29300 33158 29310 33210
rect 29310 33158 29356 33210
rect 29380 33158 29426 33210
rect 29426 33158 29436 33210
rect 29460 33158 29490 33210
rect 29490 33158 29516 33210
rect 29220 33156 29276 33158
rect 29300 33156 29356 33158
rect 29380 33156 29436 33158
rect 29460 33156 29516 33158
rect 29220 32122 29276 32124
rect 29300 32122 29356 32124
rect 29380 32122 29436 32124
rect 29460 32122 29516 32124
rect 29220 32070 29246 32122
rect 29246 32070 29276 32122
rect 29300 32070 29310 32122
rect 29310 32070 29356 32122
rect 29380 32070 29426 32122
rect 29426 32070 29436 32122
rect 29460 32070 29490 32122
rect 29490 32070 29516 32122
rect 29220 32068 29276 32070
rect 29300 32068 29356 32070
rect 29380 32068 29436 32070
rect 29460 32068 29516 32070
rect 29220 31034 29276 31036
rect 29300 31034 29356 31036
rect 29380 31034 29436 31036
rect 29460 31034 29516 31036
rect 29220 30982 29246 31034
rect 29246 30982 29276 31034
rect 29300 30982 29310 31034
rect 29310 30982 29356 31034
rect 29380 30982 29426 31034
rect 29426 30982 29436 31034
rect 29460 30982 29490 31034
rect 29490 30982 29516 31034
rect 29220 30980 29276 30982
rect 29300 30980 29356 30982
rect 29380 30980 29436 30982
rect 29460 30980 29516 30982
rect 29220 29946 29276 29948
rect 29300 29946 29356 29948
rect 29380 29946 29436 29948
rect 29460 29946 29516 29948
rect 29220 29894 29246 29946
rect 29246 29894 29276 29946
rect 29300 29894 29310 29946
rect 29310 29894 29356 29946
rect 29380 29894 29426 29946
rect 29426 29894 29436 29946
rect 29460 29894 29490 29946
rect 29490 29894 29516 29946
rect 29220 29892 29276 29894
rect 29300 29892 29356 29894
rect 29380 29892 29436 29894
rect 29460 29892 29516 29894
rect 29220 28858 29276 28860
rect 29300 28858 29356 28860
rect 29380 28858 29436 28860
rect 29460 28858 29516 28860
rect 29220 28806 29246 28858
rect 29246 28806 29276 28858
rect 29300 28806 29310 28858
rect 29310 28806 29356 28858
rect 29380 28806 29426 28858
rect 29426 28806 29436 28858
rect 29460 28806 29490 28858
rect 29490 28806 29516 28858
rect 29220 28804 29276 28806
rect 29300 28804 29356 28806
rect 29380 28804 29436 28806
rect 29460 28804 29516 28806
rect 29220 27770 29276 27772
rect 29300 27770 29356 27772
rect 29380 27770 29436 27772
rect 29460 27770 29516 27772
rect 29220 27718 29246 27770
rect 29246 27718 29276 27770
rect 29300 27718 29310 27770
rect 29310 27718 29356 27770
rect 29380 27718 29426 27770
rect 29426 27718 29436 27770
rect 29460 27718 29490 27770
rect 29490 27718 29516 27770
rect 29220 27716 29276 27718
rect 29300 27716 29356 27718
rect 29380 27716 29436 27718
rect 29460 27716 29516 27718
rect 29220 26682 29276 26684
rect 29300 26682 29356 26684
rect 29380 26682 29436 26684
rect 29460 26682 29516 26684
rect 29220 26630 29246 26682
rect 29246 26630 29276 26682
rect 29300 26630 29310 26682
rect 29310 26630 29356 26682
rect 29380 26630 29426 26682
rect 29426 26630 29436 26682
rect 29460 26630 29490 26682
rect 29490 26630 29516 26682
rect 29220 26628 29276 26630
rect 29300 26628 29356 26630
rect 29380 26628 29436 26630
rect 29460 26628 29516 26630
rect 29220 25594 29276 25596
rect 29300 25594 29356 25596
rect 29380 25594 29436 25596
rect 29460 25594 29516 25596
rect 29220 25542 29246 25594
rect 29246 25542 29276 25594
rect 29300 25542 29310 25594
rect 29310 25542 29356 25594
rect 29380 25542 29426 25594
rect 29426 25542 29436 25594
rect 29460 25542 29490 25594
rect 29490 25542 29516 25594
rect 29220 25540 29276 25542
rect 29300 25540 29356 25542
rect 29380 25540 29436 25542
rect 29460 25540 29516 25542
rect 29220 24506 29276 24508
rect 29300 24506 29356 24508
rect 29380 24506 29436 24508
rect 29460 24506 29516 24508
rect 29220 24454 29246 24506
rect 29246 24454 29276 24506
rect 29300 24454 29310 24506
rect 29310 24454 29356 24506
rect 29380 24454 29426 24506
rect 29426 24454 29436 24506
rect 29460 24454 29490 24506
rect 29490 24454 29516 24506
rect 29220 24452 29276 24454
rect 29300 24452 29356 24454
rect 29380 24452 29436 24454
rect 29460 24452 29516 24454
rect 29220 23418 29276 23420
rect 29300 23418 29356 23420
rect 29380 23418 29436 23420
rect 29460 23418 29516 23420
rect 29220 23366 29246 23418
rect 29246 23366 29276 23418
rect 29300 23366 29310 23418
rect 29310 23366 29356 23418
rect 29380 23366 29426 23418
rect 29426 23366 29436 23418
rect 29460 23366 29490 23418
rect 29490 23366 29516 23418
rect 29220 23364 29276 23366
rect 29300 23364 29356 23366
rect 29380 23364 29436 23366
rect 29460 23364 29516 23366
rect 29220 22330 29276 22332
rect 29300 22330 29356 22332
rect 29380 22330 29436 22332
rect 29460 22330 29516 22332
rect 29220 22278 29246 22330
rect 29246 22278 29276 22330
rect 29300 22278 29310 22330
rect 29310 22278 29356 22330
rect 29380 22278 29426 22330
rect 29426 22278 29436 22330
rect 29460 22278 29490 22330
rect 29490 22278 29516 22330
rect 29220 22276 29276 22278
rect 29300 22276 29356 22278
rect 29380 22276 29436 22278
rect 29460 22276 29516 22278
rect 29220 21242 29276 21244
rect 29300 21242 29356 21244
rect 29380 21242 29436 21244
rect 29460 21242 29516 21244
rect 29220 21190 29246 21242
rect 29246 21190 29276 21242
rect 29300 21190 29310 21242
rect 29310 21190 29356 21242
rect 29380 21190 29426 21242
rect 29426 21190 29436 21242
rect 29460 21190 29490 21242
rect 29490 21190 29516 21242
rect 29220 21188 29276 21190
rect 29300 21188 29356 21190
rect 29380 21188 29436 21190
rect 29460 21188 29516 21190
rect 29220 20154 29276 20156
rect 29300 20154 29356 20156
rect 29380 20154 29436 20156
rect 29460 20154 29516 20156
rect 29220 20102 29246 20154
rect 29246 20102 29276 20154
rect 29300 20102 29310 20154
rect 29310 20102 29356 20154
rect 29380 20102 29426 20154
rect 29426 20102 29436 20154
rect 29460 20102 29490 20154
rect 29490 20102 29516 20154
rect 29220 20100 29276 20102
rect 29300 20100 29356 20102
rect 29380 20100 29436 20102
rect 29460 20100 29516 20102
rect 32770 34604 32826 34640
rect 32770 34584 32772 34604
rect 32772 34584 32824 34604
rect 32824 34584 32826 34604
rect 34220 66394 34276 66396
rect 34300 66394 34356 66396
rect 34380 66394 34436 66396
rect 34460 66394 34516 66396
rect 34220 66342 34246 66394
rect 34246 66342 34276 66394
rect 34300 66342 34310 66394
rect 34310 66342 34356 66394
rect 34380 66342 34426 66394
rect 34426 66342 34436 66394
rect 34460 66342 34490 66394
rect 34490 66342 34516 66394
rect 34220 66340 34276 66342
rect 34300 66340 34356 66342
rect 34380 66340 34436 66342
rect 34460 66340 34516 66342
rect 34220 65306 34276 65308
rect 34300 65306 34356 65308
rect 34380 65306 34436 65308
rect 34460 65306 34516 65308
rect 34220 65254 34246 65306
rect 34246 65254 34276 65306
rect 34300 65254 34310 65306
rect 34310 65254 34356 65306
rect 34380 65254 34426 65306
rect 34426 65254 34436 65306
rect 34460 65254 34490 65306
rect 34490 65254 34516 65306
rect 34220 65252 34276 65254
rect 34300 65252 34356 65254
rect 34380 65252 34436 65254
rect 34460 65252 34516 65254
rect 34220 64218 34276 64220
rect 34300 64218 34356 64220
rect 34380 64218 34436 64220
rect 34460 64218 34516 64220
rect 34220 64166 34246 64218
rect 34246 64166 34276 64218
rect 34300 64166 34310 64218
rect 34310 64166 34356 64218
rect 34380 64166 34426 64218
rect 34426 64166 34436 64218
rect 34460 64166 34490 64218
rect 34490 64166 34516 64218
rect 34220 64164 34276 64166
rect 34300 64164 34356 64166
rect 34380 64164 34436 64166
rect 34460 64164 34516 64166
rect 34220 63130 34276 63132
rect 34300 63130 34356 63132
rect 34380 63130 34436 63132
rect 34460 63130 34516 63132
rect 34220 63078 34246 63130
rect 34246 63078 34276 63130
rect 34300 63078 34310 63130
rect 34310 63078 34356 63130
rect 34380 63078 34426 63130
rect 34426 63078 34436 63130
rect 34460 63078 34490 63130
rect 34490 63078 34516 63130
rect 34220 63076 34276 63078
rect 34300 63076 34356 63078
rect 34380 63076 34436 63078
rect 34460 63076 34516 63078
rect 34220 62042 34276 62044
rect 34300 62042 34356 62044
rect 34380 62042 34436 62044
rect 34460 62042 34516 62044
rect 34220 61990 34246 62042
rect 34246 61990 34276 62042
rect 34300 61990 34310 62042
rect 34310 61990 34356 62042
rect 34380 61990 34426 62042
rect 34426 61990 34436 62042
rect 34460 61990 34490 62042
rect 34490 61990 34516 62042
rect 34220 61988 34276 61990
rect 34300 61988 34356 61990
rect 34380 61988 34436 61990
rect 34460 61988 34516 61990
rect 34220 60954 34276 60956
rect 34300 60954 34356 60956
rect 34380 60954 34436 60956
rect 34460 60954 34516 60956
rect 34220 60902 34246 60954
rect 34246 60902 34276 60954
rect 34300 60902 34310 60954
rect 34310 60902 34356 60954
rect 34380 60902 34426 60954
rect 34426 60902 34436 60954
rect 34460 60902 34490 60954
rect 34490 60902 34516 60954
rect 34220 60900 34276 60902
rect 34300 60900 34356 60902
rect 34380 60900 34436 60902
rect 34460 60900 34516 60902
rect 34220 59866 34276 59868
rect 34300 59866 34356 59868
rect 34380 59866 34436 59868
rect 34460 59866 34516 59868
rect 34220 59814 34246 59866
rect 34246 59814 34276 59866
rect 34300 59814 34310 59866
rect 34310 59814 34356 59866
rect 34380 59814 34426 59866
rect 34426 59814 34436 59866
rect 34460 59814 34490 59866
rect 34490 59814 34516 59866
rect 34220 59812 34276 59814
rect 34300 59812 34356 59814
rect 34380 59812 34436 59814
rect 34460 59812 34516 59814
rect 34220 58778 34276 58780
rect 34300 58778 34356 58780
rect 34380 58778 34436 58780
rect 34460 58778 34516 58780
rect 34220 58726 34246 58778
rect 34246 58726 34276 58778
rect 34300 58726 34310 58778
rect 34310 58726 34356 58778
rect 34380 58726 34426 58778
rect 34426 58726 34436 58778
rect 34460 58726 34490 58778
rect 34490 58726 34516 58778
rect 34220 58724 34276 58726
rect 34300 58724 34356 58726
rect 34380 58724 34436 58726
rect 34460 58724 34516 58726
rect 34220 57690 34276 57692
rect 34300 57690 34356 57692
rect 34380 57690 34436 57692
rect 34460 57690 34516 57692
rect 34220 57638 34246 57690
rect 34246 57638 34276 57690
rect 34300 57638 34310 57690
rect 34310 57638 34356 57690
rect 34380 57638 34426 57690
rect 34426 57638 34436 57690
rect 34460 57638 34490 57690
rect 34490 57638 34516 57690
rect 34220 57636 34276 57638
rect 34300 57636 34356 57638
rect 34380 57636 34436 57638
rect 34460 57636 34516 57638
rect 34220 56602 34276 56604
rect 34300 56602 34356 56604
rect 34380 56602 34436 56604
rect 34460 56602 34516 56604
rect 34220 56550 34246 56602
rect 34246 56550 34276 56602
rect 34300 56550 34310 56602
rect 34310 56550 34356 56602
rect 34380 56550 34426 56602
rect 34426 56550 34436 56602
rect 34460 56550 34490 56602
rect 34490 56550 34516 56602
rect 34220 56548 34276 56550
rect 34300 56548 34356 56550
rect 34380 56548 34436 56550
rect 34460 56548 34516 56550
rect 34220 55514 34276 55516
rect 34300 55514 34356 55516
rect 34380 55514 34436 55516
rect 34460 55514 34516 55516
rect 34220 55462 34246 55514
rect 34246 55462 34276 55514
rect 34300 55462 34310 55514
rect 34310 55462 34356 55514
rect 34380 55462 34426 55514
rect 34426 55462 34436 55514
rect 34460 55462 34490 55514
rect 34490 55462 34516 55514
rect 34220 55460 34276 55462
rect 34300 55460 34356 55462
rect 34380 55460 34436 55462
rect 34460 55460 34516 55462
rect 34220 54426 34276 54428
rect 34300 54426 34356 54428
rect 34380 54426 34436 54428
rect 34460 54426 34516 54428
rect 34220 54374 34246 54426
rect 34246 54374 34276 54426
rect 34300 54374 34310 54426
rect 34310 54374 34356 54426
rect 34380 54374 34426 54426
rect 34426 54374 34436 54426
rect 34460 54374 34490 54426
rect 34490 54374 34516 54426
rect 34220 54372 34276 54374
rect 34300 54372 34356 54374
rect 34380 54372 34436 54374
rect 34460 54372 34516 54374
rect 34220 53338 34276 53340
rect 34300 53338 34356 53340
rect 34380 53338 34436 53340
rect 34460 53338 34516 53340
rect 34220 53286 34246 53338
rect 34246 53286 34276 53338
rect 34300 53286 34310 53338
rect 34310 53286 34356 53338
rect 34380 53286 34426 53338
rect 34426 53286 34436 53338
rect 34460 53286 34490 53338
rect 34490 53286 34516 53338
rect 34220 53284 34276 53286
rect 34300 53284 34356 53286
rect 34380 53284 34436 53286
rect 34460 53284 34516 53286
rect 34220 52250 34276 52252
rect 34300 52250 34356 52252
rect 34380 52250 34436 52252
rect 34460 52250 34516 52252
rect 34220 52198 34246 52250
rect 34246 52198 34276 52250
rect 34300 52198 34310 52250
rect 34310 52198 34356 52250
rect 34380 52198 34426 52250
rect 34426 52198 34436 52250
rect 34460 52198 34490 52250
rect 34490 52198 34516 52250
rect 34220 52196 34276 52198
rect 34300 52196 34356 52198
rect 34380 52196 34436 52198
rect 34460 52196 34516 52198
rect 34220 51162 34276 51164
rect 34300 51162 34356 51164
rect 34380 51162 34436 51164
rect 34460 51162 34516 51164
rect 34220 51110 34246 51162
rect 34246 51110 34276 51162
rect 34300 51110 34310 51162
rect 34310 51110 34356 51162
rect 34380 51110 34426 51162
rect 34426 51110 34436 51162
rect 34460 51110 34490 51162
rect 34490 51110 34516 51162
rect 34220 51108 34276 51110
rect 34300 51108 34356 51110
rect 34380 51108 34436 51110
rect 34460 51108 34516 51110
rect 34220 50074 34276 50076
rect 34300 50074 34356 50076
rect 34380 50074 34436 50076
rect 34460 50074 34516 50076
rect 34220 50022 34246 50074
rect 34246 50022 34276 50074
rect 34300 50022 34310 50074
rect 34310 50022 34356 50074
rect 34380 50022 34426 50074
rect 34426 50022 34436 50074
rect 34460 50022 34490 50074
rect 34490 50022 34516 50074
rect 34220 50020 34276 50022
rect 34300 50020 34356 50022
rect 34380 50020 34436 50022
rect 34460 50020 34516 50022
rect 34220 48986 34276 48988
rect 34300 48986 34356 48988
rect 34380 48986 34436 48988
rect 34460 48986 34516 48988
rect 34220 48934 34246 48986
rect 34246 48934 34276 48986
rect 34300 48934 34310 48986
rect 34310 48934 34356 48986
rect 34380 48934 34426 48986
rect 34426 48934 34436 48986
rect 34460 48934 34490 48986
rect 34490 48934 34516 48986
rect 34220 48932 34276 48934
rect 34300 48932 34356 48934
rect 34380 48932 34436 48934
rect 34460 48932 34516 48934
rect 34220 47898 34276 47900
rect 34300 47898 34356 47900
rect 34380 47898 34436 47900
rect 34460 47898 34516 47900
rect 34220 47846 34246 47898
rect 34246 47846 34276 47898
rect 34300 47846 34310 47898
rect 34310 47846 34356 47898
rect 34380 47846 34426 47898
rect 34426 47846 34436 47898
rect 34460 47846 34490 47898
rect 34490 47846 34516 47898
rect 34220 47844 34276 47846
rect 34300 47844 34356 47846
rect 34380 47844 34436 47846
rect 34460 47844 34516 47846
rect 34220 46810 34276 46812
rect 34300 46810 34356 46812
rect 34380 46810 34436 46812
rect 34460 46810 34516 46812
rect 34220 46758 34246 46810
rect 34246 46758 34276 46810
rect 34300 46758 34310 46810
rect 34310 46758 34356 46810
rect 34380 46758 34426 46810
rect 34426 46758 34436 46810
rect 34460 46758 34490 46810
rect 34490 46758 34516 46810
rect 34220 46756 34276 46758
rect 34300 46756 34356 46758
rect 34380 46756 34436 46758
rect 34460 46756 34516 46758
rect 34220 45722 34276 45724
rect 34300 45722 34356 45724
rect 34380 45722 34436 45724
rect 34460 45722 34516 45724
rect 34220 45670 34246 45722
rect 34246 45670 34276 45722
rect 34300 45670 34310 45722
rect 34310 45670 34356 45722
rect 34380 45670 34426 45722
rect 34426 45670 34436 45722
rect 34460 45670 34490 45722
rect 34490 45670 34516 45722
rect 34220 45668 34276 45670
rect 34300 45668 34356 45670
rect 34380 45668 34436 45670
rect 34460 45668 34516 45670
rect 34220 44634 34276 44636
rect 34300 44634 34356 44636
rect 34380 44634 34436 44636
rect 34460 44634 34516 44636
rect 34220 44582 34246 44634
rect 34246 44582 34276 44634
rect 34300 44582 34310 44634
rect 34310 44582 34356 44634
rect 34380 44582 34426 44634
rect 34426 44582 34436 44634
rect 34460 44582 34490 44634
rect 34490 44582 34516 44634
rect 34220 44580 34276 44582
rect 34300 44580 34356 44582
rect 34380 44580 34436 44582
rect 34460 44580 34516 44582
rect 34220 43546 34276 43548
rect 34300 43546 34356 43548
rect 34380 43546 34436 43548
rect 34460 43546 34516 43548
rect 34220 43494 34246 43546
rect 34246 43494 34276 43546
rect 34300 43494 34310 43546
rect 34310 43494 34356 43546
rect 34380 43494 34426 43546
rect 34426 43494 34436 43546
rect 34460 43494 34490 43546
rect 34490 43494 34516 43546
rect 34220 43492 34276 43494
rect 34300 43492 34356 43494
rect 34380 43492 34436 43494
rect 34460 43492 34516 43494
rect 34220 42458 34276 42460
rect 34300 42458 34356 42460
rect 34380 42458 34436 42460
rect 34460 42458 34516 42460
rect 34220 42406 34246 42458
rect 34246 42406 34276 42458
rect 34300 42406 34310 42458
rect 34310 42406 34356 42458
rect 34380 42406 34426 42458
rect 34426 42406 34436 42458
rect 34460 42406 34490 42458
rect 34490 42406 34516 42458
rect 34220 42404 34276 42406
rect 34300 42404 34356 42406
rect 34380 42404 34436 42406
rect 34460 42404 34516 42406
rect 34220 41370 34276 41372
rect 34300 41370 34356 41372
rect 34380 41370 34436 41372
rect 34460 41370 34516 41372
rect 34220 41318 34246 41370
rect 34246 41318 34276 41370
rect 34300 41318 34310 41370
rect 34310 41318 34356 41370
rect 34380 41318 34426 41370
rect 34426 41318 34436 41370
rect 34460 41318 34490 41370
rect 34490 41318 34516 41370
rect 34220 41316 34276 41318
rect 34300 41316 34356 41318
rect 34380 41316 34436 41318
rect 34460 41316 34516 41318
rect 34220 40282 34276 40284
rect 34300 40282 34356 40284
rect 34380 40282 34436 40284
rect 34460 40282 34516 40284
rect 34220 40230 34246 40282
rect 34246 40230 34276 40282
rect 34300 40230 34310 40282
rect 34310 40230 34356 40282
rect 34380 40230 34426 40282
rect 34426 40230 34436 40282
rect 34460 40230 34490 40282
rect 34490 40230 34516 40282
rect 34220 40228 34276 40230
rect 34300 40228 34356 40230
rect 34380 40228 34436 40230
rect 34460 40228 34516 40230
rect 34220 39194 34276 39196
rect 34300 39194 34356 39196
rect 34380 39194 34436 39196
rect 34460 39194 34516 39196
rect 34220 39142 34246 39194
rect 34246 39142 34276 39194
rect 34300 39142 34310 39194
rect 34310 39142 34356 39194
rect 34380 39142 34426 39194
rect 34426 39142 34436 39194
rect 34460 39142 34490 39194
rect 34490 39142 34516 39194
rect 34220 39140 34276 39142
rect 34300 39140 34356 39142
rect 34380 39140 34436 39142
rect 34460 39140 34516 39142
rect 34220 38106 34276 38108
rect 34300 38106 34356 38108
rect 34380 38106 34436 38108
rect 34460 38106 34516 38108
rect 34220 38054 34246 38106
rect 34246 38054 34276 38106
rect 34300 38054 34310 38106
rect 34310 38054 34356 38106
rect 34380 38054 34426 38106
rect 34426 38054 34436 38106
rect 34460 38054 34490 38106
rect 34490 38054 34516 38106
rect 34220 38052 34276 38054
rect 34300 38052 34356 38054
rect 34380 38052 34436 38054
rect 34460 38052 34516 38054
rect 34220 37018 34276 37020
rect 34300 37018 34356 37020
rect 34380 37018 34436 37020
rect 34460 37018 34516 37020
rect 34220 36966 34246 37018
rect 34246 36966 34276 37018
rect 34300 36966 34310 37018
rect 34310 36966 34356 37018
rect 34380 36966 34426 37018
rect 34426 36966 34436 37018
rect 34460 36966 34490 37018
rect 34490 36966 34516 37018
rect 34220 36964 34276 36966
rect 34300 36964 34356 36966
rect 34380 36964 34436 36966
rect 34460 36964 34516 36966
rect 34220 35930 34276 35932
rect 34300 35930 34356 35932
rect 34380 35930 34436 35932
rect 34460 35930 34516 35932
rect 34220 35878 34246 35930
rect 34246 35878 34276 35930
rect 34300 35878 34310 35930
rect 34310 35878 34356 35930
rect 34380 35878 34426 35930
rect 34426 35878 34436 35930
rect 34460 35878 34490 35930
rect 34490 35878 34516 35930
rect 34220 35876 34276 35878
rect 34300 35876 34356 35878
rect 34380 35876 34436 35878
rect 34460 35876 34516 35878
rect 34220 34842 34276 34844
rect 34300 34842 34356 34844
rect 34380 34842 34436 34844
rect 34460 34842 34516 34844
rect 34220 34790 34246 34842
rect 34246 34790 34276 34842
rect 34300 34790 34310 34842
rect 34310 34790 34356 34842
rect 34380 34790 34426 34842
rect 34426 34790 34436 34842
rect 34460 34790 34490 34842
rect 34490 34790 34516 34842
rect 34220 34788 34276 34790
rect 34300 34788 34356 34790
rect 34380 34788 34436 34790
rect 34460 34788 34516 34790
rect 33874 34604 33930 34640
rect 33874 34584 33876 34604
rect 33876 34584 33928 34604
rect 33928 34584 33930 34604
rect 34220 33754 34276 33756
rect 34300 33754 34356 33756
rect 34380 33754 34436 33756
rect 34460 33754 34516 33756
rect 34220 33702 34246 33754
rect 34246 33702 34276 33754
rect 34300 33702 34310 33754
rect 34310 33702 34356 33754
rect 34380 33702 34426 33754
rect 34426 33702 34436 33754
rect 34460 33702 34490 33754
rect 34490 33702 34516 33754
rect 34220 33700 34276 33702
rect 34300 33700 34356 33702
rect 34380 33700 34436 33702
rect 34460 33700 34516 33702
rect 34220 32666 34276 32668
rect 34300 32666 34356 32668
rect 34380 32666 34436 32668
rect 34460 32666 34516 32668
rect 34220 32614 34246 32666
rect 34246 32614 34276 32666
rect 34300 32614 34310 32666
rect 34310 32614 34356 32666
rect 34380 32614 34426 32666
rect 34426 32614 34436 32666
rect 34460 32614 34490 32666
rect 34490 32614 34516 32666
rect 34220 32612 34276 32614
rect 34300 32612 34356 32614
rect 34380 32612 34436 32614
rect 34460 32612 34516 32614
rect 34220 31578 34276 31580
rect 34300 31578 34356 31580
rect 34380 31578 34436 31580
rect 34460 31578 34516 31580
rect 34220 31526 34246 31578
rect 34246 31526 34276 31578
rect 34300 31526 34310 31578
rect 34310 31526 34356 31578
rect 34380 31526 34426 31578
rect 34426 31526 34436 31578
rect 34460 31526 34490 31578
rect 34490 31526 34516 31578
rect 34220 31524 34276 31526
rect 34300 31524 34356 31526
rect 34380 31524 34436 31526
rect 34460 31524 34516 31526
rect 34220 30490 34276 30492
rect 34300 30490 34356 30492
rect 34380 30490 34436 30492
rect 34460 30490 34516 30492
rect 34220 30438 34246 30490
rect 34246 30438 34276 30490
rect 34300 30438 34310 30490
rect 34310 30438 34356 30490
rect 34380 30438 34426 30490
rect 34426 30438 34436 30490
rect 34460 30438 34490 30490
rect 34490 30438 34516 30490
rect 34220 30436 34276 30438
rect 34300 30436 34356 30438
rect 34380 30436 34436 30438
rect 34460 30436 34516 30438
rect 34220 29402 34276 29404
rect 34300 29402 34356 29404
rect 34380 29402 34436 29404
rect 34460 29402 34516 29404
rect 34220 29350 34246 29402
rect 34246 29350 34276 29402
rect 34300 29350 34310 29402
rect 34310 29350 34356 29402
rect 34380 29350 34426 29402
rect 34426 29350 34436 29402
rect 34460 29350 34490 29402
rect 34490 29350 34516 29402
rect 34220 29348 34276 29350
rect 34300 29348 34356 29350
rect 34380 29348 34436 29350
rect 34460 29348 34516 29350
rect 34220 28314 34276 28316
rect 34300 28314 34356 28316
rect 34380 28314 34436 28316
rect 34460 28314 34516 28316
rect 34220 28262 34246 28314
rect 34246 28262 34276 28314
rect 34300 28262 34310 28314
rect 34310 28262 34356 28314
rect 34380 28262 34426 28314
rect 34426 28262 34436 28314
rect 34460 28262 34490 28314
rect 34490 28262 34516 28314
rect 34220 28260 34276 28262
rect 34300 28260 34356 28262
rect 34380 28260 34436 28262
rect 34460 28260 34516 28262
rect 34220 27226 34276 27228
rect 34300 27226 34356 27228
rect 34380 27226 34436 27228
rect 34460 27226 34516 27228
rect 34220 27174 34246 27226
rect 34246 27174 34276 27226
rect 34300 27174 34310 27226
rect 34310 27174 34356 27226
rect 34380 27174 34426 27226
rect 34426 27174 34436 27226
rect 34460 27174 34490 27226
rect 34490 27174 34516 27226
rect 34220 27172 34276 27174
rect 34300 27172 34356 27174
rect 34380 27172 34436 27174
rect 34460 27172 34516 27174
rect 34220 26138 34276 26140
rect 34300 26138 34356 26140
rect 34380 26138 34436 26140
rect 34460 26138 34516 26140
rect 34220 26086 34246 26138
rect 34246 26086 34276 26138
rect 34300 26086 34310 26138
rect 34310 26086 34356 26138
rect 34380 26086 34426 26138
rect 34426 26086 34436 26138
rect 34460 26086 34490 26138
rect 34490 26086 34516 26138
rect 34220 26084 34276 26086
rect 34300 26084 34356 26086
rect 34380 26084 34436 26086
rect 34460 26084 34516 26086
rect 34220 25050 34276 25052
rect 34300 25050 34356 25052
rect 34380 25050 34436 25052
rect 34460 25050 34516 25052
rect 34220 24998 34246 25050
rect 34246 24998 34276 25050
rect 34300 24998 34310 25050
rect 34310 24998 34356 25050
rect 34380 24998 34426 25050
rect 34426 24998 34436 25050
rect 34460 24998 34490 25050
rect 34490 24998 34516 25050
rect 34220 24996 34276 24998
rect 34300 24996 34356 24998
rect 34380 24996 34436 24998
rect 34460 24996 34516 24998
rect 34220 23962 34276 23964
rect 34300 23962 34356 23964
rect 34380 23962 34436 23964
rect 34460 23962 34516 23964
rect 34220 23910 34246 23962
rect 34246 23910 34276 23962
rect 34300 23910 34310 23962
rect 34310 23910 34356 23962
rect 34380 23910 34426 23962
rect 34426 23910 34436 23962
rect 34460 23910 34490 23962
rect 34490 23910 34516 23962
rect 34220 23908 34276 23910
rect 34300 23908 34356 23910
rect 34380 23908 34436 23910
rect 34460 23908 34516 23910
rect 34220 22874 34276 22876
rect 34300 22874 34356 22876
rect 34380 22874 34436 22876
rect 34460 22874 34516 22876
rect 34220 22822 34246 22874
rect 34246 22822 34276 22874
rect 34300 22822 34310 22874
rect 34310 22822 34356 22874
rect 34380 22822 34426 22874
rect 34426 22822 34436 22874
rect 34460 22822 34490 22874
rect 34490 22822 34516 22874
rect 34220 22820 34276 22822
rect 34300 22820 34356 22822
rect 34380 22820 34436 22822
rect 34460 22820 34516 22822
rect 34220 21786 34276 21788
rect 34300 21786 34356 21788
rect 34380 21786 34436 21788
rect 34460 21786 34516 21788
rect 34220 21734 34246 21786
rect 34246 21734 34276 21786
rect 34300 21734 34310 21786
rect 34310 21734 34356 21786
rect 34380 21734 34426 21786
rect 34426 21734 34436 21786
rect 34460 21734 34490 21786
rect 34490 21734 34516 21786
rect 34220 21732 34276 21734
rect 34300 21732 34356 21734
rect 34380 21732 34436 21734
rect 34460 21732 34516 21734
rect 34220 20698 34276 20700
rect 34300 20698 34356 20700
rect 34380 20698 34436 20700
rect 34460 20698 34516 20700
rect 34220 20646 34246 20698
rect 34246 20646 34276 20698
rect 34300 20646 34310 20698
rect 34310 20646 34356 20698
rect 34380 20646 34426 20698
rect 34426 20646 34436 20698
rect 34460 20646 34490 20698
rect 34490 20646 34516 20698
rect 34220 20644 34276 20646
rect 34300 20644 34356 20646
rect 34380 20644 34436 20646
rect 34460 20644 34516 20646
rect 34220 19610 34276 19612
rect 34300 19610 34356 19612
rect 34380 19610 34436 19612
rect 34460 19610 34516 19612
rect 34220 19558 34246 19610
rect 34246 19558 34276 19610
rect 34300 19558 34310 19610
rect 34310 19558 34356 19610
rect 34380 19558 34426 19610
rect 34426 19558 34436 19610
rect 34460 19558 34490 19610
rect 34490 19558 34516 19610
rect 34220 19556 34276 19558
rect 34300 19556 34356 19558
rect 34380 19556 34436 19558
rect 34460 19556 34516 19558
rect 39220 66938 39276 66940
rect 39300 66938 39356 66940
rect 39380 66938 39436 66940
rect 39460 66938 39516 66940
rect 39220 66886 39246 66938
rect 39246 66886 39276 66938
rect 39300 66886 39310 66938
rect 39310 66886 39356 66938
rect 39380 66886 39426 66938
rect 39426 66886 39436 66938
rect 39460 66886 39490 66938
rect 39490 66886 39516 66938
rect 39220 66884 39276 66886
rect 39300 66884 39356 66886
rect 39380 66884 39436 66886
rect 39460 66884 39516 66886
rect 49220 66938 49276 66940
rect 49300 66938 49356 66940
rect 49380 66938 49436 66940
rect 49460 66938 49516 66940
rect 49220 66886 49246 66938
rect 49246 66886 49276 66938
rect 49300 66886 49310 66938
rect 49310 66886 49356 66938
rect 49380 66886 49426 66938
rect 49426 66886 49436 66938
rect 49460 66886 49490 66938
rect 49490 66886 49516 66938
rect 49220 66884 49276 66886
rect 49300 66884 49356 66886
rect 49380 66884 49436 66886
rect 49460 66884 49516 66886
rect 39220 65850 39276 65852
rect 39300 65850 39356 65852
rect 39380 65850 39436 65852
rect 39460 65850 39516 65852
rect 39220 65798 39246 65850
rect 39246 65798 39276 65850
rect 39300 65798 39310 65850
rect 39310 65798 39356 65850
rect 39380 65798 39426 65850
rect 39426 65798 39436 65850
rect 39460 65798 39490 65850
rect 39490 65798 39516 65850
rect 39220 65796 39276 65798
rect 39300 65796 39356 65798
rect 39380 65796 39436 65798
rect 39460 65796 39516 65798
rect 39220 64762 39276 64764
rect 39300 64762 39356 64764
rect 39380 64762 39436 64764
rect 39460 64762 39516 64764
rect 39220 64710 39246 64762
rect 39246 64710 39276 64762
rect 39300 64710 39310 64762
rect 39310 64710 39356 64762
rect 39380 64710 39426 64762
rect 39426 64710 39436 64762
rect 39460 64710 39490 64762
rect 39490 64710 39516 64762
rect 39220 64708 39276 64710
rect 39300 64708 39356 64710
rect 39380 64708 39436 64710
rect 39460 64708 39516 64710
rect 18786 6296 18842 6352
rect 18878 5752 18934 5808
rect 18878 2896 18934 2952
rect 18878 2760 18934 2816
rect 18878 2624 18934 2680
rect 19062 3304 19118 3360
rect 19154 2896 19210 2952
rect 21178 5616 21234 5672
rect 21638 3848 21694 3904
rect 22650 3712 22706 3768
rect 23478 5888 23534 5944
rect 23938 6160 23994 6216
rect 23938 6024 23994 6080
rect 24122 4800 24178 4856
rect 27710 1808 27766 1864
rect 28078 1808 28134 1864
rect 28170 1672 28226 1728
rect 28906 1672 28962 1728
rect 29918 1808 29974 1864
rect 30194 1808 30250 1864
rect 31022 1808 31078 1864
rect 31850 3440 31906 3496
rect 31850 1128 31906 1184
rect 32402 3848 32458 3904
rect 32770 3576 32826 3632
rect 33138 5752 33194 5808
rect 33046 5072 33102 5128
rect 33046 3576 33102 3632
rect 33966 3732 34022 3768
rect 33966 3712 33968 3732
rect 33968 3712 34020 3732
rect 34020 3712 34022 3732
rect 33874 3304 33930 3360
rect 34702 3188 34758 3224
rect 34702 3168 34704 3188
rect 34704 3168 34756 3188
rect 34756 3168 34758 3188
rect 34702 2760 34758 2816
rect 35162 6840 35218 6896
rect 35070 2760 35126 2816
rect 35990 3712 36046 3768
rect 35990 3032 36046 3088
rect 36726 6432 36782 6488
rect 36634 2352 36690 2408
rect 37922 12144 37978 12200
rect 39220 63674 39276 63676
rect 39300 63674 39356 63676
rect 39380 63674 39436 63676
rect 39460 63674 39516 63676
rect 39220 63622 39246 63674
rect 39246 63622 39276 63674
rect 39300 63622 39310 63674
rect 39310 63622 39356 63674
rect 39380 63622 39426 63674
rect 39426 63622 39436 63674
rect 39460 63622 39490 63674
rect 39490 63622 39516 63674
rect 39220 63620 39276 63622
rect 39300 63620 39356 63622
rect 39380 63620 39436 63622
rect 39460 63620 39516 63622
rect 39220 62586 39276 62588
rect 39300 62586 39356 62588
rect 39380 62586 39436 62588
rect 39460 62586 39516 62588
rect 39220 62534 39246 62586
rect 39246 62534 39276 62586
rect 39300 62534 39310 62586
rect 39310 62534 39356 62586
rect 39380 62534 39426 62586
rect 39426 62534 39436 62586
rect 39460 62534 39490 62586
rect 39490 62534 39516 62586
rect 39220 62532 39276 62534
rect 39300 62532 39356 62534
rect 39380 62532 39436 62534
rect 39460 62532 39516 62534
rect 39220 61498 39276 61500
rect 39300 61498 39356 61500
rect 39380 61498 39436 61500
rect 39460 61498 39516 61500
rect 39220 61446 39246 61498
rect 39246 61446 39276 61498
rect 39300 61446 39310 61498
rect 39310 61446 39356 61498
rect 39380 61446 39426 61498
rect 39426 61446 39436 61498
rect 39460 61446 39490 61498
rect 39490 61446 39516 61498
rect 39220 61444 39276 61446
rect 39300 61444 39356 61446
rect 39380 61444 39436 61446
rect 39460 61444 39516 61446
rect 39220 60410 39276 60412
rect 39300 60410 39356 60412
rect 39380 60410 39436 60412
rect 39460 60410 39516 60412
rect 39220 60358 39246 60410
rect 39246 60358 39276 60410
rect 39300 60358 39310 60410
rect 39310 60358 39356 60410
rect 39380 60358 39426 60410
rect 39426 60358 39436 60410
rect 39460 60358 39490 60410
rect 39490 60358 39516 60410
rect 39220 60356 39276 60358
rect 39300 60356 39356 60358
rect 39380 60356 39436 60358
rect 39460 60356 39516 60358
rect 39220 59322 39276 59324
rect 39300 59322 39356 59324
rect 39380 59322 39436 59324
rect 39460 59322 39516 59324
rect 39220 59270 39246 59322
rect 39246 59270 39276 59322
rect 39300 59270 39310 59322
rect 39310 59270 39356 59322
rect 39380 59270 39426 59322
rect 39426 59270 39436 59322
rect 39460 59270 39490 59322
rect 39490 59270 39516 59322
rect 39220 59268 39276 59270
rect 39300 59268 39356 59270
rect 39380 59268 39436 59270
rect 39460 59268 39516 59270
rect 39220 58234 39276 58236
rect 39300 58234 39356 58236
rect 39380 58234 39436 58236
rect 39460 58234 39516 58236
rect 39220 58182 39246 58234
rect 39246 58182 39276 58234
rect 39300 58182 39310 58234
rect 39310 58182 39356 58234
rect 39380 58182 39426 58234
rect 39426 58182 39436 58234
rect 39460 58182 39490 58234
rect 39490 58182 39516 58234
rect 39220 58180 39276 58182
rect 39300 58180 39356 58182
rect 39380 58180 39436 58182
rect 39460 58180 39516 58182
rect 39220 57146 39276 57148
rect 39300 57146 39356 57148
rect 39380 57146 39436 57148
rect 39460 57146 39516 57148
rect 39220 57094 39246 57146
rect 39246 57094 39276 57146
rect 39300 57094 39310 57146
rect 39310 57094 39356 57146
rect 39380 57094 39426 57146
rect 39426 57094 39436 57146
rect 39460 57094 39490 57146
rect 39490 57094 39516 57146
rect 39220 57092 39276 57094
rect 39300 57092 39356 57094
rect 39380 57092 39436 57094
rect 39460 57092 39516 57094
rect 39220 56058 39276 56060
rect 39300 56058 39356 56060
rect 39380 56058 39436 56060
rect 39460 56058 39516 56060
rect 39220 56006 39246 56058
rect 39246 56006 39276 56058
rect 39300 56006 39310 56058
rect 39310 56006 39356 56058
rect 39380 56006 39426 56058
rect 39426 56006 39436 56058
rect 39460 56006 39490 56058
rect 39490 56006 39516 56058
rect 39220 56004 39276 56006
rect 39300 56004 39356 56006
rect 39380 56004 39436 56006
rect 39460 56004 39516 56006
rect 39220 54970 39276 54972
rect 39300 54970 39356 54972
rect 39380 54970 39436 54972
rect 39460 54970 39516 54972
rect 39220 54918 39246 54970
rect 39246 54918 39276 54970
rect 39300 54918 39310 54970
rect 39310 54918 39356 54970
rect 39380 54918 39426 54970
rect 39426 54918 39436 54970
rect 39460 54918 39490 54970
rect 39490 54918 39516 54970
rect 39220 54916 39276 54918
rect 39300 54916 39356 54918
rect 39380 54916 39436 54918
rect 39460 54916 39516 54918
rect 39220 53882 39276 53884
rect 39300 53882 39356 53884
rect 39380 53882 39436 53884
rect 39460 53882 39516 53884
rect 39220 53830 39246 53882
rect 39246 53830 39276 53882
rect 39300 53830 39310 53882
rect 39310 53830 39356 53882
rect 39380 53830 39426 53882
rect 39426 53830 39436 53882
rect 39460 53830 39490 53882
rect 39490 53830 39516 53882
rect 39220 53828 39276 53830
rect 39300 53828 39356 53830
rect 39380 53828 39436 53830
rect 39460 53828 39516 53830
rect 39220 52794 39276 52796
rect 39300 52794 39356 52796
rect 39380 52794 39436 52796
rect 39460 52794 39516 52796
rect 39220 52742 39246 52794
rect 39246 52742 39276 52794
rect 39300 52742 39310 52794
rect 39310 52742 39356 52794
rect 39380 52742 39426 52794
rect 39426 52742 39436 52794
rect 39460 52742 39490 52794
rect 39490 52742 39516 52794
rect 39220 52740 39276 52742
rect 39300 52740 39356 52742
rect 39380 52740 39436 52742
rect 39460 52740 39516 52742
rect 39220 51706 39276 51708
rect 39300 51706 39356 51708
rect 39380 51706 39436 51708
rect 39460 51706 39516 51708
rect 39220 51654 39246 51706
rect 39246 51654 39276 51706
rect 39300 51654 39310 51706
rect 39310 51654 39356 51706
rect 39380 51654 39426 51706
rect 39426 51654 39436 51706
rect 39460 51654 39490 51706
rect 39490 51654 39516 51706
rect 39220 51652 39276 51654
rect 39300 51652 39356 51654
rect 39380 51652 39436 51654
rect 39460 51652 39516 51654
rect 39220 50618 39276 50620
rect 39300 50618 39356 50620
rect 39380 50618 39436 50620
rect 39460 50618 39516 50620
rect 39220 50566 39246 50618
rect 39246 50566 39276 50618
rect 39300 50566 39310 50618
rect 39310 50566 39356 50618
rect 39380 50566 39426 50618
rect 39426 50566 39436 50618
rect 39460 50566 39490 50618
rect 39490 50566 39516 50618
rect 39220 50564 39276 50566
rect 39300 50564 39356 50566
rect 39380 50564 39436 50566
rect 39460 50564 39516 50566
rect 39220 49530 39276 49532
rect 39300 49530 39356 49532
rect 39380 49530 39436 49532
rect 39460 49530 39516 49532
rect 39220 49478 39246 49530
rect 39246 49478 39276 49530
rect 39300 49478 39310 49530
rect 39310 49478 39356 49530
rect 39380 49478 39426 49530
rect 39426 49478 39436 49530
rect 39460 49478 39490 49530
rect 39490 49478 39516 49530
rect 39220 49476 39276 49478
rect 39300 49476 39356 49478
rect 39380 49476 39436 49478
rect 39460 49476 39516 49478
rect 39220 48442 39276 48444
rect 39300 48442 39356 48444
rect 39380 48442 39436 48444
rect 39460 48442 39516 48444
rect 39220 48390 39246 48442
rect 39246 48390 39276 48442
rect 39300 48390 39310 48442
rect 39310 48390 39356 48442
rect 39380 48390 39426 48442
rect 39426 48390 39436 48442
rect 39460 48390 39490 48442
rect 39490 48390 39516 48442
rect 39220 48388 39276 48390
rect 39300 48388 39356 48390
rect 39380 48388 39436 48390
rect 39460 48388 39516 48390
rect 39220 47354 39276 47356
rect 39300 47354 39356 47356
rect 39380 47354 39436 47356
rect 39460 47354 39516 47356
rect 39220 47302 39246 47354
rect 39246 47302 39276 47354
rect 39300 47302 39310 47354
rect 39310 47302 39356 47354
rect 39380 47302 39426 47354
rect 39426 47302 39436 47354
rect 39460 47302 39490 47354
rect 39490 47302 39516 47354
rect 39220 47300 39276 47302
rect 39300 47300 39356 47302
rect 39380 47300 39436 47302
rect 39460 47300 39516 47302
rect 39220 46266 39276 46268
rect 39300 46266 39356 46268
rect 39380 46266 39436 46268
rect 39460 46266 39516 46268
rect 39220 46214 39246 46266
rect 39246 46214 39276 46266
rect 39300 46214 39310 46266
rect 39310 46214 39356 46266
rect 39380 46214 39426 46266
rect 39426 46214 39436 46266
rect 39460 46214 39490 46266
rect 39490 46214 39516 46266
rect 39220 46212 39276 46214
rect 39300 46212 39356 46214
rect 39380 46212 39436 46214
rect 39460 46212 39516 46214
rect 39220 45178 39276 45180
rect 39300 45178 39356 45180
rect 39380 45178 39436 45180
rect 39460 45178 39516 45180
rect 39220 45126 39246 45178
rect 39246 45126 39276 45178
rect 39300 45126 39310 45178
rect 39310 45126 39356 45178
rect 39380 45126 39426 45178
rect 39426 45126 39436 45178
rect 39460 45126 39490 45178
rect 39490 45126 39516 45178
rect 39220 45124 39276 45126
rect 39300 45124 39356 45126
rect 39380 45124 39436 45126
rect 39460 45124 39516 45126
rect 39220 44090 39276 44092
rect 39300 44090 39356 44092
rect 39380 44090 39436 44092
rect 39460 44090 39516 44092
rect 39220 44038 39246 44090
rect 39246 44038 39276 44090
rect 39300 44038 39310 44090
rect 39310 44038 39356 44090
rect 39380 44038 39426 44090
rect 39426 44038 39436 44090
rect 39460 44038 39490 44090
rect 39490 44038 39516 44090
rect 39220 44036 39276 44038
rect 39300 44036 39356 44038
rect 39380 44036 39436 44038
rect 39460 44036 39516 44038
rect 39220 43002 39276 43004
rect 39300 43002 39356 43004
rect 39380 43002 39436 43004
rect 39460 43002 39516 43004
rect 39220 42950 39246 43002
rect 39246 42950 39276 43002
rect 39300 42950 39310 43002
rect 39310 42950 39356 43002
rect 39380 42950 39426 43002
rect 39426 42950 39436 43002
rect 39460 42950 39490 43002
rect 39490 42950 39516 43002
rect 39220 42948 39276 42950
rect 39300 42948 39356 42950
rect 39380 42948 39436 42950
rect 39460 42948 39516 42950
rect 39220 41914 39276 41916
rect 39300 41914 39356 41916
rect 39380 41914 39436 41916
rect 39460 41914 39516 41916
rect 39220 41862 39246 41914
rect 39246 41862 39276 41914
rect 39300 41862 39310 41914
rect 39310 41862 39356 41914
rect 39380 41862 39426 41914
rect 39426 41862 39436 41914
rect 39460 41862 39490 41914
rect 39490 41862 39516 41914
rect 39220 41860 39276 41862
rect 39300 41860 39356 41862
rect 39380 41860 39436 41862
rect 39460 41860 39516 41862
rect 39220 40826 39276 40828
rect 39300 40826 39356 40828
rect 39380 40826 39436 40828
rect 39460 40826 39516 40828
rect 39220 40774 39246 40826
rect 39246 40774 39276 40826
rect 39300 40774 39310 40826
rect 39310 40774 39356 40826
rect 39380 40774 39426 40826
rect 39426 40774 39436 40826
rect 39460 40774 39490 40826
rect 39490 40774 39516 40826
rect 39220 40772 39276 40774
rect 39300 40772 39356 40774
rect 39380 40772 39436 40774
rect 39460 40772 39516 40774
rect 39220 39738 39276 39740
rect 39300 39738 39356 39740
rect 39380 39738 39436 39740
rect 39460 39738 39516 39740
rect 39220 39686 39246 39738
rect 39246 39686 39276 39738
rect 39300 39686 39310 39738
rect 39310 39686 39356 39738
rect 39380 39686 39426 39738
rect 39426 39686 39436 39738
rect 39460 39686 39490 39738
rect 39490 39686 39516 39738
rect 39220 39684 39276 39686
rect 39300 39684 39356 39686
rect 39380 39684 39436 39686
rect 39460 39684 39516 39686
rect 39220 38650 39276 38652
rect 39300 38650 39356 38652
rect 39380 38650 39436 38652
rect 39460 38650 39516 38652
rect 39220 38598 39246 38650
rect 39246 38598 39276 38650
rect 39300 38598 39310 38650
rect 39310 38598 39356 38650
rect 39380 38598 39426 38650
rect 39426 38598 39436 38650
rect 39460 38598 39490 38650
rect 39490 38598 39516 38650
rect 39220 38596 39276 38598
rect 39300 38596 39356 38598
rect 39380 38596 39436 38598
rect 39460 38596 39516 38598
rect 39220 37562 39276 37564
rect 39300 37562 39356 37564
rect 39380 37562 39436 37564
rect 39460 37562 39516 37564
rect 39220 37510 39246 37562
rect 39246 37510 39276 37562
rect 39300 37510 39310 37562
rect 39310 37510 39356 37562
rect 39380 37510 39426 37562
rect 39426 37510 39436 37562
rect 39460 37510 39490 37562
rect 39490 37510 39516 37562
rect 39220 37508 39276 37510
rect 39300 37508 39356 37510
rect 39380 37508 39436 37510
rect 39460 37508 39516 37510
rect 39220 36474 39276 36476
rect 39300 36474 39356 36476
rect 39380 36474 39436 36476
rect 39460 36474 39516 36476
rect 39220 36422 39246 36474
rect 39246 36422 39276 36474
rect 39300 36422 39310 36474
rect 39310 36422 39356 36474
rect 39380 36422 39426 36474
rect 39426 36422 39436 36474
rect 39460 36422 39490 36474
rect 39490 36422 39516 36474
rect 39220 36420 39276 36422
rect 39300 36420 39356 36422
rect 39380 36420 39436 36422
rect 39460 36420 39516 36422
rect 39220 35386 39276 35388
rect 39300 35386 39356 35388
rect 39380 35386 39436 35388
rect 39460 35386 39516 35388
rect 39220 35334 39246 35386
rect 39246 35334 39276 35386
rect 39300 35334 39310 35386
rect 39310 35334 39356 35386
rect 39380 35334 39426 35386
rect 39426 35334 39436 35386
rect 39460 35334 39490 35386
rect 39490 35334 39516 35386
rect 39220 35332 39276 35334
rect 39300 35332 39356 35334
rect 39380 35332 39436 35334
rect 39460 35332 39516 35334
rect 39220 34298 39276 34300
rect 39300 34298 39356 34300
rect 39380 34298 39436 34300
rect 39460 34298 39516 34300
rect 39220 34246 39246 34298
rect 39246 34246 39276 34298
rect 39300 34246 39310 34298
rect 39310 34246 39356 34298
rect 39380 34246 39426 34298
rect 39426 34246 39436 34298
rect 39460 34246 39490 34298
rect 39490 34246 39516 34298
rect 39220 34244 39276 34246
rect 39300 34244 39356 34246
rect 39380 34244 39436 34246
rect 39460 34244 39516 34246
rect 39220 33210 39276 33212
rect 39300 33210 39356 33212
rect 39380 33210 39436 33212
rect 39460 33210 39516 33212
rect 39220 33158 39246 33210
rect 39246 33158 39276 33210
rect 39300 33158 39310 33210
rect 39310 33158 39356 33210
rect 39380 33158 39426 33210
rect 39426 33158 39436 33210
rect 39460 33158 39490 33210
rect 39490 33158 39516 33210
rect 39220 33156 39276 33158
rect 39300 33156 39356 33158
rect 39380 33156 39436 33158
rect 39460 33156 39516 33158
rect 39220 32122 39276 32124
rect 39300 32122 39356 32124
rect 39380 32122 39436 32124
rect 39460 32122 39516 32124
rect 39220 32070 39246 32122
rect 39246 32070 39276 32122
rect 39300 32070 39310 32122
rect 39310 32070 39356 32122
rect 39380 32070 39426 32122
rect 39426 32070 39436 32122
rect 39460 32070 39490 32122
rect 39490 32070 39516 32122
rect 39220 32068 39276 32070
rect 39300 32068 39356 32070
rect 39380 32068 39436 32070
rect 39460 32068 39516 32070
rect 39220 31034 39276 31036
rect 39300 31034 39356 31036
rect 39380 31034 39436 31036
rect 39460 31034 39516 31036
rect 39220 30982 39246 31034
rect 39246 30982 39276 31034
rect 39300 30982 39310 31034
rect 39310 30982 39356 31034
rect 39380 30982 39426 31034
rect 39426 30982 39436 31034
rect 39460 30982 39490 31034
rect 39490 30982 39516 31034
rect 39220 30980 39276 30982
rect 39300 30980 39356 30982
rect 39380 30980 39436 30982
rect 39460 30980 39516 30982
rect 37922 6316 37978 6352
rect 37922 6296 37924 6316
rect 37924 6296 37976 6316
rect 37976 6296 37978 6316
rect 38290 12008 38346 12064
rect 38750 7384 38806 7440
rect 38658 6024 38714 6080
rect 38566 5888 38622 5944
rect 38658 4120 38714 4176
rect 39220 29946 39276 29948
rect 39300 29946 39356 29948
rect 39380 29946 39436 29948
rect 39460 29946 39516 29948
rect 39220 29894 39246 29946
rect 39246 29894 39276 29946
rect 39300 29894 39310 29946
rect 39310 29894 39356 29946
rect 39380 29894 39426 29946
rect 39426 29894 39436 29946
rect 39460 29894 39490 29946
rect 39490 29894 39516 29946
rect 39220 29892 39276 29894
rect 39300 29892 39356 29894
rect 39380 29892 39436 29894
rect 39460 29892 39516 29894
rect 39220 28858 39276 28860
rect 39300 28858 39356 28860
rect 39380 28858 39436 28860
rect 39460 28858 39516 28860
rect 39220 28806 39246 28858
rect 39246 28806 39276 28858
rect 39300 28806 39310 28858
rect 39310 28806 39356 28858
rect 39380 28806 39426 28858
rect 39426 28806 39436 28858
rect 39460 28806 39490 28858
rect 39490 28806 39516 28858
rect 39220 28804 39276 28806
rect 39300 28804 39356 28806
rect 39380 28804 39436 28806
rect 39460 28804 39516 28806
rect 39220 27770 39276 27772
rect 39300 27770 39356 27772
rect 39380 27770 39436 27772
rect 39460 27770 39516 27772
rect 39220 27718 39246 27770
rect 39246 27718 39276 27770
rect 39300 27718 39310 27770
rect 39310 27718 39356 27770
rect 39380 27718 39426 27770
rect 39426 27718 39436 27770
rect 39460 27718 39490 27770
rect 39490 27718 39516 27770
rect 39220 27716 39276 27718
rect 39300 27716 39356 27718
rect 39380 27716 39436 27718
rect 39460 27716 39516 27718
rect 39220 26682 39276 26684
rect 39300 26682 39356 26684
rect 39380 26682 39436 26684
rect 39460 26682 39516 26684
rect 39220 26630 39246 26682
rect 39246 26630 39276 26682
rect 39300 26630 39310 26682
rect 39310 26630 39356 26682
rect 39380 26630 39426 26682
rect 39426 26630 39436 26682
rect 39460 26630 39490 26682
rect 39490 26630 39516 26682
rect 39220 26628 39276 26630
rect 39300 26628 39356 26630
rect 39380 26628 39436 26630
rect 39460 26628 39516 26630
rect 39220 25594 39276 25596
rect 39300 25594 39356 25596
rect 39380 25594 39436 25596
rect 39460 25594 39516 25596
rect 39220 25542 39246 25594
rect 39246 25542 39276 25594
rect 39300 25542 39310 25594
rect 39310 25542 39356 25594
rect 39380 25542 39426 25594
rect 39426 25542 39436 25594
rect 39460 25542 39490 25594
rect 39490 25542 39516 25594
rect 39220 25540 39276 25542
rect 39300 25540 39356 25542
rect 39380 25540 39436 25542
rect 39460 25540 39516 25542
rect 39220 24506 39276 24508
rect 39300 24506 39356 24508
rect 39380 24506 39436 24508
rect 39460 24506 39516 24508
rect 39220 24454 39246 24506
rect 39246 24454 39276 24506
rect 39300 24454 39310 24506
rect 39310 24454 39356 24506
rect 39380 24454 39426 24506
rect 39426 24454 39436 24506
rect 39460 24454 39490 24506
rect 39490 24454 39516 24506
rect 39220 24452 39276 24454
rect 39300 24452 39356 24454
rect 39380 24452 39436 24454
rect 39460 24452 39516 24454
rect 39220 23418 39276 23420
rect 39300 23418 39356 23420
rect 39380 23418 39436 23420
rect 39460 23418 39516 23420
rect 39220 23366 39246 23418
rect 39246 23366 39276 23418
rect 39300 23366 39310 23418
rect 39310 23366 39356 23418
rect 39380 23366 39426 23418
rect 39426 23366 39436 23418
rect 39460 23366 39490 23418
rect 39490 23366 39516 23418
rect 39220 23364 39276 23366
rect 39300 23364 39356 23366
rect 39380 23364 39436 23366
rect 39460 23364 39516 23366
rect 39220 22330 39276 22332
rect 39300 22330 39356 22332
rect 39380 22330 39436 22332
rect 39460 22330 39516 22332
rect 39220 22278 39246 22330
rect 39246 22278 39276 22330
rect 39300 22278 39310 22330
rect 39310 22278 39356 22330
rect 39380 22278 39426 22330
rect 39426 22278 39436 22330
rect 39460 22278 39490 22330
rect 39490 22278 39516 22330
rect 39220 22276 39276 22278
rect 39300 22276 39356 22278
rect 39380 22276 39436 22278
rect 39460 22276 39516 22278
rect 39220 21242 39276 21244
rect 39300 21242 39356 21244
rect 39380 21242 39436 21244
rect 39460 21242 39516 21244
rect 39220 21190 39246 21242
rect 39246 21190 39276 21242
rect 39300 21190 39310 21242
rect 39310 21190 39356 21242
rect 39380 21190 39426 21242
rect 39426 21190 39436 21242
rect 39460 21190 39490 21242
rect 39490 21190 39516 21242
rect 39220 21188 39276 21190
rect 39300 21188 39356 21190
rect 39380 21188 39436 21190
rect 39460 21188 39516 21190
rect 39220 20154 39276 20156
rect 39300 20154 39356 20156
rect 39380 20154 39436 20156
rect 39460 20154 39516 20156
rect 39220 20102 39246 20154
rect 39246 20102 39276 20154
rect 39300 20102 39310 20154
rect 39310 20102 39356 20154
rect 39380 20102 39426 20154
rect 39426 20102 39436 20154
rect 39460 20102 39490 20154
rect 39490 20102 39516 20154
rect 39220 20100 39276 20102
rect 39300 20100 39356 20102
rect 39380 20100 39436 20102
rect 39460 20100 39516 20102
rect 39220 19066 39276 19068
rect 39300 19066 39356 19068
rect 39380 19066 39436 19068
rect 39460 19066 39516 19068
rect 39220 19014 39246 19066
rect 39246 19014 39276 19066
rect 39300 19014 39310 19066
rect 39310 19014 39356 19066
rect 39380 19014 39426 19066
rect 39426 19014 39436 19066
rect 39460 19014 39490 19066
rect 39490 19014 39516 19066
rect 39220 19012 39276 19014
rect 39300 19012 39356 19014
rect 39380 19012 39436 19014
rect 39460 19012 39516 19014
rect 39220 17978 39276 17980
rect 39300 17978 39356 17980
rect 39380 17978 39436 17980
rect 39460 17978 39516 17980
rect 39220 17926 39246 17978
rect 39246 17926 39276 17978
rect 39300 17926 39310 17978
rect 39310 17926 39356 17978
rect 39380 17926 39426 17978
rect 39426 17926 39436 17978
rect 39460 17926 39490 17978
rect 39490 17926 39516 17978
rect 39220 17924 39276 17926
rect 39300 17924 39356 17926
rect 39380 17924 39436 17926
rect 39460 17924 39516 17926
rect 39220 16890 39276 16892
rect 39300 16890 39356 16892
rect 39380 16890 39436 16892
rect 39460 16890 39516 16892
rect 39220 16838 39246 16890
rect 39246 16838 39276 16890
rect 39300 16838 39310 16890
rect 39310 16838 39356 16890
rect 39380 16838 39426 16890
rect 39426 16838 39436 16890
rect 39460 16838 39490 16890
rect 39490 16838 39516 16890
rect 39220 16836 39276 16838
rect 39300 16836 39356 16838
rect 39380 16836 39436 16838
rect 39460 16836 39516 16838
rect 39220 15802 39276 15804
rect 39300 15802 39356 15804
rect 39380 15802 39436 15804
rect 39460 15802 39516 15804
rect 39220 15750 39246 15802
rect 39246 15750 39276 15802
rect 39300 15750 39310 15802
rect 39310 15750 39356 15802
rect 39380 15750 39426 15802
rect 39426 15750 39436 15802
rect 39460 15750 39490 15802
rect 39490 15750 39516 15802
rect 39220 15748 39276 15750
rect 39300 15748 39356 15750
rect 39380 15748 39436 15750
rect 39460 15748 39516 15750
rect 39220 14714 39276 14716
rect 39300 14714 39356 14716
rect 39380 14714 39436 14716
rect 39460 14714 39516 14716
rect 39220 14662 39246 14714
rect 39246 14662 39276 14714
rect 39300 14662 39310 14714
rect 39310 14662 39356 14714
rect 39380 14662 39426 14714
rect 39426 14662 39436 14714
rect 39460 14662 39490 14714
rect 39490 14662 39516 14714
rect 39220 14660 39276 14662
rect 39300 14660 39356 14662
rect 39380 14660 39436 14662
rect 39460 14660 39516 14662
rect 39220 13626 39276 13628
rect 39300 13626 39356 13628
rect 39380 13626 39436 13628
rect 39460 13626 39516 13628
rect 39220 13574 39246 13626
rect 39246 13574 39276 13626
rect 39300 13574 39310 13626
rect 39310 13574 39356 13626
rect 39380 13574 39426 13626
rect 39426 13574 39436 13626
rect 39460 13574 39490 13626
rect 39490 13574 39516 13626
rect 39220 13572 39276 13574
rect 39300 13572 39356 13574
rect 39380 13572 39436 13574
rect 39460 13572 39516 13574
rect 39210 13132 39212 13152
rect 39212 13132 39264 13152
rect 39264 13132 39266 13152
rect 39210 13096 39266 13132
rect 39220 12538 39276 12540
rect 39300 12538 39356 12540
rect 39380 12538 39436 12540
rect 39460 12538 39516 12540
rect 39220 12486 39246 12538
rect 39246 12486 39276 12538
rect 39300 12486 39310 12538
rect 39310 12486 39356 12538
rect 39380 12486 39426 12538
rect 39426 12486 39436 12538
rect 39460 12486 39490 12538
rect 39490 12486 39516 12538
rect 39220 12484 39276 12486
rect 39300 12484 39356 12486
rect 39380 12484 39436 12486
rect 39460 12484 39516 12486
rect 38658 3576 38714 3632
rect 38658 3304 38714 3360
rect 38750 2488 38806 2544
rect 38658 1944 38714 2000
rect 39220 11450 39276 11452
rect 39300 11450 39356 11452
rect 39380 11450 39436 11452
rect 39460 11450 39516 11452
rect 39220 11398 39246 11450
rect 39246 11398 39276 11450
rect 39300 11398 39310 11450
rect 39310 11398 39356 11450
rect 39380 11398 39426 11450
rect 39426 11398 39436 11450
rect 39460 11398 39490 11450
rect 39490 11398 39516 11450
rect 39220 11396 39276 11398
rect 39300 11396 39356 11398
rect 39380 11396 39436 11398
rect 39460 11396 39516 11398
rect 39220 10362 39276 10364
rect 39300 10362 39356 10364
rect 39380 10362 39436 10364
rect 39460 10362 39516 10364
rect 39220 10310 39246 10362
rect 39246 10310 39276 10362
rect 39300 10310 39310 10362
rect 39310 10310 39356 10362
rect 39380 10310 39426 10362
rect 39426 10310 39436 10362
rect 39460 10310 39490 10362
rect 39490 10310 39516 10362
rect 39220 10308 39276 10310
rect 39300 10308 39356 10310
rect 39380 10308 39436 10310
rect 39460 10308 39516 10310
rect 39486 9424 39542 9480
rect 39220 9274 39276 9276
rect 39300 9274 39356 9276
rect 39380 9274 39436 9276
rect 39460 9274 39516 9276
rect 39220 9222 39246 9274
rect 39246 9222 39276 9274
rect 39300 9222 39310 9274
rect 39310 9222 39356 9274
rect 39380 9222 39426 9274
rect 39426 9222 39436 9274
rect 39460 9222 39490 9274
rect 39490 9222 39516 9274
rect 39220 9220 39276 9222
rect 39300 9220 39356 9222
rect 39380 9220 39436 9222
rect 39460 9220 39516 9222
rect 39026 9036 39082 9072
rect 39026 9016 39028 9036
rect 39028 9016 39080 9036
rect 39080 9016 39082 9036
rect 39394 8472 39450 8528
rect 39220 8186 39276 8188
rect 39300 8186 39356 8188
rect 39380 8186 39436 8188
rect 39460 8186 39516 8188
rect 39220 8134 39246 8186
rect 39246 8134 39276 8186
rect 39300 8134 39310 8186
rect 39310 8134 39356 8186
rect 39380 8134 39426 8186
rect 39426 8134 39436 8186
rect 39460 8134 39490 8186
rect 39490 8134 39516 8186
rect 39220 8132 39276 8134
rect 39300 8132 39356 8134
rect 39380 8132 39436 8134
rect 39460 8132 39516 8134
rect 39220 7098 39276 7100
rect 39300 7098 39356 7100
rect 39380 7098 39436 7100
rect 39460 7098 39516 7100
rect 39220 7046 39246 7098
rect 39246 7046 39276 7098
rect 39300 7046 39310 7098
rect 39310 7046 39356 7098
rect 39380 7046 39426 7098
rect 39426 7046 39436 7098
rect 39460 7046 39490 7098
rect 39490 7046 39516 7098
rect 39220 7044 39276 7046
rect 39300 7044 39356 7046
rect 39380 7044 39436 7046
rect 39460 7044 39516 7046
rect 39220 6010 39276 6012
rect 39300 6010 39356 6012
rect 39380 6010 39436 6012
rect 39460 6010 39516 6012
rect 39220 5958 39246 6010
rect 39246 5958 39276 6010
rect 39300 5958 39310 6010
rect 39310 5958 39356 6010
rect 39380 5958 39426 6010
rect 39426 5958 39436 6010
rect 39460 5958 39490 6010
rect 39490 5958 39516 6010
rect 39220 5956 39276 5958
rect 39300 5956 39356 5958
rect 39380 5956 39436 5958
rect 39460 5956 39516 5958
rect 39210 5636 39266 5672
rect 39210 5616 39212 5636
rect 39212 5616 39264 5636
rect 39264 5616 39266 5636
rect 39220 4922 39276 4924
rect 39300 4922 39356 4924
rect 39380 4922 39436 4924
rect 39460 4922 39516 4924
rect 39220 4870 39246 4922
rect 39246 4870 39276 4922
rect 39300 4870 39310 4922
rect 39310 4870 39356 4922
rect 39380 4870 39426 4922
rect 39426 4870 39436 4922
rect 39460 4870 39490 4922
rect 39490 4870 39516 4922
rect 39220 4868 39276 4870
rect 39300 4868 39356 4870
rect 39380 4868 39436 4870
rect 39460 4868 39516 4870
rect 39026 4664 39082 4720
rect 39762 12416 39818 12472
rect 39762 12180 39764 12200
rect 39764 12180 39816 12200
rect 39816 12180 39818 12200
rect 39762 12144 39818 12180
rect 39946 12980 40002 13016
rect 39946 12960 39948 12980
rect 39948 12960 40000 12980
rect 40000 12960 40002 12980
rect 39670 11328 39726 11384
rect 39670 11056 39726 11112
rect 39670 6976 39726 7032
rect 39854 8880 39910 8936
rect 39854 6568 39910 6624
rect 39026 3712 39082 3768
rect 39670 4528 39726 4584
rect 39394 4120 39450 4176
rect 39220 3834 39276 3836
rect 39300 3834 39356 3836
rect 39380 3834 39436 3836
rect 39460 3834 39516 3836
rect 39220 3782 39246 3834
rect 39246 3782 39276 3834
rect 39300 3782 39310 3834
rect 39310 3782 39356 3834
rect 39380 3782 39426 3834
rect 39426 3782 39436 3834
rect 39460 3782 39490 3834
rect 39490 3782 39516 3834
rect 39220 3780 39276 3782
rect 39300 3780 39356 3782
rect 39380 3780 39436 3782
rect 39460 3780 39516 3782
rect 39854 4684 39910 4720
rect 39854 4664 39856 4684
rect 39856 4664 39908 4684
rect 39908 4664 39910 4684
rect 39210 3304 39266 3360
rect 39486 3304 39542 3360
rect 39220 2746 39276 2748
rect 39300 2746 39356 2748
rect 39380 2746 39436 2748
rect 39460 2746 39516 2748
rect 39220 2694 39246 2746
rect 39246 2694 39276 2746
rect 39300 2694 39310 2746
rect 39310 2694 39356 2746
rect 39380 2694 39426 2746
rect 39426 2694 39436 2746
rect 39460 2694 39490 2746
rect 39490 2694 39516 2746
rect 39220 2692 39276 2694
rect 39300 2692 39356 2694
rect 39380 2692 39436 2694
rect 39460 2692 39516 2694
rect 39210 2216 39266 2272
rect 39762 3440 39818 3496
rect 40130 10512 40186 10568
rect 40038 5480 40094 5536
rect 40498 9152 40554 9208
rect 40406 6568 40462 6624
rect 40130 2796 40132 2816
rect 40132 2796 40184 2816
rect 40184 2796 40186 2816
rect 40130 2760 40186 2796
rect 39486 1264 39542 1320
rect 40498 6024 40554 6080
rect 40498 3052 40554 3088
rect 40498 3032 40500 3052
rect 40500 3032 40552 3052
rect 40552 3032 40554 3052
rect 40866 12588 40868 12608
rect 40868 12588 40920 12608
rect 40920 12588 40922 12608
rect 40866 12552 40922 12588
rect 40866 9968 40922 10024
rect 40682 3032 40738 3088
rect 44220 66394 44276 66396
rect 44300 66394 44356 66396
rect 44380 66394 44436 66396
rect 44460 66394 44516 66396
rect 44220 66342 44246 66394
rect 44246 66342 44276 66394
rect 44300 66342 44310 66394
rect 44310 66342 44356 66394
rect 44380 66342 44426 66394
rect 44426 66342 44436 66394
rect 44460 66342 44490 66394
rect 44490 66342 44516 66394
rect 44220 66340 44276 66342
rect 44300 66340 44356 66342
rect 44380 66340 44436 66342
rect 44460 66340 44516 66342
rect 49220 65850 49276 65852
rect 49300 65850 49356 65852
rect 49380 65850 49436 65852
rect 49460 65850 49516 65852
rect 49220 65798 49246 65850
rect 49246 65798 49276 65850
rect 49300 65798 49310 65850
rect 49310 65798 49356 65850
rect 49380 65798 49426 65850
rect 49426 65798 49436 65850
rect 49460 65798 49490 65850
rect 49490 65798 49516 65850
rect 49220 65796 49276 65798
rect 49300 65796 49356 65798
rect 49380 65796 49436 65798
rect 49460 65796 49516 65798
rect 44220 65306 44276 65308
rect 44300 65306 44356 65308
rect 44380 65306 44436 65308
rect 44460 65306 44516 65308
rect 44220 65254 44246 65306
rect 44246 65254 44276 65306
rect 44300 65254 44310 65306
rect 44310 65254 44356 65306
rect 44380 65254 44426 65306
rect 44426 65254 44436 65306
rect 44460 65254 44490 65306
rect 44490 65254 44516 65306
rect 44220 65252 44276 65254
rect 44300 65252 44356 65254
rect 44380 65252 44436 65254
rect 44460 65252 44516 65254
rect 49220 64762 49276 64764
rect 49300 64762 49356 64764
rect 49380 64762 49436 64764
rect 49460 64762 49516 64764
rect 49220 64710 49246 64762
rect 49246 64710 49276 64762
rect 49300 64710 49310 64762
rect 49310 64710 49356 64762
rect 49380 64710 49426 64762
rect 49426 64710 49436 64762
rect 49460 64710 49490 64762
rect 49490 64710 49516 64762
rect 49220 64708 49276 64710
rect 49300 64708 49356 64710
rect 49380 64708 49436 64710
rect 49460 64708 49516 64710
rect 44220 64218 44276 64220
rect 44300 64218 44356 64220
rect 44380 64218 44436 64220
rect 44460 64218 44516 64220
rect 44220 64166 44246 64218
rect 44246 64166 44276 64218
rect 44300 64166 44310 64218
rect 44310 64166 44356 64218
rect 44380 64166 44426 64218
rect 44426 64166 44436 64218
rect 44460 64166 44490 64218
rect 44490 64166 44516 64218
rect 44220 64164 44276 64166
rect 44300 64164 44356 64166
rect 44380 64164 44436 64166
rect 44460 64164 44516 64166
rect 49220 63674 49276 63676
rect 49300 63674 49356 63676
rect 49380 63674 49436 63676
rect 49460 63674 49516 63676
rect 49220 63622 49246 63674
rect 49246 63622 49276 63674
rect 49300 63622 49310 63674
rect 49310 63622 49356 63674
rect 49380 63622 49426 63674
rect 49426 63622 49436 63674
rect 49460 63622 49490 63674
rect 49490 63622 49516 63674
rect 49220 63620 49276 63622
rect 49300 63620 49356 63622
rect 49380 63620 49436 63622
rect 49460 63620 49516 63622
rect 44220 63130 44276 63132
rect 44300 63130 44356 63132
rect 44380 63130 44436 63132
rect 44460 63130 44516 63132
rect 44220 63078 44246 63130
rect 44246 63078 44276 63130
rect 44300 63078 44310 63130
rect 44310 63078 44356 63130
rect 44380 63078 44426 63130
rect 44426 63078 44436 63130
rect 44460 63078 44490 63130
rect 44490 63078 44516 63130
rect 44220 63076 44276 63078
rect 44300 63076 44356 63078
rect 44380 63076 44436 63078
rect 44460 63076 44516 63078
rect 44220 62042 44276 62044
rect 44300 62042 44356 62044
rect 44380 62042 44436 62044
rect 44460 62042 44516 62044
rect 44220 61990 44246 62042
rect 44246 61990 44276 62042
rect 44300 61990 44310 62042
rect 44310 61990 44356 62042
rect 44380 61990 44426 62042
rect 44426 61990 44436 62042
rect 44460 61990 44490 62042
rect 44490 61990 44516 62042
rect 44220 61988 44276 61990
rect 44300 61988 44356 61990
rect 44380 61988 44436 61990
rect 44460 61988 44516 61990
rect 44220 60954 44276 60956
rect 44300 60954 44356 60956
rect 44380 60954 44436 60956
rect 44460 60954 44516 60956
rect 44220 60902 44246 60954
rect 44246 60902 44276 60954
rect 44300 60902 44310 60954
rect 44310 60902 44356 60954
rect 44380 60902 44426 60954
rect 44426 60902 44436 60954
rect 44460 60902 44490 60954
rect 44490 60902 44516 60954
rect 44220 60900 44276 60902
rect 44300 60900 44356 60902
rect 44380 60900 44436 60902
rect 44460 60900 44516 60902
rect 44220 59866 44276 59868
rect 44300 59866 44356 59868
rect 44380 59866 44436 59868
rect 44460 59866 44516 59868
rect 44220 59814 44246 59866
rect 44246 59814 44276 59866
rect 44300 59814 44310 59866
rect 44310 59814 44356 59866
rect 44380 59814 44426 59866
rect 44426 59814 44436 59866
rect 44460 59814 44490 59866
rect 44490 59814 44516 59866
rect 44220 59812 44276 59814
rect 44300 59812 44356 59814
rect 44380 59812 44436 59814
rect 44460 59812 44516 59814
rect 44220 58778 44276 58780
rect 44300 58778 44356 58780
rect 44380 58778 44436 58780
rect 44460 58778 44516 58780
rect 44220 58726 44246 58778
rect 44246 58726 44276 58778
rect 44300 58726 44310 58778
rect 44310 58726 44356 58778
rect 44380 58726 44426 58778
rect 44426 58726 44436 58778
rect 44460 58726 44490 58778
rect 44490 58726 44516 58778
rect 44220 58724 44276 58726
rect 44300 58724 44356 58726
rect 44380 58724 44436 58726
rect 44460 58724 44516 58726
rect 41510 14456 41566 14512
rect 41326 8200 41382 8256
rect 41970 10784 42026 10840
rect 41142 6060 41144 6080
rect 41144 6060 41196 6080
rect 41196 6060 41198 6080
rect 41142 6024 41198 6060
rect 41142 4528 41198 4584
rect 41050 2896 41106 2952
rect 41694 6432 41750 6488
rect 41418 3032 41474 3088
rect 41786 5208 41842 5264
rect 41694 3304 41750 3360
rect 42338 11056 42394 11112
rect 42338 8880 42394 8936
rect 42338 5888 42394 5944
rect 42706 11076 42762 11112
rect 42706 11056 42708 11076
rect 42708 11056 42760 11076
rect 42760 11056 42762 11076
rect 42890 9016 42946 9072
rect 42890 6860 42946 6896
rect 42890 6840 42892 6860
rect 42892 6840 42944 6860
rect 42944 6840 42946 6860
rect 42614 4684 42670 4720
rect 42614 4664 42616 4684
rect 42616 4664 42668 4684
rect 42668 4664 42670 4684
rect 42062 3304 42118 3360
rect 41602 2488 41658 2544
rect 41970 2760 42026 2816
rect 42430 2624 42486 2680
rect 42338 2352 42394 2408
rect 42706 3032 42762 3088
rect 42890 3168 42946 3224
rect 43074 6024 43130 6080
rect 44220 57690 44276 57692
rect 44300 57690 44356 57692
rect 44380 57690 44436 57692
rect 44460 57690 44516 57692
rect 44220 57638 44246 57690
rect 44246 57638 44276 57690
rect 44300 57638 44310 57690
rect 44310 57638 44356 57690
rect 44380 57638 44426 57690
rect 44426 57638 44436 57690
rect 44460 57638 44490 57690
rect 44490 57638 44516 57690
rect 44220 57636 44276 57638
rect 44300 57636 44356 57638
rect 44380 57636 44436 57638
rect 44460 57636 44516 57638
rect 44220 56602 44276 56604
rect 44300 56602 44356 56604
rect 44380 56602 44436 56604
rect 44460 56602 44516 56604
rect 44220 56550 44246 56602
rect 44246 56550 44276 56602
rect 44300 56550 44310 56602
rect 44310 56550 44356 56602
rect 44380 56550 44426 56602
rect 44426 56550 44436 56602
rect 44460 56550 44490 56602
rect 44490 56550 44516 56602
rect 44220 56548 44276 56550
rect 44300 56548 44356 56550
rect 44380 56548 44436 56550
rect 44460 56548 44516 56550
rect 44220 55514 44276 55516
rect 44300 55514 44356 55516
rect 44380 55514 44436 55516
rect 44460 55514 44516 55516
rect 44220 55462 44246 55514
rect 44246 55462 44276 55514
rect 44300 55462 44310 55514
rect 44310 55462 44356 55514
rect 44380 55462 44426 55514
rect 44426 55462 44436 55514
rect 44460 55462 44490 55514
rect 44490 55462 44516 55514
rect 44220 55460 44276 55462
rect 44300 55460 44356 55462
rect 44380 55460 44436 55462
rect 44460 55460 44516 55462
rect 44220 54426 44276 54428
rect 44300 54426 44356 54428
rect 44380 54426 44436 54428
rect 44460 54426 44516 54428
rect 44220 54374 44246 54426
rect 44246 54374 44276 54426
rect 44300 54374 44310 54426
rect 44310 54374 44356 54426
rect 44380 54374 44426 54426
rect 44426 54374 44436 54426
rect 44460 54374 44490 54426
rect 44490 54374 44516 54426
rect 44220 54372 44276 54374
rect 44300 54372 44356 54374
rect 44380 54372 44436 54374
rect 44460 54372 44516 54374
rect 44220 53338 44276 53340
rect 44300 53338 44356 53340
rect 44380 53338 44436 53340
rect 44460 53338 44516 53340
rect 44220 53286 44246 53338
rect 44246 53286 44276 53338
rect 44300 53286 44310 53338
rect 44310 53286 44356 53338
rect 44380 53286 44426 53338
rect 44426 53286 44436 53338
rect 44460 53286 44490 53338
rect 44490 53286 44516 53338
rect 44220 53284 44276 53286
rect 44300 53284 44356 53286
rect 44380 53284 44436 53286
rect 44460 53284 44516 53286
rect 44220 52250 44276 52252
rect 44300 52250 44356 52252
rect 44380 52250 44436 52252
rect 44460 52250 44516 52252
rect 44220 52198 44246 52250
rect 44246 52198 44276 52250
rect 44300 52198 44310 52250
rect 44310 52198 44356 52250
rect 44380 52198 44426 52250
rect 44426 52198 44436 52250
rect 44460 52198 44490 52250
rect 44490 52198 44516 52250
rect 44220 52196 44276 52198
rect 44300 52196 44356 52198
rect 44380 52196 44436 52198
rect 44460 52196 44516 52198
rect 44220 51162 44276 51164
rect 44300 51162 44356 51164
rect 44380 51162 44436 51164
rect 44460 51162 44516 51164
rect 44220 51110 44246 51162
rect 44246 51110 44276 51162
rect 44300 51110 44310 51162
rect 44310 51110 44356 51162
rect 44380 51110 44426 51162
rect 44426 51110 44436 51162
rect 44460 51110 44490 51162
rect 44490 51110 44516 51162
rect 44220 51108 44276 51110
rect 44300 51108 44356 51110
rect 44380 51108 44436 51110
rect 44460 51108 44516 51110
rect 44220 50074 44276 50076
rect 44300 50074 44356 50076
rect 44380 50074 44436 50076
rect 44460 50074 44516 50076
rect 44220 50022 44246 50074
rect 44246 50022 44276 50074
rect 44300 50022 44310 50074
rect 44310 50022 44356 50074
rect 44380 50022 44426 50074
rect 44426 50022 44436 50074
rect 44460 50022 44490 50074
rect 44490 50022 44516 50074
rect 44220 50020 44276 50022
rect 44300 50020 44356 50022
rect 44380 50020 44436 50022
rect 44460 50020 44516 50022
rect 44220 48986 44276 48988
rect 44300 48986 44356 48988
rect 44380 48986 44436 48988
rect 44460 48986 44516 48988
rect 44220 48934 44246 48986
rect 44246 48934 44276 48986
rect 44300 48934 44310 48986
rect 44310 48934 44356 48986
rect 44380 48934 44426 48986
rect 44426 48934 44436 48986
rect 44460 48934 44490 48986
rect 44490 48934 44516 48986
rect 44220 48932 44276 48934
rect 44300 48932 44356 48934
rect 44380 48932 44436 48934
rect 44460 48932 44516 48934
rect 44220 47898 44276 47900
rect 44300 47898 44356 47900
rect 44380 47898 44436 47900
rect 44460 47898 44516 47900
rect 44220 47846 44246 47898
rect 44246 47846 44276 47898
rect 44300 47846 44310 47898
rect 44310 47846 44356 47898
rect 44380 47846 44426 47898
rect 44426 47846 44436 47898
rect 44460 47846 44490 47898
rect 44490 47846 44516 47898
rect 44220 47844 44276 47846
rect 44300 47844 44356 47846
rect 44380 47844 44436 47846
rect 44460 47844 44516 47846
rect 44220 46810 44276 46812
rect 44300 46810 44356 46812
rect 44380 46810 44436 46812
rect 44460 46810 44516 46812
rect 44220 46758 44246 46810
rect 44246 46758 44276 46810
rect 44300 46758 44310 46810
rect 44310 46758 44356 46810
rect 44380 46758 44426 46810
rect 44426 46758 44436 46810
rect 44460 46758 44490 46810
rect 44490 46758 44516 46810
rect 44220 46756 44276 46758
rect 44300 46756 44356 46758
rect 44380 46756 44436 46758
rect 44460 46756 44516 46758
rect 44220 45722 44276 45724
rect 44300 45722 44356 45724
rect 44380 45722 44436 45724
rect 44460 45722 44516 45724
rect 44220 45670 44246 45722
rect 44246 45670 44276 45722
rect 44300 45670 44310 45722
rect 44310 45670 44356 45722
rect 44380 45670 44426 45722
rect 44426 45670 44436 45722
rect 44460 45670 44490 45722
rect 44490 45670 44516 45722
rect 44220 45668 44276 45670
rect 44300 45668 44356 45670
rect 44380 45668 44436 45670
rect 44460 45668 44516 45670
rect 44220 44634 44276 44636
rect 44300 44634 44356 44636
rect 44380 44634 44436 44636
rect 44460 44634 44516 44636
rect 44220 44582 44246 44634
rect 44246 44582 44276 44634
rect 44300 44582 44310 44634
rect 44310 44582 44356 44634
rect 44380 44582 44426 44634
rect 44426 44582 44436 44634
rect 44460 44582 44490 44634
rect 44490 44582 44516 44634
rect 44220 44580 44276 44582
rect 44300 44580 44356 44582
rect 44380 44580 44436 44582
rect 44460 44580 44516 44582
rect 44220 43546 44276 43548
rect 44300 43546 44356 43548
rect 44380 43546 44436 43548
rect 44460 43546 44516 43548
rect 44220 43494 44246 43546
rect 44246 43494 44276 43546
rect 44300 43494 44310 43546
rect 44310 43494 44356 43546
rect 44380 43494 44426 43546
rect 44426 43494 44436 43546
rect 44460 43494 44490 43546
rect 44490 43494 44516 43546
rect 44220 43492 44276 43494
rect 44300 43492 44356 43494
rect 44380 43492 44436 43494
rect 44460 43492 44516 43494
rect 44220 42458 44276 42460
rect 44300 42458 44356 42460
rect 44380 42458 44436 42460
rect 44460 42458 44516 42460
rect 44220 42406 44246 42458
rect 44246 42406 44276 42458
rect 44300 42406 44310 42458
rect 44310 42406 44356 42458
rect 44380 42406 44426 42458
rect 44426 42406 44436 42458
rect 44460 42406 44490 42458
rect 44490 42406 44516 42458
rect 44220 42404 44276 42406
rect 44300 42404 44356 42406
rect 44380 42404 44436 42406
rect 44460 42404 44516 42406
rect 44220 41370 44276 41372
rect 44300 41370 44356 41372
rect 44380 41370 44436 41372
rect 44460 41370 44516 41372
rect 44220 41318 44246 41370
rect 44246 41318 44276 41370
rect 44300 41318 44310 41370
rect 44310 41318 44356 41370
rect 44380 41318 44426 41370
rect 44426 41318 44436 41370
rect 44460 41318 44490 41370
rect 44490 41318 44516 41370
rect 44220 41316 44276 41318
rect 44300 41316 44356 41318
rect 44380 41316 44436 41318
rect 44460 41316 44516 41318
rect 44220 40282 44276 40284
rect 44300 40282 44356 40284
rect 44380 40282 44436 40284
rect 44460 40282 44516 40284
rect 44220 40230 44246 40282
rect 44246 40230 44276 40282
rect 44300 40230 44310 40282
rect 44310 40230 44356 40282
rect 44380 40230 44426 40282
rect 44426 40230 44436 40282
rect 44460 40230 44490 40282
rect 44490 40230 44516 40282
rect 44220 40228 44276 40230
rect 44300 40228 44356 40230
rect 44380 40228 44436 40230
rect 44460 40228 44516 40230
rect 44220 39194 44276 39196
rect 44300 39194 44356 39196
rect 44380 39194 44436 39196
rect 44460 39194 44516 39196
rect 44220 39142 44246 39194
rect 44246 39142 44276 39194
rect 44300 39142 44310 39194
rect 44310 39142 44356 39194
rect 44380 39142 44426 39194
rect 44426 39142 44436 39194
rect 44460 39142 44490 39194
rect 44490 39142 44516 39194
rect 44220 39140 44276 39142
rect 44300 39140 44356 39142
rect 44380 39140 44436 39142
rect 44460 39140 44516 39142
rect 44220 38106 44276 38108
rect 44300 38106 44356 38108
rect 44380 38106 44436 38108
rect 44460 38106 44516 38108
rect 44220 38054 44246 38106
rect 44246 38054 44276 38106
rect 44300 38054 44310 38106
rect 44310 38054 44356 38106
rect 44380 38054 44426 38106
rect 44426 38054 44436 38106
rect 44460 38054 44490 38106
rect 44490 38054 44516 38106
rect 44220 38052 44276 38054
rect 44300 38052 44356 38054
rect 44380 38052 44436 38054
rect 44460 38052 44516 38054
rect 44220 37018 44276 37020
rect 44300 37018 44356 37020
rect 44380 37018 44436 37020
rect 44460 37018 44516 37020
rect 44220 36966 44246 37018
rect 44246 36966 44276 37018
rect 44300 36966 44310 37018
rect 44310 36966 44356 37018
rect 44380 36966 44426 37018
rect 44426 36966 44436 37018
rect 44460 36966 44490 37018
rect 44490 36966 44516 37018
rect 44220 36964 44276 36966
rect 44300 36964 44356 36966
rect 44380 36964 44436 36966
rect 44460 36964 44516 36966
rect 44220 35930 44276 35932
rect 44300 35930 44356 35932
rect 44380 35930 44436 35932
rect 44460 35930 44516 35932
rect 44220 35878 44246 35930
rect 44246 35878 44276 35930
rect 44300 35878 44310 35930
rect 44310 35878 44356 35930
rect 44380 35878 44426 35930
rect 44426 35878 44436 35930
rect 44460 35878 44490 35930
rect 44490 35878 44516 35930
rect 44220 35876 44276 35878
rect 44300 35876 44356 35878
rect 44380 35876 44436 35878
rect 44460 35876 44516 35878
rect 44220 34842 44276 34844
rect 44300 34842 44356 34844
rect 44380 34842 44436 34844
rect 44460 34842 44516 34844
rect 44220 34790 44246 34842
rect 44246 34790 44276 34842
rect 44300 34790 44310 34842
rect 44310 34790 44356 34842
rect 44380 34790 44426 34842
rect 44426 34790 44436 34842
rect 44460 34790 44490 34842
rect 44490 34790 44516 34842
rect 44220 34788 44276 34790
rect 44300 34788 44356 34790
rect 44380 34788 44436 34790
rect 44460 34788 44516 34790
rect 44220 33754 44276 33756
rect 44300 33754 44356 33756
rect 44380 33754 44436 33756
rect 44460 33754 44516 33756
rect 44220 33702 44246 33754
rect 44246 33702 44276 33754
rect 44300 33702 44310 33754
rect 44310 33702 44356 33754
rect 44380 33702 44426 33754
rect 44426 33702 44436 33754
rect 44460 33702 44490 33754
rect 44490 33702 44516 33754
rect 44220 33700 44276 33702
rect 44300 33700 44356 33702
rect 44380 33700 44436 33702
rect 44460 33700 44516 33702
rect 44220 32666 44276 32668
rect 44300 32666 44356 32668
rect 44380 32666 44436 32668
rect 44460 32666 44516 32668
rect 44220 32614 44246 32666
rect 44246 32614 44276 32666
rect 44300 32614 44310 32666
rect 44310 32614 44356 32666
rect 44380 32614 44426 32666
rect 44426 32614 44436 32666
rect 44460 32614 44490 32666
rect 44490 32614 44516 32666
rect 44220 32612 44276 32614
rect 44300 32612 44356 32614
rect 44380 32612 44436 32614
rect 44460 32612 44516 32614
rect 44220 31578 44276 31580
rect 44300 31578 44356 31580
rect 44380 31578 44436 31580
rect 44460 31578 44516 31580
rect 44220 31526 44246 31578
rect 44246 31526 44276 31578
rect 44300 31526 44310 31578
rect 44310 31526 44356 31578
rect 44380 31526 44426 31578
rect 44426 31526 44436 31578
rect 44460 31526 44490 31578
rect 44490 31526 44516 31578
rect 44220 31524 44276 31526
rect 44300 31524 44356 31526
rect 44380 31524 44436 31526
rect 44460 31524 44516 31526
rect 44220 30490 44276 30492
rect 44300 30490 44356 30492
rect 44380 30490 44436 30492
rect 44460 30490 44516 30492
rect 44220 30438 44246 30490
rect 44246 30438 44276 30490
rect 44300 30438 44310 30490
rect 44310 30438 44356 30490
rect 44380 30438 44426 30490
rect 44426 30438 44436 30490
rect 44460 30438 44490 30490
rect 44490 30438 44516 30490
rect 44220 30436 44276 30438
rect 44300 30436 44356 30438
rect 44380 30436 44436 30438
rect 44460 30436 44516 30438
rect 44220 29402 44276 29404
rect 44300 29402 44356 29404
rect 44380 29402 44436 29404
rect 44460 29402 44516 29404
rect 44220 29350 44246 29402
rect 44246 29350 44276 29402
rect 44300 29350 44310 29402
rect 44310 29350 44356 29402
rect 44380 29350 44426 29402
rect 44426 29350 44436 29402
rect 44460 29350 44490 29402
rect 44490 29350 44516 29402
rect 44220 29348 44276 29350
rect 44300 29348 44356 29350
rect 44380 29348 44436 29350
rect 44460 29348 44516 29350
rect 44220 28314 44276 28316
rect 44300 28314 44356 28316
rect 44380 28314 44436 28316
rect 44460 28314 44516 28316
rect 44220 28262 44246 28314
rect 44246 28262 44276 28314
rect 44300 28262 44310 28314
rect 44310 28262 44356 28314
rect 44380 28262 44426 28314
rect 44426 28262 44436 28314
rect 44460 28262 44490 28314
rect 44490 28262 44516 28314
rect 44220 28260 44276 28262
rect 44300 28260 44356 28262
rect 44380 28260 44436 28262
rect 44460 28260 44516 28262
rect 44220 27226 44276 27228
rect 44300 27226 44356 27228
rect 44380 27226 44436 27228
rect 44460 27226 44516 27228
rect 44220 27174 44246 27226
rect 44246 27174 44276 27226
rect 44300 27174 44310 27226
rect 44310 27174 44356 27226
rect 44380 27174 44426 27226
rect 44426 27174 44436 27226
rect 44460 27174 44490 27226
rect 44490 27174 44516 27226
rect 44220 27172 44276 27174
rect 44300 27172 44356 27174
rect 44380 27172 44436 27174
rect 44460 27172 44516 27174
rect 44220 26138 44276 26140
rect 44300 26138 44356 26140
rect 44380 26138 44436 26140
rect 44460 26138 44516 26140
rect 44220 26086 44246 26138
rect 44246 26086 44276 26138
rect 44300 26086 44310 26138
rect 44310 26086 44356 26138
rect 44380 26086 44426 26138
rect 44426 26086 44436 26138
rect 44460 26086 44490 26138
rect 44490 26086 44516 26138
rect 44220 26084 44276 26086
rect 44300 26084 44356 26086
rect 44380 26084 44436 26086
rect 44460 26084 44516 26086
rect 44220 25050 44276 25052
rect 44300 25050 44356 25052
rect 44380 25050 44436 25052
rect 44460 25050 44516 25052
rect 44220 24998 44246 25050
rect 44246 24998 44276 25050
rect 44300 24998 44310 25050
rect 44310 24998 44356 25050
rect 44380 24998 44426 25050
rect 44426 24998 44436 25050
rect 44460 24998 44490 25050
rect 44490 24998 44516 25050
rect 44220 24996 44276 24998
rect 44300 24996 44356 24998
rect 44380 24996 44436 24998
rect 44460 24996 44516 24998
rect 44220 23962 44276 23964
rect 44300 23962 44356 23964
rect 44380 23962 44436 23964
rect 44460 23962 44516 23964
rect 44220 23910 44246 23962
rect 44246 23910 44276 23962
rect 44300 23910 44310 23962
rect 44310 23910 44356 23962
rect 44380 23910 44426 23962
rect 44426 23910 44436 23962
rect 44460 23910 44490 23962
rect 44490 23910 44516 23962
rect 44220 23908 44276 23910
rect 44300 23908 44356 23910
rect 44380 23908 44436 23910
rect 44460 23908 44516 23910
rect 44220 22874 44276 22876
rect 44300 22874 44356 22876
rect 44380 22874 44436 22876
rect 44460 22874 44516 22876
rect 44220 22822 44246 22874
rect 44246 22822 44276 22874
rect 44300 22822 44310 22874
rect 44310 22822 44356 22874
rect 44380 22822 44426 22874
rect 44426 22822 44436 22874
rect 44460 22822 44490 22874
rect 44490 22822 44516 22874
rect 44220 22820 44276 22822
rect 44300 22820 44356 22822
rect 44380 22820 44436 22822
rect 44460 22820 44516 22822
rect 44220 21786 44276 21788
rect 44300 21786 44356 21788
rect 44380 21786 44436 21788
rect 44460 21786 44516 21788
rect 44220 21734 44246 21786
rect 44246 21734 44276 21786
rect 44300 21734 44310 21786
rect 44310 21734 44356 21786
rect 44380 21734 44426 21786
rect 44426 21734 44436 21786
rect 44460 21734 44490 21786
rect 44490 21734 44516 21786
rect 44220 21732 44276 21734
rect 44300 21732 44356 21734
rect 44380 21732 44436 21734
rect 44460 21732 44516 21734
rect 44220 20698 44276 20700
rect 44300 20698 44356 20700
rect 44380 20698 44436 20700
rect 44460 20698 44516 20700
rect 44220 20646 44246 20698
rect 44246 20646 44276 20698
rect 44300 20646 44310 20698
rect 44310 20646 44356 20698
rect 44380 20646 44426 20698
rect 44426 20646 44436 20698
rect 44460 20646 44490 20698
rect 44490 20646 44516 20698
rect 44220 20644 44276 20646
rect 44300 20644 44356 20646
rect 44380 20644 44436 20646
rect 44460 20644 44516 20646
rect 44220 19610 44276 19612
rect 44300 19610 44356 19612
rect 44380 19610 44436 19612
rect 44460 19610 44516 19612
rect 44220 19558 44246 19610
rect 44246 19558 44276 19610
rect 44300 19558 44310 19610
rect 44310 19558 44356 19610
rect 44380 19558 44426 19610
rect 44426 19558 44436 19610
rect 44460 19558 44490 19610
rect 44490 19558 44516 19610
rect 44220 19556 44276 19558
rect 44300 19556 44356 19558
rect 44380 19556 44436 19558
rect 44460 19556 44516 19558
rect 44220 18522 44276 18524
rect 44300 18522 44356 18524
rect 44380 18522 44436 18524
rect 44460 18522 44516 18524
rect 44220 18470 44246 18522
rect 44246 18470 44276 18522
rect 44300 18470 44310 18522
rect 44310 18470 44356 18522
rect 44380 18470 44426 18522
rect 44426 18470 44436 18522
rect 44460 18470 44490 18522
rect 44490 18470 44516 18522
rect 44220 18468 44276 18470
rect 44300 18468 44356 18470
rect 44380 18468 44436 18470
rect 44460 18468 44516 18470
rect 44220 17434 44276 17436
rect 44300 17434 44356 17436
rect 44380 17434 44436 17436
rect 44460 17434 44516 17436
rect 44220 17382 44246 17434
rect 44246 17382 44276 17434
rect 44300 17382 44310 17434
rect 44310 17382 44356 17434
rect 44380 17382 44426 17434
rect 44426 17382 44436 17434
rect 44460 17382 44490 17434
rect 44490 17382 44516 17434
rect 44220 17380 44276 17382
rect 44300 17380 44356 17382
rect 44380 17380 44436 17382
rect 44460 17380 44516 17382
rect 43810 11328 43866 11384
rect 43626 9152 43682 9208
rect 44220 16346 44276 16348
rect 44300 16346 44356 16348
rect 44380 16346 44436 16348
rect 44460 16346 44516 16348
rect 44220 16294 44246 16346
rect 44246 16294 44276 16346
rect 44300 16294 44310 16346
rect 44310 16294 44356 16346
rect 44380 16294 44426 16346
rect 44426 16294 44436 16346
rect 44460 16294 44490 16346
rect 44490 16294 44516 16346
rect 44220 16292 44276 16294
rect 44300 16292 44356 16294
rect 44380 16292 44436 16294
rect 44460 16292 44516 16294
rect 44220 15258 44276 15260
rect 44300 15258 44356 15260
rect 44380 15258 44436 15260
rect 44460 15258 44516 15260
rect 44220 15206 44246 15258
rect 44246 15206 44276 15258
rect 44300 15206 44310 15258
rect 44310 15206 44356 15258
rect 44380 15206 44426 15258
rect 44426 15206 44436 15258
rect 44460 15206 44490 15258
rect 44490 15206 44516 15258
rect 44220 15204 44276 15206
rect 44300 15204 44356 15206
rect 44380 15204 44436 15206
rect 44460 15204 44516 15206
rect 44220 14170 44276 14172
rect 44300 14170 44356 14172
rect 44380 14170 44436 14172
rect 44460 14170 44516 14172
rect 44220 14118 44246 14170
rect 44246 14118 44276 14170
rect 44300 14118 44310 14170
rect 44310 14118 44356 14170
rect 44380 14118 44426 14170
rect 44426 14118 44436 14170
rect 44460 14118 44490 14170
rect 44490 14118 44516 14170
rect 44220 14116 44276 14118
rect 44300 14116 44356 14118
rect 44380 14116 44436 14118
rect 44460 14116 44516 14118
rect 44220 13082 44276 13084
rect 44300 13082 44356 13084
rect 44380 13082 44436 13084
rect 44460 13082 44516 13084
rect 44220 13030 44246 13082
rect 44246 13030 44276 13082
rect 44300 13030 44310 13082
rect 44310 13030 44356 13082
rect 44380 13030 44426 13082
rect 44426 13030 44436 13082
rect 44460 13030 44490 13082
rect 44490 13030 44516 13082
rect 44220 13028 44276 13030
rect 44300 13028 44356 13030
rect 44380 13028 44436 13030
rect 44460 13028 44516 13030
rect 44220 11994 44276 11996
rect 44300 11994 44356 11996
rect 44380 11994 44436 11996
rect 44460 11994 44516 11996
rect 44220 11942 44246 11994
rect 44246 11942 44276 11994
rect 44300 11942 44310 11994
rect 44310 11942 44356 11994
rect 44380 11942 44426 11994
rect 44426 11942 44436 11994
rect 44460 11942 44490 11994
rect 44490 11942 44516 11994
rect 44220 11940 44276 11942
rect 44300 11940 44356 11942
rect 44380 11940 44436 11942
rect 44460 11940 44516 11942
rect 44086 10920 44142 10976
rect 44220 10906 44276 10908
rect 44300 10906 44356 10908
rect 44380 10906 44436 10908
rect 44460 10906 44516 10908
rect 44220 10854 44246 10906
rect 44246 10854 44276 10906
rect 44300 10854 44310 10906
rect 44310 10854 44356 10906
rect 44380 10854 44426 10906
rect 44426 10854 44436 10906
rect 44460 10854 44490 10906
rect 44490 10854 44516 10906
rect 44220 10852 44276 10854
rect 44300 10852 44356 10854
rect 44380 10852 44436 10854
rect 44460 10852 44516 10854
rect 44220 9818 44276 9820
rect 44300 9818 44356 9820
rect 44380 9818 44436 9820
rect 44460 9818 44516 9820
rect 44220 9766 44246 9818
rect 44246 9766 44276 9818
rect 44300 9766 44310 9818
rect 44310 9766 44356 9818
rect 44380 9766 44426 9818
rect 44426 9766 44436 9818
rect 44460 9766 44490 9818
rect 44490 9766 44516 9818
rect 44220 9764 44276 9766
rect 44300 9764 44356 9766
rect 44380 9764 44436 9766
rect 44460 9764 44516 9766
rect 43994 9424 44050 9480
rect 43350 5344 43406 5400
rect 43350 4392 43406 4448
rect 43258 3984 43314 4040
rect 43166 2760 43222 2816
rect 43626 4664 43682 4720
rect 43534 2760 43590 2816
rect 44270 8880 44326 8936
rect 43718 3712 43774 3768
rect 43718 3032 43774 3088
rect 44220 8730 44276 8732
rect 44300 8730 44356 8732
rect 44380 8730 44436 8732
rect 44460 8730 44516 8732
rect 44220 8678 44246 8730
rect 44246 8678 44276 8730
rect 44300 8678 44310 8730
rect 44310 8678 44356 8730
rect 44380 8678 44426 8730
rect 44426 8678 44436 8730
rect 44460 8678 44490 8730
rect 44490 8678 44516 8730
rect 44220 8676 44276 8678
rect 44300 8676 44356 8678
rect 44380 8676 44436 8678
rect 44460 8676 44516 8678
rect 44220 7642 44276 7644
rect 44300 7642 44356 7644
rect 44380 7642 44436 7644
rect 44460 7642 44516 7644
rect 44220 7590 44246 7642
rect 44246 7590 44276 7642
rect 44300 7590 44310 7642
rect 44310 7590 44356 7642
rect 44380 7590 44426 7642
rect 44426 7590 44436 7642
rect 44460 7590 44490 7642
rect 44490 7590 44516 7642
rect 44220 7588 44276 7590
rect 44300 7588 44356 7590
rect 44380 7588 44436 7590
rect 44460 7588 44516 7590
rect 44220 6554 44276 6556
rect 44300 6554 44356 6556
rect 44380 6554 44436 6556
rect 44460 6554 44516 6556
rect 44220 6502 44246 6554
rect 44246 6502 44276 6554
rect 44300 6502 44310 6554
rect 44310 6502 44356 6554
rect 44380 6502 44426 6554
rect 44426 6502 44436 6554
rect 44460 6502 44490 6554
rect 44490 6502 44516 6554
rect 44220 6500 44276 6502
rect 44300 6500 44356 6502
rect 44380 6500 44436 6502
rect 44460 6500 44516 6502
rect 44220 5466 44276 5468
rect 44300 5466 44356 5468
rect 44380 5466 44436 5468
rect 44460 5466 44516 5468
rect 44220 5414 44246 5466
rect 44246 5414 44276 5466
rect 44300 5414 44310 5466
rect 44310 5414 44356 5466
rect 44380 5414 44426 5466
rect 44426 5414 44436 5466
rect 44460 5414 44490 5466
rect 44490 5414 44516 5466
rect 44220 5412 44276 5414
rect 44300 5412 44356 5414
rect 44380 5412 44436 5414
rect 44460 5412 44516 5414
rect 44178 4528 44234 4584
rect 44220 4378 44276 4380
rect 44300 4378 44356 4380
rect 44380 4378 44436 4380
rect 44460 4378 44516 4380
rect 44220 4326 44246 4378
rect 44246 4326 44276 4378
rect 44300 4326 44310 4378
rect 44310 4326 44356 4378
rect 44380 4326 44426 4378
rect 44426 4326 44436 4378
rect 44460 4326 44490 4378
rect 44490 4326 44516 4378
rect 44220 4324 44276 4326
rect 44300 4324 44356 4326
rect 44380 4324 44436 4326
rect 44460 4324 44516 4326
rect 44546 3576 44602 3632
rect 44220 3290 44276 3292
rect 44300 3290 44356 3292
rect 44380 3290 44436 3292
rect 44460 3290 44516 3292
rect 44220 3238 44246 3290
rect 44246 3238 44276 3290
rect 44300 3238 44310 3290
rect 44310 3238 44356 3290
rect 44380 3238 44426 3290
rect 44426 3238 44436 3290
rect 44460 3238 44490 3290
rect 44490 3238 44516 3290
rect 44220 3236 44276 3238
rect 44300 3236 44356 3238
rect 44380 3236 44436 3238
rect 44460 3236 44516 3238
rect 45374 11192 45430 11248
rect 44546 2760 44602 2816
rect 44220 2202 44276 2204
rect 44300 2202 44356 2204
rect 44380 2202 44436 2204
rect 44460 2202 44516 2204
rect 44220 2150 44246 2202
rect 44246 2150 44276 2202
rect 44300 2150 44310 2202
rect 44310 2150 44356 2202
rect 44380 2150 44426 2202
rect 44426 2150 44436 2202
rect 44460 2150 44490 2202
rect 44490 2150 44516 2202
rect 44220 2148 44276 2150
rect 44300 2148 44356 2150
rect 44380 2148 44436 2150
rect 44460 2148 44516 2150
rect 45098 8472 45154 8528
rect 45098 3440 45154 3496
rect 45466 3304 45522 3360
rect 45650 3612 45652 3632
rect 45652 3612 45704 3632
rect 45704 3612 45706 3632
rect 45650 3576 45706 3612
rect 46202 4392 46258 4448
rect 46662 5772 46718 5808
rect 46662 5752 46664 5772
rect 46664 5752 46716 5772
rect 46716 5752 46718 5772
rect 46938 12280 46994 12336
rect 46846 7792 46902 7848
rect 46570 3848 46626 3904
rect 47582 3168 47638 3224
rect 47858 3848 47914 3904
rect 47766 2896 47822 2952
rect 48502 4392 48558 4448
rect 48410 3440 48466 3496
rect 48502 2488 48558 2544
rect 48686 3032 48742 3088
rect 49220 62586 49276 62588
rect 49300 62586 49356 62588
rect 49380 62586 49436 62588
rect 49460 62586 49516 62588
rect 49220 62534 49246 62586
rect 49246 62534 49276 62586
rect 49300 62534 49310 62586
rect 49310 62534 49356 62586
rect 49380 62534 49426 62586
rect 49426 62534 49436 62586
rect 49460 62534 49490 62586
rect 49490 62534 49516 62586
rect 49220 62532 49276 62534
rect 49300 62532 49356 62534
rect 49380 62532 49436 62534
rect 49460 62532 49516 62534
rect 49220 61498 49276 61500
rect 49300 61498 49356 61500
rect 49380 61498 49436 61500
rect 49460 61498 49516 61500
rect 49220 61446 49246 61498
rect 49246 61446 49276 61498
rect 49300 61446 49310 61498
rect 49310 61446 49356 61498
rect 49380 61446 49426 61498
rect 49426 61446 49436 61498
rect 49460 61446 49490 61498
rect 49490 61446 49516 61498
rect 49220 61444 49276 61446
rect 49300 61444 49356 61446
rect 49380 61444 49436 61446
rect 49460 61444 49516 61446
rect 49220 60410 49276 60412
rect 49300 60410 49356 60412
rect 49380 60410 49436 60412
rect 49460 60410 49516 60412
rect 49220 60358 49246 60410
rect 49246 60358 49276 60410
rect 49300 60358 49310 60410
rect 49310 60358 49356 60410
rect 49380 60358 49426 60410
rect 49426 60358 49436 60410
rect 49460 60358 49490 60410
rect 49490 60358 49516 60410
rect 49220 60356 49276 60358
rect 49300 60356 49356 60358
rect 49380 60356 49436 60358
rect 49460 60356 49516 60358
rect 49220 59322 49276 59324
rect 49300 59322 49356 59324
rect 49380 59322 49436 59324
rect 49460 59322 49516 59324
rect 49220 59270 49246 59322
rect 49246 59270 49276 59322
rect 49300 59270 49310 59322
rect 49310 59270 49356 59322
rect 49380 59270 49426 59322
rect 49426 59270 49436 59322
rect 49460 59270 49490 59322
rect 49490 59270 49516 59322
rect 49220 59268 49276 59270
rect 49300 59268 49356 59270
rect 49380 59268 49436 59270
rect 49460 59268 49516 59270
rect 49220 58234 49276 58236
rect 49300 58234 49356 58236
rect 49380 58234 49436 58236
rect 49460 58234 49516 58236
rect 49220 58182 49246 58234
rect 49246 58182 49276 58234
rect 49300 58182 49310 58234
rect 49310 58182 49356 58234
rect 49380 58182 49426 58234
rect 49426 58182 49436 58234
rect 49460 58182 49490 58234
rect 49490 58182 49516 58234
rect 49220 58180 49276 58182
rect 49300 58180 49356 58182
rect 49380 58180 49436 58182
rect 49460 58180 49516 58182
rect 49220 57146 49276 57148
rect 49300 57146 49356 57148
rect 49380 57146 49436 57148
rect 49460 57146 49516 57148
rect 49220 57094 49246 57146
rect 49246 57094 49276 57146
rect 49300 57094 49310 57146
rect 49310 57094 49356 57146
rect 49380 57094 49426 57146
rect 49426 57094 49436 57146
rect 49460 57094 49490 57146
rect 49490 57094 49516 57146
rect 49220 57092 49276 57094
rect 49300 57092 49356 57094
rect 49380 57092 49436 57094
rect 49460 57092 49516 57094
rect 49220 56058 49276 56060
rect 49300 56058 49356 56060
rect 49380 56058 49436 56060
rect 49460 56058 49516 56060
rect 49220 56006 49246 56058
rect 49246 56006 49276 56058
rect 49300 56006 49310 56058
rect 49310 56006 49356 56058
rect 49380 56006 49426 56058
rect 49426 56006 49436 56058
rect 49460 56006 49490 56058
rect 49490 56006 49516 56058
rect 49220 56004 49276 56006
rect 49300 56004 49356 56006
rect 49380 56004 49436 56006
rect 49460 56004 49516 56006
rect 49220 54970 49276 54972
rect 49300 54970 49356 54972
rect 49380 54970 49436 54972
rect 49460 54970 49516 54972
rect 49220 54918 49246 54970
rect 49246 54918 49276 54970
rect 49300 54918 49310 54970
rect 49310 54918 49356 54970
rect 49380 54918 49426 54970
rect 49426 54918 49436 54970
rect 49460 54918 49490 54970
rect 49490 54918 49516 54970
rect 49220 54916 49276 54918
rect 49300 54916 49356 54918
rect 49380 54916 49436 54918
rect 49460 54916 49516 54918
rect 49220 53882 49276 53884
rect 49300 53882 49356 53884
rect 49380 53882 49436 53884
rect 49460 53882 49516 53884
rect 49220 53830 49246 53882
rect 49246 53830 49276 53882
rect 49300 53830 49310 53882
rect 49310 53830 49356 53882
rect 49380 53830 49426 53882
rect 49426 53830 49436 53882
rect 49460 53830 49490 53882
rect 49490 53830 49516 53882
rect 49220 53828 49276 53830
rect 49300 53828 49356 53830
rect 49380 53828 49436 53830
rect 49460 53828 49516 53830
rect 49220 52794 49276 52796
rect 49300 52794 49356 52796
rect 49380 52794 49436 52796
rect 49460 52794 49516 52796
rect 49220 52742 49246 52794
rect 49246 52742 49276 52794
rect 49300 52742 49310 52794
rect 49310 52742 49356 52794
rect 49380 52742 49426 52794
rect 49426 52742 49436 52794
rect 49460 52742 49490 52794
rect 49490 52742 49516 52794
rect 49220 52740 49276 52742
rect 49300 52740 49356 52742
rect 49380 52740 49436 52742
rect 49460 52740 49516 52742
rect 49220 51706 49276 51708
rect 49300 51706 49356 51708
rect 49380 51706 49436 51708
rect 49460 51706 49516 51708
rect 49220 51654 49246 51706
rect 49246 51654 49276 51706
rect 49300 51654 49310 51706
rect 49310 51654 49356 51706
rect 49380 51654 49426 51706
rect 49426 51654 49436 51706
rect 49460 51654 49490 51706
rect 49490 51654 49516 51706
rect 49220 51652 49276 51654
rect 49300 51652 49356 51654
rect 49380 51652 49436 51654
rect 49460 51652 49516 51654
rect 49220 50618 49276 50620
rect 49300 50618 49356 50620
rect 49380 50618 49436 50620
rect 49460 50618 49516 50620
rect 49220 50566 49246 50618
rect 49246 50566 49276 50618
rect 49300 50566 49310 50618
rect 49310 50566 49356 50618
rect 49380 50566 49426 50618
rect 49426 50566 49436 50618
rect 49460 50566 49490 50618
rect 49490 50566 49516 50618
rect 49220 50564 49276 50566
rect 49300 50564 49356 50566
rect 49380 50564 49436 50566
rect 49460 50564 49516 50566
rect 49220 49530 49276 49532
rect 49300 49530 49356 49532
rect 49380 49530 49436 49532
rect 49460 49530 49516 49532
rect 49220 49478 49246 49530
rect 49246 49478 49276 49530
rect 49300 49478 49310 49530
rect 49310 49478 49356 49530
rect 49380 49478 49426 49530
rect 49426 49478 49436 49530
rect 49460 49478 49490 49530
rect 49490 49478 49516 49530
rect 49220 49476 49276 49478
rect 49300 49476 49356 49478
rect 49380 49476 49436 49478
rect 49460 49476 49516 49478
rect 49220 48442 49276 48444
rect 49300 48442 49356 48444
rect 49380 48442 49436 48444
rect 49460 48442 49516 48444
rect 49220 48390 49246 48442
rect 49246 48390 49276 48442
rect 49300 48390 49310 48442
rect 49310 48390 49356 48442
rect 49380 48390 49426 48442
rect 49426 48390 49436 48442
rect 49460 48390 49490 48442
rect 49490 48390 49516 48442
rect 49220 48388 49276 48390
rect 49300 48388 49356 48390
rect 49380 48388 49436 48390
rect 49460 48388 49516 48390
rect 49220 47354 49276 47356
rect 49300 47354 49356 47356
rect 49380 47354 49436 47356
rect 49460 47354 49516 47356
rect 49220 47302 49246 47354
rect 49246 47302 49276 47354
rect 49300 47302 49310 47354
rect 49310 47302 49356 47354
rect 49380 47302 49426 47354
rect 49426 47302 49436 47354
rect 49460 47302 49490 47354
rect 49490 47302 49516 47354
rect 49220 47300 49276 47302
rect 49300 47300 49356 47302
rect 49380 47300 49436 47302
rect 49460 47300 49516 47302
rect 49220 46266 49276 46268
rect 49300 46266 49356 46268
rect 49380 46266 49436 46268
rect 49460 46266 49516 46268
rect 49220 46214 49246 46266
rect 49246 46214 49276 46266
rect 49300 46214 49310 46266
rect 49310 46214 49356 46266
rect 49380 46214 49426 46266
rect 49426 46214 49436 46266
rect 49460 46214 49490 46266
rect 49490 46214 49516 46266
rect 49220 46212 49276 46214
rect 49300 46212 49356 46214
rect 49380 46212 49436 46214
rect 49460 46212 49516 46214
rect 49220 45178 49276 45180
rect 49300 45178 49356 45180
rect 49380 45178 49436 45180
rect 49460 45178 49516 45180
rect 49220 45126 49246 45178
rect 49246 45126 49276 45178
rect 49300 45126 49310 45178
rect 49310 45126 49356 45178
rect 49380 45126 49426 45178
rect 49426 45126 49436 45178
rect 49460 45126 49490 45178
rect 49490 45126 49516 45178
rect 49220 45124 49276 45126
rect 49300 45124 49356 45126
rect 49380 45124 49436 45126
rect 49460 45124 49516 45126
rect 49220 44090 49276 44092
rect 49300 44090 49356 44092
rect 49380 44090 49436 44092
rect 49460 44090 49516 44092
rect 49220 44038 49246 44090
rect 49246 44038 49276 44090
rect 49300 44038 49310 44090
rect 49310 44038 49356 44090
rect 49380 44038 49426 44090
rect 49426 44038 49436 44090
rect 49460 44038 49490 44090
rect 49490 44038 49516 44090
rect 49220 44036 49276 44038
rect 49300 44036 49356 44038
rect 49380 44036 49436 44038
rect 49460 44036 49516 44038
rect 49220 43002 49276 43004
rect 49300 43002 49356 43004
rect 49380 43002 49436 43004
rect 49460 43002 49516 43004
rect 49220 42950 49246 43002
rect 49246 42950 49276 43002
rect 49300 42950 49310 43002
rect 49310 42950 49356 43002
rect 49380 42950 49426 43002
rect 49426 42950 49436 43002
rect 49460 42950 49490 43002
rect 49490 42950 49516 43002
rect 49220 42948 49276 42950
rect 49300 42948 49356 42950
rect 49380 42948 49436 42950
rect 49460 42948 49516 42950
rect 49220 41914 49276 41916
rect 49300 41914 49356 41916
rect 49380 41914 49436 41916
rect 49460 41914 49516 41916
rect 49220 41862 49246 41914
rect 49246 41862 49276 41914
rect 49300 41862 49310 41914
rect 49310 41862 49356 41914
rect 49380 41862 49426 41914
rect 49426 41862 49436 41914
rect 49460 41862 49490 41914
rect 49490 41862 49516 41914
rect 49220 41860 49276 41862
rect 49300 41860 49356 41862
rect 49380 41860 49436 41862
rect 49460 41860 49516 41862
rect 49220 40826 49276 40828
rect 49300 40826 49356 40828
rect 49380 40826 49436 40828
rect 49460 40826 49516 40828
rect 49220 40774 49246 40826
rect 49246 40774 49276 40826
rect 49300 40774 49310 40826
rect 49310 40774 49356 40826
rect 49380 40774 49426 40826
rect 49426 40774 49436 40826
rect 49460 40774 49490 40826
rect 49490 40774 49516 40826
rect 49220 40772 49276 40774
rect 49300 40772 49356 40774
rect 49380 40772 49436 40774
rect 49460 40772 49516 40774
rect 49220 39738 49276 39740
rect 49300 39738 49356 39740
rect 49380 39738 49436 39740
rect 49460 39738 49516 39740
rect 49220 39686 49246 39738
rect 49246 39686 49276 39738
rect 49300 39686 49310 39738
rect 49310 39686 49356 39738
rect 49380 39686 49426 39738
rect 49426 39686 49436 39738
rect 49460 39686 49490 39738
rect 49490 39686 49516 39738
rect 49220 39684 49276 39686
rect 49300 39684 49356 39686
rect 49380 39684 49436 39686
rect 49460 39684 49516 39686
rect 49220 38650 49276 38652
rect 49300 38650 49356 38652
rect 49380 38650 49436 38652
rect 49460 38650 49516 38652
rect 49220 38598 49246 38650
rect 49246 38598 49276 38650
rect 49300 38598 49310 38650
rect 49310 38598 49356 38650
rect 49380 38598 49426 38650
rect 49426 38598 49436 38650
rect 49460 38598 49490 38650
rect 49490 38598 49516 38650
rect 49220 38596 49276 38598
rect 49300 38596 49356 38598
rect 49380 38596 49436 38598
rect 49460 38596 49516 38598
rect 49220 37562 49276 37564
rect 49300 37562 49356 37564
rect 49380 37562 49436 37564
rect 49460 37562 49516 37564
rect 49220 37510 49246 37562
rect 49246 37510 49276 37562
rect 49300 37510 49310 37562
rect 49310 37510 49356 37562
rect 49380 37510 49426 37562
rect 49426 37510 49436 37562
rect 49460 37510 49490 37562
rect 49490 37510 49516 37562
rect 49220 37508 49276 37510
rect 49300 37508 49356 37510
rect 49380 37508 49436 37510
rect 49460 37508 49516 37510
rect 49220 36474 49276 36476
rect 49300 36474 49356 36476
rect 49380 36474 49436 36476
rect 49460 36474 49516 36476
rect 49220 36422 49246 36474
rect 49246 36422 49276 36474
rect 49300 36422 49310 36474
rect 49310 36422 49356 36474
rect 49380 36422 49426 36474
rect 49426 36422 49436 36474
rect 49460 36422 49490 36474
rect 49490 36422 49516 36474
rect 49220 36420 49276 36422
rect 49300 36420 49356 36422
rect 49380 36420 49436 36422
rect 49460 36420 49516 36422
rect 49220 35386 49276 35388
rect 49300 35386 49356 35388
rect 49380 35386 49436 35388
rect 49460 35386 49516 35388
rect 49220 35334 49246 35386
rect 49246 35334 49276 35386
rect 49300 35334 49310 35386
rect 49310 35334 49356 35386
rect 49380 35334 49426 35386
rect 49426 35334 49436 35386
rect 49460 35334 49490 35386
rect 49490 35334 49516 35386
rect 49220 35332 49276 35334
rect 49300 35332 49356 35334
rect 49380 35332 49436 35334
rect 49460 35332 49516 35334
rect 49220 34298 49276 34300
rect 49300 34298 49356 34300
rect 49380 34298 49436 34300
rect 49460 34298 49516 34300
rect 49220 34246 49246 34298
rect 49246 34246 49276 34298
rect 49300 34246 49310 34298
rect 49310 34246 49356 34298
rect 49380 34246 49426 34298
rect 49426 34246 49436 34298
rect 49460 34246 49490 34298
rect 49490 34246 49516 34298
rect 49220 34244 49276 34246
rect 49300 34244 49356 34246
rect 49380 34244 49436 34246
rect 49460 34244 49516 34246
rect 49220 33210 49276 33212
rect 49300 33210 49356 33212
rect 49380 33210 49436 33212
rect 49460 33210 49516 33212
rect 49220 33158 49246 33210
rect 49246 33158 49276 33210
rect 49300 33158 49310 33210
rect 49310 33158 49356 33210
rect 49380 33158 49426 33210
rect 49426 33158 49436 33210
rect 49460 33158 49490 33210
rect 49490 33158 49516 33210
rect 49220 33156 49276 33158
rect 49300 33156 49356 33158
rect 49380 33156 49436 33158
rect 49460 33156 49516 33158
rect 49220 32122 49276 32124
rect 49300 32122 49356 32124
rect 49380 32122 49436 32124
rect 49460 32122 49516 32124
rect 49220 32070 49246 32122
rect 49246 32070 49276 32122
rect 49300 32070 49310 32122
rect 49310 32070 49356 32122
rect 49380 32070 49426 32122
rect 49426 32070 49436 32122
rect 49460 32070 49490 32122
rect 49490 32070 49516 32122
rect 49220 32068 49276 32070
rect 49300 32068 49356 32070
rect 49380 32068 49436 32070
rect 49460 32068 49516 32070
rect 49220 31034 49276 31036
rect 49300 31034 49356 31036
rect 49380 31034 49436 31036
rect 49460 31034 49516 31036
rect 49220 30982 49246 31034
rect 49246 30982 49276 31034
rect 49300 30982 49310 31034
rect 49310 30982 49356 31034
rect 49380 30982 49426 31034
rect 49426 30982 49436 31034
rect 49460 30982 49490 31034
rect 49490 30982 49516 31034
rect 49220 30980 49276 30982
rect 49300 30980 49356 30982
rect 49380 30980 49436 30982
rect 49460 30980 49516 30982
rect 49220 29946 49276 29948
rect 49300 29946 49356 29948
rect 49380 29946 49436 29948
rect 49460 29946 49516 29948
rect 49220 29894 49246 29946
rect 49246 29894 49276 29946
rect 49300 29894 49310 29946
rect 49310 29894 49356 29946
rect 49380 29894 49426 29946
rect 49426 29894 49436 29946
rect 49460 29894 49490 29946
rect 49490 29894 49516 29946
rect 49220 29892 49276 29894
rect 49300 29892 49356 29894
rect 49380 29892 49436 29894
rect 49460 29892 49516 29894
rect 49220 28858 49276 28860
rect 49300 28858 49356 28860
rect 49380 28858 49436 28860
rect 49460 28858 49516 28860
rect 49220 28806 49246 28858
rect 49246 28806 49276 28858
rect 49300 28806 49310 28858
rect 49310 28806 49356 28858
rect 49380 28806 49426 28858
rect 49426 28806 49436 28858
rect 49460 28806 49490 28858
rect 49490 28806 49516 28858
rect 49220 28804 49276 28806
rect 49300 28804 49356 28806
rect 49380 28804 49436 28806
rect 49460 28804 49516 28806
rect 49220 27770 49276 27772
rect 49300 27770 49356 27772
rect 49380 27770 49436 27772
rect 49460 27770 49516 27772
rect 49220 27718 49246 27770
rect 49246 27718 49276 27770
rect 49300 27718 49310 27770
rect 49310 27718 49356 27770
rect 49380 27718 49426 27770
rect 49426 27718 49436 27770
rect 49460 27718 49490 27770
rect 49490 27718 49516 27770
rect 49220 27716 49276 27718
rect 49300 27716 49356 27718
rect 49380 27716 49436 27718
rect 49460 27716 49516 27718
rect 49220 26682 49276 26684
rect 49300 26682 49356 26684
rect 49380 26682 49436 26684
rect 49460 26682 49516 26684
rect 49220 26630 49246 26682
rect 49246 26630 49276 26682
rect 49300 26630 49310 26682
rect 49310 26630 49356 26682
rect 49380 26630 49426 26682
rect 49426 26630 49436 26682
rect 49460 26630 49490 26682
rect 49490 26630 49516 26682
rect 49220 26628 49276 26630
rect 49300 26628 49356 26630
rect 49380 26628 49436 26630
rect 49460 26628 49516 26630
rect 49220 25594 49276 25596
rect 49300 25594 49356 25596
rect 49380 25594 49436 25596
rect 49460 25594 49516 25596
rect 49220 25542 49246 25594
rect 49246 25542 49276 25594
rect 49300 25542 49310 25594
rect 49310 25542 49356 25594
rect 49380 25542 49426 25594
rect 49426 25542 49436 25594
rect 49460 25542 49490 25594
rect 49490 25542 49516 25594
rect 49220 25540 49276 25542
rect 49300 25540 49356 25542
rect 49380 25540 49436 25542
rect 49460 25540 49516 25542
rect 49220 24506 49276 24508
rect 49300 24506 49356 24508
rect 49380 24506 49436 24508
rect 49460 24506 49516 24508
rect 49220 24454 49246 24506
rect 49246 24454 49276 24506
rect 49300 24454 49310 24506
rect 49310 24454 49356 24506
rect 49380 24454 49426 24506
rect 49426 24454 49436 24506
rect 49460 24454 49490 24506
rect 49490 24454 49516 24506
rect 49220 24452 49276 24454
rect 49300 24452 49356 24454
rect 49380 24452 49436 24454
rect 49460 24452 49516 24454
rect 49220 23418 49276 23420
rect 49300 23418 49356 23420
rect 49380 23418 49436 23420
rect 49460 23418 49516 23420
rect 49220 23366 49246 23418
rect 49246 23366 49276 23418
rect 49300 23366 49310 23418
rect 49310 23366 49356 23418
rect 49380 23366 49426 23418
rect 49426 23366 49436 23418
rect 49460 23366 49490 23418
rect 49490 23366 49516 23418
rect 49220 23364 49276 23366
rect 49300 23364 49356 23366
rect 49380 23364 49436 23366
rect 49460 23364 49516 23366
rect 49220 22330 49276 22332
rect 49300 22330 49356 22332
rect 49380 22330 49436 22332
rect 49460 22330 49516 22332
rect 49220 22278 49246 22330
rect 49246 22278 49276 22330
rect 49300 22278 49310 22330
rect 49310 22278 49356 22330
rect 49380 22278 49426 22330
rect 49426 22278 49436 22330
rect 49460 22278 49490 22330
rect 49490 22278 49516 22330
rect 49220 22276 49276 22278
rect 49300 22276 49356 22278
rect 49380 22276 49436 22278
rect 49460 22276 49516 22278
rect 49220 21242 49276 21244
rect 49300 21242 49356 21244
rect 49380 21242 49436 21244
rect 49460 21242 49516 21244
rect 49220 21190 49246 21242
rect 49246 21190 49276 21242
rect 49300 21190 49310 21242
rect 49310 21190 49356 21242
rect 49380 21190 49426 21242
rect 49426 21190 49436 21242
rect 49460 21190 49490 21242
rect 49490 21190 49516 21242
rect 49220 21188 49276 21190
rect 49300 21188 49356 21190
rect 49380 21188 49436 21190
rect 49460 21188 49516 21190
rect 49220 20154 49276 20156
rect 49300 20154 49356 20156
rect 49380 20154 49436 20156
rect 49460 20154 49516 20156
rect 49220 20102 49246 20154
rect 49246 20102 49276 20154
rect 49300 20102 49310 20154
rect 49310 20102 49356 20154
rect 49380 20102 49426 20154
rect 49426 20102 49436 20154
rect 49460 20102 49490 20154
rect 49490 20102 49516 20154
rect 49220 20100 49276 20102
rect 49300 20100 49356 20102
rect 49380 20100 49436 20102
rect 49460 20100 49516 20102
rect 49220 19066 49276 19068
rect 49300 19066 49356 19068
rect 49380 19066 49436 19068
rect 49460 19066 49516 19068
rect 49220 19014 49246 19066
rect 49246 19014 49276 19066
rect 49300 19014 49310 19066
rect 49310 19014 49356 19066
rect 49380 19014 49426 19066
rect 49426 19014 49436 19066
rect 49460 19014 49490 19066
rect 49490 19014 49516 19066
rect 49220 19012 49276 19014
rect 49300 19012 49356 19014
rect 49380 19012 49436 19014
rect 49460 19012 49516 19014
rect 49220 17978 49276 17980
rect 49300 17978 49356 17980
rect 49380 17978 49436 17980
rect 49460 17978 49516 17980
rect 49220 17926 49246 17978
rect 49246 17926 49276 17978
rect 49300 17926 49310 17978
rect 49310 17926 49356 17978
rect 49380 17926 49426 17978
rect 49426 17926 49436 17978
rect 49460 17926 49490 17978
rect 49490 17926 49516 17978
rect 49220 17924 49276 17926
rect 49300 17924 49356 17926
rect 49380 17924 49436 17926
rect 49460 17924 49516 17926
rect 49220 16890 49276 16892
rect 49300 16890 49356 16892
rect 49380 16890 49436 16892
rect 49460 16890 49516 16892
rect 49220 16838 49246 16890
rect 49246 16838 49276 16890
rect 49300 16838 49310 16890
rect 49310 16838 49356 16890
rect 49380 16838 49426 16890
rect 49426 16838 49436 16890
rect 49460 16838 49490 16890
rect 49490 16838 49516 16890
rect 49220 16836 49276 16838
rect 49300 16836 49356 16838
rect 49380 16836 49436 16838
rect 49460 16836 49516 16838
rect 49220 15802 49276 15804
rect 49300 15802 49356 15804
rect 49380 15802 49436 15804
rect 49460 15802 49516 15804
rect 49220 15750 49246 15802
rect 49246 15750 49276 15802
rect 49300 15750 49310 15802
rect 49310 15750 49356 15802
rect 49380 15750 49426 15802
rect 49426 15750 49436 15802
rect 49460 15750 49490 15802
rect 49490 15750 49516 15802
rect 49220 15748 49276 15750
rect 49300 15748 49356 15750
rect 49380 15748 49436 15750
rect 49460 15748 49516 15750
rect 49220 14714 49276 14716
rect 49300 14714 49356 14716
rect 49380 14714 49436 14716
rect 49460 14714 49516 14716
rect 49220 14662 49246 14714
rect 49246 14662 49276 14714
rect 49300 14662 49310 14714
rect 49310 14662 49356 14714
rect 49380 14662 49426 14714
rect 49426 14662 49436 14714
rect 49460 14662 49490 14714
rect 49490 14662 49516 14714
rect 49220 14660 49276 14662
rect 49300 14660 49356 14662
rect 49380 14660 49436 14662
rect 49460 14660 49516 14662
rect 49220 13626 49276 13628
rect 49300 13626 49356 13628
rect 49380 13626 49436 13628
rect 49460 13626 49516 13628
rect 49220 13574 49246 13626
rect 49246 13574 49276 13626
rect 49300 13574 49310 13626
rect 49310 13574 49356 13626
rect 49380 13574 49426 13626
rect 49426 13574 49436 13626
rect 49460 13574 49490 13626
rect 49490 13574 49516 13626
rect 49220 13572 49276 13574
rect 49300 13572 49356 13574
rect 49380 13572 49436 13574
rect 49460 13572 49516 13574
rect 49220 12538 49276 12540
rect 49300 12538 49356 12540
rect 49380 12538 49436 12540
rect 49460 12538 49516 12540
rect 49220 12486 49246 12538
rect 49246 12486 49276 12538
rect 49300 12486 49310 12538
rect 49310 12486 49356 12538
rect 49380 12486 49426 12538
rect 49426 12486 49436 12538
rect 49460 12486 49490 12538
rect 49490 12486 49516 12538
rect 49220 12484 49276 12486
rect 49300 12484 49356 12486
rect 49380 12484 49436 12486
rect 49460 12484 49516 12486
rect 49220 11450 49276 11452
rect 49300 11450 49356 11452
rect 49380 11450 49436 11452
rect 49460 11450 49516 11452
rect 49220 11398 49246 11450
rect 49246 11398 49276 11450
rect 49300 11398 49310 11450
rect 49310 11398 49356 11450
rect 49380 11398 49426 11450
rect 49426 11398 49436 11450
rect 49460 11398 49490 11450
rect 49490 11398 49516 11450
rect 49220 11396 49276 11398
rect 49300 11396 49356 11398
rect 49380 11396 49436 11398
rect 49460 11396 49516 11398
rect 49220 10362 49276 10364
rect 49300 10362 49356 10364
rect 49380 10362 49436 10364
rect 49460 10362 49516 10364
rect 49220 10310 49246 10362
rect 49246 10310 49276 10362
rect 49300 10310 49310 10362
rect 49310 10310 49356 10362
rect 49380 10310 49426 10362
rect 49426 10310 49436 10362
rect 49460 10310 49490 10362
rect 49490 10310 49516 10362
rect 49220 10308 49276 10310
rect 49300 10308 49356 10310
rect 49380 10308 49436 10310
rect 49460 10308 49516 10310
rect 49220 9274 49276 9276
rect 49300 9274 49356 9276
rect 49380 9274 49436 9276
rect 49460 9274 49516 9276
rect 49220 9222 49246 9274
rect 49246 9222 49276 9274
rect 49300 9222 49310 9274
rect 49310 9222 49356 9274
rect 49380 9222 49426 9274
rect 49426 9222 49436 9274
rect 49460 9222 49490 9274
rect 49490 9222 49516 9274
rect 49220 9220 49276 9222
rect 49300 9220 49356 9222
rect 49380 9220 49436 9222
rect 49460 9220 49516 9222
rect 49220 8186 49276 8188
rect 49300 8186 49356 8188
rect 49380 8186 49436 8188
rect 49460 8186 49516 8188
rect 49220 8134 49246 8186
rect 49246 8134 49276 8186
rect 49300 8134 49310 8186
rect 49310 8134 49356 8186
rect 49380 8134 49426 8186
rect 49426 8134 49436 8186
rect 49460 8134 49490 8186
rect 49490 8134 49516 8186
rect 49220 8132 49276 8134
rect 49300 8132 49356 8134
rect 49380 8132 49436 8134
rect 49460 8132 49516 8134
rect 49220 7098 49276 7100
rect 49300 7098 49356 7100
rect 49380 7098 49436 7100
rect 49460 7098 49516 7100
rect 49220 7046 49246 7098
rect 49246 7046 49276 7098
rect 49300 7046 49310 7098
rect 49310 7046 49356 7098
rect 49380 7046 49426 7098
rect 49426 7046 49436 7098
rect 49460 7046 49490 7098
rect 49490 7046 49516 7098
rect 49220 7044 49276 7046
rect 49300 7044 49356 7046
rect 49380 7044 49436 7046
rect 49460 7044 49516 7046
rect 49220 6010 49276 6012
rect 49300 6010 49356 6012
rect 49380 6010 49436 6012
rect 49460 6010 49516 6012
rect 49220 5958 49246 6010
rect 49246 5958 49276 6010
rect 49300 5958 49310 6010
rect 49310 5958 49356 6010
rect 49380 5958 49426 6010
rect 49426 5958 49436 6010
rect 49460 5958 49490 6010
rect 49490 5958 49516 6010
rect 49220 5956 49276 5958
rect 49300 5956 49356 5958
rect 49380 5956 49436 5958
rect 49460 5956 49516 5958
rect 49220 4922 49276 4924
rect 49300 4922 49356 4924
rect 49380 4922 49436 4924
rect 49460 4922 49516 4924
rect 49220 4870 49246 4922
rect 49246 4870 49276 4922
rect 49300 4870 49310 4922
rect 49310 4870 49356 4922
rect 49380 4870 49426 4922
rect 49426 4870 49436 4922
rect 49460 4870 49490 4922
rect 49490 4870 49516 4922
rect 49220 4868 49276 4870
rect 49300 4868 49356 4870
rect 49380 4868 49436 4870
rect 49460 4868 49516 4870
rect 49220 3834 49276 3836
rect 49300 3834 49356 3836
rect 49380 3834 49436 3836
rect 49460 3834 49516 3836
rect 49220 3782 49246 3834
rect 49246 3782 49276 3834
rect 49300 3782 49310 3834
rect 49310 3782 49356 3834
rect 49380 3782 49426 3834
rect 49426 3782 49436 3834
rect 49460 3782 49490 3834
rect 49490 3782 49516 3834
rect 49220 3780 49276 3782
rect 49300 3780 49356 3782
rect 49380 3780 49436 3782
rect 49460 3780 49516 3782
rect 48870 2352 48926 2408
rect 49054 2760 49110 2816
rect 49220 2746 49276 2748
rect 49300 2746 49356 2748
rect 49380 2746 49436 2748
rect 49460 2746 49516 2748
rect 49220 2694 49246 2746
rect 49246 2694 49276 2746
rect 49300 2694 49310 2746
rect 49310 2694 49356 2746
rect 49380 2694 49426 2746
rect 49426 2694 49436 2746
rect 49460 2694 49490 2746
rect 49490 2694 49516 2746
rect 49220 2692 49276 2694
rect 49300 2692 49356 2694
rect 49380 2692 49436 2694
rect 49460 2692 49516 2694
rect 49422 2216 49478 2272
rect 49882 4020 49884 4040
rect 49884 4020 49936 4040
rect 49936 4020 49938 4040
rect 49882 3984 49938 4020
rect 49882 3848 49938 3904
rect 49790 2488 49846 2544
rect 49974 2896 50030 2952
rect 54220 66394 54276 66396
rect 54300 66394 54356 66396
rect 54380 66394 54436 66396
rect 54460 66394 54516 66396
rect 54220 66342 54246 66394
rect 54246 66342 54276 66394
rect 54300 66342 54310 66394
rect 54310 66342 54356 66394
rect 54380 66342 54426 66394
rect 54426 66342 54436 66394
rect 54460 66342 54490 66394
rect 54490 66342 54516 66394
rect 54220 66340 54276 66342
rect 54300 66340 54356 66342
rect 54380 66340 54436 66342
rect 54460 66340 54516 66342
rect 54220 65306 54276 65308
rect 54300 65306 54356 65308
rect 54380 65306 54436 65308
rect 54460 65306 54516 65308
rect 54220 65254 54246 65306
rect 54246 65254 54276 65306
rect 54300 65254 54310 65306
rect 54310 65254 54356 65306
rect 54380 65254 54426 65306
rect 54426 65254 54436 65306
rect 54460 65254 54490 65306
rect 54490 65254 54516 65306
rect 54220 65252 54276 65254
rect 54300 65252 54356 65254
rect 54380 65252 54436 65254
rect 54460 65252 54516 65254
rect 54220 64218 54276 64220
rect 54300 64218 54356 64220
rect 54380 64218 54436 64220
rect 54460 64218 54516 64220
rect 54220 64166 54246 64218
rect 54246 64166 54276 64218
rect 54300 64166 54310 64218
rect 54310 64166 54356 64218
rect 54380 64166 54426 64218
rect 54426 64166 54436 64218
rect 54460 64166 54490 64218
rect 54490 64166 54516 64218
rect 54220 64164 54276 64166
rect 54300 64164 54356 64166
rect 54380 64164 54436 64166
rect 54460 64164 54516 64166
rect 54220 63130 54276 63132
rect 54300 63130 54356 63132
rect 54380 63130 54436 63132
rect 54460 63130 54516 63132
rect 54220 63078 54246 63130
rect 54246 63078 54276 63130
rect 54300 63078 54310 63130
rect 54310 63078 54356 63130
rect 54380 63078 54426 63130
rect 54426 63078 54436 63130
rect 54460 63078 54490 63130
rect 54490 63078 54516 63130
rect 54220 63076 54276 63078
rect 54300 63076 54356 63078
rect 54380 63076 54436 63078
rect 54460 63076 54516 63078
rect 54220 62042 54276 62044
rect 54300 62042 54356 62044
rect 54380 62042 54436 62044
rect 54460 62042 54516 62044
rect 54220 61990 54246 62042
rect 54246 61990 54276 62042
rect 54300 61990 54310 62042
rect 54310 61990 54356 62042
rect 54380 61990 54426 62042
rect 54426 61990 54436 62042
rect 54460 61990 54490 62042
rect 54490 61990 54516 62042
rect 54220 61988 54276 61990
rect 54300 61988 54356 61990
rect 54380 61988 54436 61990
rect 54460 61988 54516 61990
rect 54220 60954 54276 60956
rect 54300 60954 54356 60956
rect 54380 60954 54436 60956
rect 54460 60954 54516 60956
rect 54220 60902 54246 60954
rect 54246 60902 54276 60954
rect 54300 60902 54310 60954
rect 54310 60902 54356 60954
rect 54380 60902 54426 60954
rect 54426 60902 54436 60954
rect 54460 60902 54490 60954
rect 54490 60902 54516 60954
rect 54220 60900 54276 60902
rect 54300 60900 54356 60902
rect 54380 60900 54436 60902
rect 54460 60900 54516 60902
rect 50710 3848 50766 3904
rect 50894 3168 50950 3224
rect 51078 3168 51134 3224
rect 54220 59866 54276 59868
rect 54300 59866 54356 59868
rect 54380 59866 54436 59868
rect 54460 59866 54516 59868
rect 54220 59814 54246 59866
rect 54246 59814 54276 59866
rect 54300 59814 54310 59866
rect 54310 59814 54356 59866
rect 54380 59814 54426 59866
rect 54426 59814 54436 59866
rect 54460 59814 54490 59866
rect 54490 59814 54516 59866
rect 54220 59812 54276 59814
rect 54300 59812 54356 59814
rect 54380 59812 54436 59814
rect 54460 59812 54516 59814
rect 54220 58778 54276 58780
rect 54300 58778 54356 58780
rect 54380 58778 54436 58780
rect 54460 58778 54516 58780
rect 54220 58726 54246 58778
rect 54246 58726 54276 58778
rect 54300 58726 54310 58778
rect 54310 58726 54356 58778
rect 54380 58726 54426 58778
rect 54426 58726 54436 58778
rect 54460 58726 54490 58778
rect 54490 58726 54516 58778
rect 54220 58724 54276 58726
rect 54300 58724 54356 58726
rect 54380 58724 54436 58726
rect 54460 58724 54516 58726
rect 54220 57690 54276 57692
rect 54300 57690 54356 57692
rect 54380 57690 54436 57692
rect 54460 57690 54516 57692
rect 54220 57638 54246 57690
rect 54246 57638 54276 57690
rect 54300 57638 54310 57690
rect 54310 57638 54356 57690
rect 54380 57638 54426 57690
rect 54426 57638 54436 57690
rect 54460 57638 54490 57690
rect 54490 57638 54516 57690
rect 54220 57636 54276 57638
rect 54300 57636 54356 57638
rect 54380 57636 54436 57638
rect 54460 57636 54516 57638
rect 54220 56602 54276 56604
rect 54300 56602 54356 56604
rect 54380 56602 54436 56604
rect 54460 56602 54516 56604
rect 54220 56550 54246 56602
rect 54246 56550 54276 56602
rect 54300 56550 54310 56602
rect 54310 56550 54356 56602
rect 54380 56550 54426 56602
rect 54426 56550 54436 56602
rect 54460 56550 54490 56602
rect 54490 56550 54516 56602
rect 54220 56548 54276 56550
rect 54300 56548 54356 56550
rect 54380 56548 54436 56550
rect 54460 56548 54516 56550
rect 54220 55514 54276 55516
rect 54300 55514 54356 55516
rect 54380 55514 54436 55516
rect 54460 55514 54516 55516
rect 54220 55462 54246 55514
rect 54246 55462 54276 55514
rect 54300 55462 54310 55514
rect 54310 55462 54356 55514
rect 54380 55462 54426 55514
rect 54426 55462 54436 55514
rect 54460 55462 54490 55514
rect 54490 55462 54516 55514
rect 54220 55460 54276 55462
rect 54300 55460 54356 55462
rect 54380 55460 54436 55462
rect 54460 55460 54516 55462
rect 54220 54426 54276 54428
rect 54300 54426 54356 54428
rect 54380 54426 54436 54428
rect 54460 54426 54516 54428
rect 54220 54374 54246 54426
rect 54246 54374 54276 54426
rect 54300 54374 54310 54426
rect 54310 54374 54356 54426
rect 54380 54374 54426 54426
rect 54426 54374 54436 54426
rect 54460 54374 54490 54426
rect 54490 54374 54516 54426
rect 54220 54372 54276 54374
rect 54300 54372 54356 54374
rect 54380 54372 54436 54374
rect 54460 54372 54516 54374
rect 54220 53338 54276 53340
rect 54300 53338 54356 53340
rect 54380 53338 54436 53340
rect 54460 53338 54516 53340
rect 54220 53286 54246 53338
rect 54246 53286 54276 53338
rect 54300 53286 54310 53338
rect 54310 53286 54356 53338
rect 54380 53286 54426 53338
rect 54426 53286 54436 53338
rect 54460 53286 54490 53338
rect 54490 53286 54516 53338
rect 54220 53284 54276 53286
rect 54300 53284 54356 53286
rect 54380 53284 54436 53286
rect 54460 53284 54516 53286
rect 54220 52250 54276 52252
rect 54300 52250 54356 52252
rect 54380 52250 54436 52252
rect 54460 52250 54516 52252
rect 54220 52198 54246 52250
rect 54246 52198 54276 52250
rect 54300 52198 54310 52250
rect 54310 52198 54356 52250
rect 54380 52198 54426 52250
rect 54426 52198 54436 52250
rect 54460 52198 54490 52250
rect 54490 52198 54516 52250
rect 54220 52196 54276 52198
rect 54300 52196 54356 52198
rect 54380 52196 54436 52198
rect 54460 52196 54516 52198
rect 54220 51162 54276 51164
rect 54300 51162 54356 51164
rect 54380 51162 54436 51164
rect 54460 51162 54516 51164
rect 54220 51110 54246 51162
rect 54246 51110 54276 51162
rect 54300 51110 54310 51162
rect 54310 51110 54356 51162
rect 54380 51110 54426 51162
rect 54426 51110 54436 51162
rect 54460 51110 54490 51162
rect 54490 51110 54516 51162
rect 54220 51108 54276 51110
rect 54300 51108 54356 51110
rect 54380 51108 54436 51110
rect 54460 51108 54516 51110
rect 54220 50074 54276 50076
rect 54300 50074 54356 50076
rect 54380 50074 54436 50076
rect 54460 50074 54516 50076
rect 54220 50022 54246 50074
rect 54246 50022 54276 50074
rect 54300 50022 54310 50074
rect 54310 50022 54356 50074
rect 54380 50022 54426 50074
rect 54426 50022 54436 50074
rect 54460 50022 54490 50074
rect 54490 50022 54516 50074
rect 54220 50020 54276 50022
rect 54300 50020 54356 50022
rect 54380 50020 54436 50022
rect 54460 50020 54516 50022
rect 54220 48986 54276 48988
rect 54300 48986 54356 48988
rect 54380 48986 54436 48988
rect 54460 48986 54516 48988
rect 54220 48934 54246 48986
rect 54246 48934 54276 48986
rect 54300 48934 54310 48986
rect 54310 48934 54356 48986
rect 54380 48934 54426 48986
rect 54426 48934 54436 48986
rect 54460 48934 54490 48986
rect 54490 48934 54516 48986
rect 54220 48932 54276 48934
rect 54300 48932 54356 48934
rect 54380 48932 54436 48934
rect 54460 48932 54516 48934
rect 54220 47898 54276 47900
rect 54300 47898 54356 47900
rect 54380 47898 54436 47900
rect 54460 47898 54516 47900
rect 54220 47846 54246 47898
rect 54246 47846 54276 47898
rect 54300 47846 54310 47898
rect 54310 47846 54356 47898
rect 54380 47846 54426 47898
rect 54426 47846 54436 47898
rect 54460 47846 54490 47898
rect 54490 47846 54516 47898
rect 54220 47844 54276 47846
rect 54300 47844 54356 47846
rect 54380 47844 54436 47846
rect 54460 47844 54516 47846
rect 54220 46810 54276 46812
rect 54300 46810 54356 46812
rect 54380 46810 54436 46812
rect 54460 46810 54516 46812
rect 54220 46758 54246 46810
rect 54246 46758 54276 46810
rect 54300 46758 54310 46810
rect 54310 46758 54356 46810
rect 54380 46758 54426 46810
rect 54426 46758 54436 46810
rect 54460 46758 54490 46810
rect 54490 46758 54516 46810
rect 54220 46756 54276 46758
rect 54300 46756 54356 46758
rect 54380 46756 54436 46758
rect 54460 46756 54516 46758
rect 54220 45722 54276 45724
rect 54300 45722 54356 45724
rect 54380 45722 54436 45724
rect 54460 45722 54516 45724
rect 54220 45670 54246 45722
rect 54246 45670 54276 45722
rect 54300 45670 54310 45722
rect 54310 45670 54356 45722
rect 54380 45670 54426 45722
rect 54426 45670 54436 45722
rect 54460 45670 54490 45722
rect 54490 45670 54516 45722
rect 54220 45668 54276 45670
rect 54300 45668 54356 45670
rect 54380 45668 54436 45670
rect 54460 45668 54516 45670
rect 54220 44634 54276 44636
rect 54300 44634 54356 44636
rect 54380 44634 54436 44636
rect 54460 44634 54516 44636
rect 54220 44582 54246 44634
rect 54246 44582 54276 44634
rect 54300 44582 54310 44634
rect 54310 44582 54356 44634
rect 54380 44582 54426 44634
rect 54426 44582 54436 44634
rect 54460 44582 54490 44634
rect 54490 44582 54516 44634
rect 54220 44580 54276 44582
rect 54300 44580 54356 44582
rect 54380 44580 54436 44582
rect 54460 44580 54516 44582
rect 54220 43546 54276 43548
rect 54300 43546 54356 43548
rect 54380 43546 54436 43548
rect 54460 43546 54516 43548
rect 54220 43494 54246 43546
rect 54246 43494 54276 43546
rect 54300 43494 54310 43546
rect 54310 43494 54356 43546
rect 54380 43494 54426 43546
rect 54426 43494 54436 43546
rect 54460 43494 54490 43546
rect 54490 43494 54516 43546
rect 54220 43492 54276 43494
rect 54300 43492 54356 43494
rect 54380 43492 54436 43494
rect 54460 43492 54516 43494
rect 54220 42458 54276 42460
rect 54300 42458 54356 42460
rect 54380 42458 54436 42460
rect 54460 42458 54516 42460
rect 54220 42406 54246 42458
rect 54246 42406 54276 42458
rect 54300 42406 54310 42458
rect 54310 42406 54356 42458
rect 54380 42406 54426 42458
rect 54426 42406 54436 42458
rect 54460 42406 54490 42458
rect 54490 42406 54516 42458
rect 54220 42404 54276 42406
rect 54300 42404 54356 42406
rect 54380 42404 54436 42406
rect 54460 42404 54516 42406
rect 54220 41370 54276 41372
rect 54300 41370 54356 41372
rect 54380 41370 54436 41372
rect 54460 41370 54516 41372
rect 54220 41318 54246 41370
rect 54246 41318 54276 41370
rect 54300 41318 54310 41370
rect 54310 41318 54356 41370
rect 54380 41318 54426 41370
rect 54426 41318 54436 41370
rect 54460 41318 54490 41370
rect 54490 41318 54516 41370
rect 54220 41316 54276 41318
rect 54300 41316 54356 41318
rect 54380 41316 54436 41318
rect 54460 41316 54516 41318
rect 54220 40282 54276 40284
rect 54300 40282 54356 40284
rect 54380 40282 54436 40284
rect 54460 40282 54516 40284
rect 54220 40230 54246 40282
rect 54246 40230 54276 40282
rect 54300 40230 54310 40282
rect 54310 40230 54356 40282
rect 54380 40230 54426 40282
rect 54426 40230 54436 40282
rect 54460 40230 54490 40282
rect 54490 40230 54516 40282
rect 54220 40228 54276 40230
rect 54300 40228 54356 40230
rect 54380 40228 54436 40230
rect 54460 40228 54516 40230
rect 54220 39194 54276 39196
rect 54300 39194 54356 39196
rect 54380 39194 54436 39196
rect 54460 39194 54516 39196
rect 54220 39142 54246 39194
rect 54246 39142 54276 39194
rect 54300 39142 54310 39194
rect 54310 39142 54356 39194
rect 54380 39142 54426 39194
rect 54426 39142 54436 39194
rect 54460 39142 54490 39194
rect 54490 39142 54516 39194
rect 54220 39140 54276 39142
rect 54300 39140 54356 39142
rect 54380 39140 54436 39142
rect 54460 39140 54516 39142
rect 54220 38106 54276 38108
rect 54300 38106 54356 38108
rect 54380 38106 54436 38108
rect 54460 38106 54516 38108
rect 54220 38054 54246 38106
rect 54246 38054 54276 38106
rect 54300 38054 54310 38106
rect 54310 38054 54356 38106
rect 54380 38054 54426 38106
rect 54426 38054 54436 38106
rect 54460 38054 54490 38106
rect 54490 38054 54516 38106
rect 54220 38052 54276 38054
rect 54300 38052 54356 38054
rect 54380 38052 54436 38054
rect 54460 38052 54516 38054
rect 54220 37018 54276 37020
rect 54300 37018 54356 37020
rect 54380 37018 54436 37020
rect 54460 37018 54516 37020
rect 54220 36966 54246 37018
rect 54246 36966 54276 37018
rect 54300 36966 54310 37018
rect 54310 36966 54356 37018
rect 54380 36966 54426 37018
rect 54426 36966 54436 37018
rect 54460 36966 54490 37018
rect 54490 36966 54516 37018
rect 54220 36964 54276 36966
rect 54300 36964 54356 36966
rect 54380 36964 54436 36966
rect 54460 36964 54516 36966
rect 54220 35930 54276 35932
rect 54300 35930 54356 35932
rect 54380 35930 54436 35932
rect 54460 35930 54516 35932
rect 54220 35878 54246 35930
rect 54246 35878 54276 35930
rect 54300 35878 54310 35930
rect 54310 35878 54356 35930
rect 54380 35878 54426 35930
rect 54426 35878 54436 35930
rect 54460 35878 54490 35930
rect 54490 35878 54516 35930
rect 54220 35876 54276 35878
rect 54300 35876 54356 35878
rect 54380 35876 54436 35878
rect 54460 35876 54516 35878
rect 54220 34842 54276 34844
rect 54300 34842 54356 34844
rect 54380 34842 54436 34844
rect 54460 34842 54516 34844
rect 54220 34790 54246 34842
rect 54246 34790 54276 34842
rect 54300 34790 54310 34842
rect 54310 34790 54356 34842
rect 54380 34790 54426 34842
rect 54426 34790 54436 34842
rect 54460 34790 54490 34842
rect 54490 34790 54516 34842
rect 54220 34788 54276 34790
rect 54300 34788 54356 34790
rect 54380 34788 54436 34790
rect 54460 34788 54516 34790
rect 54220 33754 54276 33756
rect 54300 33754 54356 33756
rect 54380 33754 54436 33756
rect 54460 33754 54516 33756
rect 54220 33702 54246 33754
rect 54246 33702 54276 33754
rect 54300 33702 54310 33754
rect 54310 33702 54356 33754
rect 54380 33702 54426 33754
rect 54426 33702 54436 33754
rect 54460 33702 54490 33754
rect 54490 33702 54516 33754
rect 54220 33700 54276 33702
rect 54300 33700 54356 33702
rect 54380 33700 54436 33702
rect 54460 33700 54516 33702
rect 54220 32666 54276 32668
rect 54300 32666 54356 32668
rect 54380 32666 54436 32668
rect 54460 32666 54516 32668
rect 54220 32614 54246 32666
rect 54246 32614 54276 32666
rect 54300 32614 54310 32666
rect 54310 32614 54356 32666
rect 54380 32614 54426 32666
rect 54426 32614 54436 32666
rect 54460 32614 54490 32666
rect 54490 32614 54516 32666
rect 54220 32612 54276 32614
rect 54300 32612 54356 32614
rect 54380 32612 54436 32614
rect 54460 32612 54516 32614
rect 54220 31578 54276 31580
rect 54300 31578 54356 31580
rect 54380 31578 54436 31580
rect 54460 31578 54516 31580
rect 54220 31526 54246 31578
rect 54246 31526 54276 31578
rect 54300 31526 54310 31578
rect 54310 31526 54356 31578
rect 54380 31526 54426 31578
rect 54426 31526 54436 31578
rect 54460 31526 54490 31578
rect 54490 31526 54516 31578
rect 54220 31524 54276 31526
rect 54300 31524 54356 31526
rect 54380 31524 54436 31526
rect 54460 31524 54516 31526
rect 54220 30490 54276 30492
rect 54300 30490 54356 30492
rect 54380 30490 54436 30492
rect 54460 30490 54516 30492
rect 54220 30438 54246 30490
rect 54246 30438 54276 30490
rect 54300 30438 54310 30490
rect 54310 30438 54356 30490
rect 54380 30438 54426 30490
rect 54426 30438 54436 30490
rect 54460 30438 54490 30490
rect 54490 30438 54516 30490
rect 54220 30436 54276 30438
rect 54300 30436 54356 30438
rect 54380 30436 54436 30438
rect 54460 30436 54516 30438
rect 54220 29402 54276 29404
rect 54300 29402 54356 29404
rect 54380 29402 54436 29404
rect 54460 29402 54516 29404
rect 54220 29350 54246 29402
rect 54246 29350 54276 29402
rect 54300 29350 54310 29402
rect 54310 29350 54356 29402
rect 54380 29350 54426 29402
rect 54426 29350 54436 29402
rect 54460 29350 54490 29402
rect 54490 29350 54516 29402
rect 54220 29348 54276 29350
rect 54300 29348 54356 29350
rect 54380 29348 54436 29350
rect 54460 29348 54516 29350
rect 54220 28314 54276 28316
rect 54300 28314 54356 28316
rect 54380 28314 54436 28316
rect 54460 28314 54516 28316
rect 54220 28262 54246 28314
rect 54246 28262 54276 28314
rect 54300 28262 54310 28314
rect 54310 28262 54356 28314
rect 54380 28262 54426 28314
rect 54426 28262 54436 28314
rect 54460 28262 54490 28314
rect 54490 28262 54516 28314
rect 54220 28260 54276 28262
rect 54300 28260 54356 28262
rect 54380 28260 54436 28262
rect 54460 28260 54516 28262
rect 54220 27226 54276 27228
rect 54300 27226 54356 27228
rect 54380 27226 54436 27228
rect 54460 27226 54516 27228
rect 54220 27174 54246 27226
rect 54246 27174 54276 27226
rect 54300 27174 54310 27226
rect 54310 27174 54356 27226
rect 54380 27174 54426 27226
rect 54426 27174 54436 27226
rect 54460 27174 54490 27226
rect 54490 27174 54516 27226
rect 54220 27172 54276 27174
rect 54300 27172 54356 27174
rect 54380 27172 54436 27174
rect 54460 27172 54516 27174
rect 54220 26138 54276 26140
rect 54300 26138 54356 26140
rect 54380 26138 54436 26140
rect 54460 26138 54516 26140
rect 54220 26086 54246 26138
rect 54246 26086 54276 26138
rect 54300 26086 54310 26138
rect 54310 26086 54356 26138
rect 54380 26086 54426 26138
rect 54426 26086 54436 26138
rect 54460 26086 54490 26138
rect 54490 26086 54516 26138
rect 54220 26084 54276 26086
rect 54300 26084 54356 26086
rect 54380 26084 54436 26086
rect 54460 26084 54516 26086
rect 54220 25050 54276 25052
rect 54300 25050 54356 25052
rect 54380 25050 54436 25052
rect 54460 25050 54516 25052
rect 54220 24998 54246 25050
rect 54246 24998 54276 25050
rect 54300 24998 54310 25050
rect 54310 24998 54356 25050
rect 54380 24998 54426 25050
rect 54426 24998 54436 25050
rect 54460 24998 54490 25050
rect 54490 24998 54516 25050
rect 54220 24996 54276 24998
rect 54300 24996 54356 24998
rect 54380 24996 54436 24998
rect 54460 24996 54516 24998
rect 54220 23962 54276 23964
rect 54300 23962 54356 23964
rect 54380 23962 54436 23964
rect 54460 23962 54516 23964
rect 54220 23910 54246 23962
rect 54246 23910 54276 23962
rect 54300 23910 54310 23962
rect 54310 23910 54356 23962
rect 54380 23910 54426 23962
rect 54426 23910 54436 23962
rect 54460 23910 54490 23962
rect 54490 23910 54516 23962
rect 54220 23908 54276 23910
rect 54300 23908 54356 23910
rect 54380 23908 54436 23910
rect 54460 23908 54516 23910
rect 52274 2488 52330 2544
rect 54220 22874 54276 22876
rect 54300 22874 54356 22876
rect 54380 22874 54436 22876
rect 54460 22874 54516 22876
rect 54220 22822 54246 22874
rect 54246 22822 54276 22874
rect 54300 22822 54310 22874
rect 54310 22822 54356 22874
rect 54380 22822 54426 22874
rect 54426 22822 54436 22874
rect 54460 22822 54490 22874
rect 54490 22822 54516 22874
rect 54220 22820 54276 22822
rect 54300 22820 54356 22822
rect 54380 22820 54436 22822
rect 54460 22820 54516 22822
rect 54220 21786 54276 21788
rect 54300 21786 54356 21788
rect 54380 21786 54436 21788
rect 54460 21786 54516 21788
rect 54220 21734 54246 21786
rect 54246 21734 54276 21786
rect 54300 21734 54310 21786
rect 54310 21734 54356 21786
rect 54380 21734 54426 21786
rect 54426 21734 54436 21786
rect 54460 21734 54490 21786
rect 54490 21734 54516 21786
rect 54220 21732 54276 21734
rect 54300 21732 54356 21734
rect 54380 21732 54436 21734
rect 54460 21732 54516 21734
rect 54220 20698 54276 20700
rect 54300 20698 54356 20700
rect 54380 20698 54436 20700
rect 54460 20698 54516 20700
rect 54220 20646 54246 20698
rect 54246 20646 54276 20698
rect 54300 20646 54310 20698
rect 54310 20646 54356 20698
rect 54380 20646 54426 20698
rect 54426 20646 54436 20698
rect 54460 20646 54490 20698
rect 54490 20646 54516 20698
rect 54220 20644 54276 20646
rect 54300 20644 54356 20646
rect 54380 20644 54436 20646
rect 54460 20644 54516 20646
rect 54220 19610 54276 19612
rect 54300 19610 54356 19612
rect 54380 19610 54436 19612
rect 54460 19610 54516 19612
rect 54220 19558 54246 19610
rect 54246 19558 54276 19610
rect 54300 19558 54310 19610
rect 54310 19558 54356 19610
rect 54380 19558 54426 19610
rect 54426 19558 54436 19610
rect 54460 19558 54490 19610
rect 54490 19558 54516 19610
rect 54220 19556 54276 19558
rect 54300 19556 54356 19558
rect 54380 19556 54436 19558
rect 54460 19556 54516 19558
rect 54220 18522 54276 18524
rect 54300 18522 54356 18524
rect 54380 18522 54436 18524
rect 54460 18522 54516 18524
rect 54220 18470 54246 18522
rect 54246 18470 54276 18522
rect 54300 18470 54310 18522
rect 54310 18470 54356 18522
rect 54380 18470 54426 18522
rect 54426 18470 54436 18522
rect 54460 18470 54490 18522
rect 54490 18470 54516 18522
rect 54220 18468 54276 18470
rect 54300 18468 54356 18470
rect 54380 18468 54436 18470
rect 54460 18468 54516 18470
rect 54220 17434 54276 17436
rect 54300 17434 54356 17436
rect 54380 17434 54436 17436
rect 54460 17434 54516 17436
rect 54220 17382 54246 17434
rect 54246 17382 54276 17434
rect 54300 17382 54310 17434
rect 54310 17382 54356 17434
rect 54380 17382 54426 17434
rect 54426 17382 54436 17434
rect 54460 17382 54490 17434
rect 54490 17382 54516 17434
rect 54220 17380 54276 17382
rect 54300 17380 54356 17382
rect 54380 17380 54436 17382
rect 54460 17380 54516 17382
rect 54220 16346 54276 16348
rect 54300 16346 54356 16348
rect 54380 16346 54436 16348
rect 54460 16346 54516 16348
rect 54220 16294 54246 16346
rect 54246 16294 54276 16346
rect 54300 16294 54310 16346
rect 54310 16294 54356 16346
rect 54380 16294 54426 16346
rect 54426 16294 54436 16346
rect 54460 16294 54490 16346
rect 54490 16294 54516 16346
rect 54220 16292 54276 16294
rect 54300 16292 54356 16294
rect 54380 16292 54436 16294
rect 54460 16292 54516 16294
rect 54220 15258 54276 15260
rect 54300 15258 54356 15260
rect 54380 15258 54436 15260
rect 54460 15258 54516 15260
rect 54220 15206 54246 15258
rect 54246 15206 54276 15258
rect 54300 15206 54310 15258
rect 54310 15206 54356 15258
rect 54380 15206 54426 15258
rect 54426 15206 54436 15258
rect 54460 15206 54490 15258
rect 54490 15206 54516 15258
rect 54220 15204 54276 15206
rect 54300 15204 54356 15206
rect 54380 15204 54436 15206
rect 54460 15204 54516 15206
rect 54220 14170 54276 14172
rect 54300 14170 54356 14172
rect 54380 14170 54436 14172
rect 54460 14170 54516 14172
rect 54220 14118 54246 14170
rect 54246 14118 54276 14170
rect 54300 14118 54310 14170
rect 54310 14118 54356 14170
rect 54380 14118 54426 14170
rect 54426 14118 54436 14170
rect 54460 14118 54490 14170
rect 54490 14118 54516 14170
rect 54220 14116 54276 14118
rect 54300 14116 54356 14118
rect 54380 14116 54436 14118
rect 54460 14116 54516 14118
rect 54220 13082 54276 13084
rect 54300 13082 54356 13084
rect 54380 13082 54436 13084
rect 54460 13082 54516 13084
rect 54220 13030 54246 13082
rect 54246 13030 54276 13082
rect 54300 13030 54310 13082
rect 54310 13030 54356 13082
rect 54380 13030 54426 13082
rect 54426 13030 54436 13082
rect 54460 13030 54490 13082
rect 54490 13030 54516 13082
rect 54220 13028 54276 13030
rect 54300 13028 54356 13030
rect 54380 13028 54436 13030
rect 54460 13028 54516 13030
rect 54220 11994 54276 11996
rect 54300 11994 54356 11996
rect 54380 11994 54436 11996
rect 54460 11994 54516 11996
rect 54220 11942 54246 11994
rect 54246 11942 54276 11994
rect 54300 11942 54310 11994
rect 54310 11942 54356 11994
rect 54380 11942 54426 11994
rect 54426 11942 54436 11994
rect 54460 11942 54490 11994
rect 54490 11942 54516 11994
rect 54220 11940 54276 11942
rect 54300 11940 54356 11942
rect 54380 11940 54436 11942
rect 54460 11940 54516 11942
rect 54220 10906 54276 10908
rect 54300 10906 54356 10908
rect 54380 10906 54436 10908
rect 54460 10906 54516 10908
rect 54220 10854 54246 10906
rect 54246 10854 54276 10906
rect 54300 10854 54310 10906
rect 54310 10854 54356 10906
rect 54380 10854 54426 10906
rect 54426 10854 54436 10906
rect 54460 10854 54490 10906
rect 54490 10854 54516 10906
rect 54220 10852 54276 10854
rect 54300 10852 54356 10854
rect 54380 10852 54436 10854
rect 54460 10852 54516 10854
rect 54220 9818 54276 9820
rect 54300 9818 54356 9820
rect 54380 9818 54436 9820
rect 54460 9818 54516 9820
rect 54220 9766 54246 9818
rect 54246 9766 54276 9818
rect 54300 9766 54310 9818
rect 54310 9766 54356 9818
rect 54380 9766 54426 9818
rect 54426 9766 54436 9818
rect 54460 9766 54490 9818
rect 54490 9766 54516 9818
rect 54220 9764 54276 9766
rect 54300 9764 54356 9766
rect 54380 9764 54436 9766
rect 54460 9764 54516 9766
rect 53746 4936 53802 4992
rect 54220 8730 54276 8732
rect 54300 8730 54356 8732
rect 54380 8730 54436 8732
rect 54460 8730 54516 8732
rect 54220 8678 54246 8730
rect 54246 8678 54276 8730
rect 54300 8678 54310 8730
rect 54310 8678 54356 8730
rect 54380 8678 54426 8730
rect 54426 8678 54436 8730
rect 54460 8678 54490 8730
rect 54490 8678 54516 8730
rect 54220 8676 54276 8678
rect 54300 8676 54356 8678
rect 54380 8676 54436 8678
rect 54460 8676 54516 8678
rect 54220 7642 54276 7644
rect 54300 7642 54356 7644
rect 54380 7642 54436 7644
rect 54460 7642 54516 7644
rect 54220 7590 54246 7642
rect 54246 7590 54276 7642
rect 54300 7590 54310 7642
rect 54310 7590 54356 7642
rect 54380 7590 54426 7642
rect 54426 7590 54436 7642
rect 54460 7590 54490 7642
rect 54490 7590 54516 7642
rect 54220 7588 54276 7590
rect 54300 7588 54356 7590
rect 54380 7588 54436 7590
rect 54460 7588 54516 7590
rect 54220 6554 54276 6556
rect 54300 6554 54356 6556
rect 54380 6554 54436 6556
rect 54460 6554 54516 6556
rect 54220 6502 54246 6554
rect 54246 6502 54276 6554
rect 54300 6502 54310 6554
rect 54310 6502 54356 6554
rect 54380 6502 54426 6554
rect 54426 6502 54436 6554
rect 54460 6502 54490 6554
rect 54490 6502 54516 6554
rect 54220 6500 54276 6502
rect 54300 6500 54356 6502
rect 54380 6500 54436 6502
rect 54460 6500 54516 6502
rect 54220 5466 54276 5468
rect 54300 5466 54356 5468
rect 54380 5466 54436 5468
rect 54460 5466 54516 5468
rect 54220 5414 54246 5466
rect 54246 5414 54276 5466
rect 54300 5414 54310 5466
rect 54310 5414 54356 5466
rect 54380 5414 54426 5466
rect 54426 5414 54436 5466
rect 54460 5414 54490 5466
rect 54490 5414 54516 5466
rect 54220 5412 54276 5414
rect 54300 5412 54356 5414
rect 54380 5412 54436 5414
rect 54460 5412 54516 5414
rect 54220 4378 54276 4380
rect 54300 4378 54356 4380
rect 54380 4378 54436 4380
rect 54460 4378 54516 4380
rect 54220 4326 54246 4378
rect 54246 4326 54276 4378
rect 54300 4326 54310 4378
rect 54310 4326 54356 4378
rect 54380 4326 54426 4378
rect 54426 4326 54436 4378
rect 54460 4326 54490 4378
rect 54490 4326 54516 4378
rect 54220 4324 54276 4326
rect 54300 4324 54356 4326
rect 54380 4324 54436 4326
rect 54460 4324 54516 4326
rect 54220 3290 54276 3292
rect 54300 3290 54356 3292
rect 54380 3290 54436 3292
rect 54460 3290 54516 3292
rect 54220 3238 54246 3290
rect 54246 3238 54276 3290
rect 54300 3238 54310 3290
rect 54310 3238 54356 3290
rect 54380 3238 54426 3290
rect 54426 3238 54436 3290
rect 54460 3238 54490 3290
rect 54490 3238 54516 3290
rect 54220 3236 54276 3238
rect 54300 3236 54356 3238
rect 54380 3236 54436 3238
rect 54460 3236 54516 3238
rect 54220 2202 54276 2204
rect 54300 2202 54356 2204
rect 54380 2202 54436 2204
rect 54460 2202 54516 2204
rect 54220 2150 54246 2202
rect 54246 2150 54276 2202
rect 54300 2150 54310 2202
rect 54310 2150 54356 2202
rect 54380 2150 54426 2202
rect 54426 2150 54436 2202
rect 54460 2150 54490 2202
rect 54490 2150 54516 2202
rect 54220 2148 54276 2150
rect 54300 2148 54356 2150
rect 54380 2148 54436 2150
rect 54460 2148 54516 2150
rect 54390 1944 54446 2000
rect 59220 66938 59276 66940
rect 59300 66938 59356 66940
rect 59380 66938 59436 66940
rect 59460 66938 59516 66940
rect 59220 66886 59246 66938
rect 59246 66886 59276 66938
rect 59300 66886 59310 66938
rect 59310 66886 59356 66938
rect 59380 66886 59426 66938
rect 59426 66886 59436 66938
rect 59460 66886 59490 66938
rect 59490 66886 59516 66938
rect 59220 66884 59276 66886
rect 59300 66884 59356 66886
rect 59380 66884 59436 66886
rect 59460 66884 59516 66886
rect 64220 66394 64276 66396
rect 64300 66394 64356 66396
rect 64380 66394 64436 66396
rect 64460 66394 64516 66396
rect 64220 66342 64246 66394
rect 64246 66342 64276 66394
rect 64300 66342 64310 66394
rect 64310 66342 64356 66394
rect 64380 66342 64426 66394
rect 64426 66342 64436 66394
rect 64460 66342 64490 66394
rect 64490 66342 64516 66394
rect 64220 66340 64276 66342
rect 64300 66340 64356 66342
rect 64380 66340 64436 66342
rect 64460 66340 64516 66342
rect 59220 65850 59276 65852
rect 59300 65850 59356 65852
rect 59380 65850 59436 65852
rect 59460 65850 59516 65852
rect 59220 65798 59246 65850
rect 59246 65798 59276 65850
rect 59300 65798 59310 65850
rect 59310 65798 59356 65850
rect 59380 65798 59426 65850
rect 59426 65798 59436 65850
rect 59460 65798 59490 65850
rect 59490 65798 59516 65850
rect 59220 65796 59276 65798
rect 59300 65796 59356 65798
rect 59380 65796 59436 65798
rect 59460 65796 59516 65798
rect 54942 4936 54998 4992
rect 55954 5208 56010 5264
rect 55954 3712 56010 3768
rect 59220 64762 59276 64764
rect 59300 64762 59356 64764
rect 59380 64762 59436 64764
rect 59460 64762 59516 64764
rect 59220 64710 59246 64762
rect 59246 64710 59276 64762
rect 59300 64710 59310 64762
rect 59310 64710 59356 64762
rect 59380 64710 59426 64762
rect 59426 64710 59436 64762
rect 59460 64710 59490 64762
rect 59490 64710 59516 64762
rect 59220 64708 59276 64710
rect 59300 64708 59356 64710
rect 59380 64708 59436 64710
rect 59460 64708 59516 64710
rect 59220 63674 59276 63676
rect 59300 63674 59356 63676
rect 59380 63674 59436 63676
rect 59460 63674 59516 63676
rect 59220 63622 59246 63674
rect 59246 63622 59276 63674
rect 59300 63622 59310 63674
rect 59310 63622 59356 63674
rect 59380 63622 59426 63674
rect 59426 63622 59436 63674
rect 59460 63622 59490 63674
rect 59490 63622 59516 63674
rect 59220 63620 59276 63622
rect 59300 63620 59356 63622
rect 59380 63620 59436 63622
rect 59460 63620 59516 63622
rect 59220 62586 59276 62588
rect 59300 62586 59356 62588
rect 59380 62586 59436 62588
rect 59460 62586 59516 62588
rect 59220 62534 59246 62586
rect 59246 62534 59276 62586
rect 59300 62534 59310 62586
rect 59310 62534 59356 62586
rect 59380 62534 59426 62586
rect 59426 62534 59436 62586
rect 59460 62534 59490 62586
rect 59490 62534 59516 62586
rect 59220 62532 59276 62534
rect 59300 62532 59356 62534
rect 59380 62532 59436 62534
rect 59460 62532 59516 62534
rect 59220 61498 59276 61500
rect 59300 61498 59356 61500
rect 59380 61498 59436 61500
rect 59460 61498 59516 61500
rect 59220 61446 59246 61498
rect 59246 61446 59276 61498
rect 59300 61446 59310 61498
rect 59310 61446 59356 61498
rect 59380 61446 59426 61498
rect 59426 61446 59436 61498
rect 59460 61446 59490 61498
rect 59490 61446 59516 61498
rect 59220 61444 59276 61446
rect 59300 61444 59356 61446
rect 59380 61444 59436 61446
rect 59460 61444 59516 61446
rect 59220 60410 59276 60412
rect 59300 60410 59356 60412
rect 59380 60410 59436 60412
rect 59460 60410 59516 60412
rect 59220 60358 59246 60410
rect 59246 60358 59276 60410
rect 59300 60358 59310 60410
rect 59310 60358 59356 60410
rect 59380 60358 59426 60410
rect 59426 60358 59436 60410
rect 59460 60358 59490 60410
rect 59490 60358 59516 60410
rect 59220 60356 59276 60358
rect 59300 60356 59356 60358
rect 59380 60356 59436 60358
rect 59460 60356 59516 60358
rect 59220 59322 59276 59324
rect 59300 59322 59356 59324
rect 59380 59322 59436 59324
rect 59460 59322 59516 59324
rect 59220 59270 59246 59322
rect 59246 59270 59276 59322
rect 59300 59270 59310 59322
rect 59310 59270 59356 59322
rect 59380 59270 59426 59322
rect 59426 59270 59436 59322
rect 59460 59270 59490 59322
rect 59490 59270 59516 59322
rect 59220 59268 59276 59270
rect 59300 59268 59356 59270
rect 59380 59268 59436 59270
rect 59460 59268 59516 59270
rect 59220 58234 59276 58236
rect 59300 58234 59356 58236
rect 59380 58234 59436 58236
rect 59460 58234 59516 58236
rect 59220 58182 59246 58234
rect 59246 58182 59276 58234
rect 59300 58182 59310 58234
rect 59310 58182 59356 58234
rect 59380 58182 59426 58234
rect 59426 58182 59436 58234
rect 59460 58182 59490 58234
rect 59490 58182 59516 58234
rect 59220 58180 59276 58182
rect 59300 58180 59356 58182
rect 59380 58180 59436 58182
rect 59460 58180 59516 58182
rect 59220 57146 59276 57148
rect 59300 57146 59356 57148
rect 59380 57146 59436 57148
rect 59460 57146 59516 57148
rect 59220 57094 59246 57146
rect 59246 57094 59276 57146
rect 59300 57094 59310 57146
rect 59310 57094 59356 57146
rect 59380 57094 59426 57146
rect 59426 57094 59436 57146
rect 59460 57094 59490 57146
rect 59490 57094 59516 57146
rect 59220 57092 59276 57094
rect 59300 57092 59356 57094
rect 59380 57092 59436 57094
rect 59460 57092 59516 57094
rect 59220 56058 59276 56060
rect 59300 56058 59356 56060
rect 59380 56058 59436 56060
rect 59460 56058 59516 56060
rect 59220 56006 59246 56058
rect 59246 56006 59276 56058
rect 59300 56006 59310 56058
rect 59310 56006 59356 56058
rect 59380 56006 59426 56058
rect 59426 56006 59436 56058
rect 59460 56006 59490 56058
rect 59490 56006 59516 56058
rect 59220 56004 59276 56006
rect 59300 56004 59356 56006
rect 59380 56004 59436 56006
rect 59460 56004 59516 56006
rect 59220 54970 59276 54972
rect 59300 54970 59356 54972
rect 59380 54970 59436 54972
rect 59460 54970 59516 54972
rect 59220 54918 59246 54970
rect 59246 54918 59276 54970
rect 59300 54918 59310 54970
rect 59310 54918 59356 54970
rect 59380 54918 59426 54970
rect 59426 54918 59436 54970
rect 59460 54918 59490 54970
rect 59490 54918 59516 54970
rect 59220 54916 59276 54918
rect 59300 54916 59356 54918
rect 59380 54916 59436 54918
rect 59460 54916 59516 54918
rect 59220 53882 59276 53884
rect 59300 53882 59356 53884
rect 59380 53882 59436 53884
rect 59460 53882 59516 53884
rect 59220 53830 59246 53882
rect 59246 53830 59276 53882
rect 59300 53830 59310 53882
rect 59310 53830 59356 53882
rect 59380 53830 59426 53882
rect 59426 53830 59436 53882
rect 59460 53830 59490 53882
rect 59490 53830 59516 53882
rect 59220 53828 59276 53830
rect 59300 53828 59356 53830
rect 59380 53828 59436 53830
rect 59460 53828 59516 53830
rect 59220 52794 59276 52796
rect 59300 52794 59356 52796
rect 59380 52794 59436 52796
rect 59460 52794 59516 52796
rect 59220 52742 59246 52794
rect 59246 52742 59276 52794
rect 59300 52742 59310 52794
rect 59310 52742 59356 52794
rect 59380 52742 59426 52794
rect 59426 52742 59436 52794
rect 59460 52742 59490 52794
rect 59490 52742 59516 52794
rect 59220 52740 59276 52742
rect 59300 52740 59356 52742
rect 59380 52740 59436 52742
rect 59460 52740 59516 52742
rect 59220 51706 59276 51708
rect 59300 51706 59356 51708
rect 59380 51706 59436 51708
rect 59460 51706 59516 51708
rect 59220 51654 59246 51706
rect 59246 51654 59276 51706
rect 59300 51654 59310 51706
rect 59310 51654 59356 51706
rect 59380 51654 59426 51706
rect 59426 51654 59436 51706
rect 59460 51654 59490 51706
rect 59490 51654 59516 51706
rect 59220 51652 59276 51654
rect 59300 51652 59356 51654
rect 59380 51652 59436 51654
rect 59460 51652 59516 51654
rect 59220 50618 59276 50620
rect 59300 50618 59356 50620
rect 59380 50618 59436 50620
rect 59460 50618 59516 50620
rect 59220 50566 59246 50618
rect 59246 50566 59276 50618
rect 59300 50566 59310 50618
rect 59310 50566 59356 50618
rect 59380 50566 59426 50618
rect 59426 50566 59436 50618
rect 59460 50566 59490 50618
rect 59490 50566 59516 50618
rect 59220 50564 59276 50566
rect 59300 50564 59356 50566
rect 59380 50564 59436 50566
rect 59460 50564 59516 50566
rect 59220 49530 59276 49532
rect 59300 49530 59356 49532
rect 59380 49530 59436 49532
rect 59460 49530 59516 49532
rect 59220 49478 59246 49530
rect 59246 49478 59276 49530
rect 59300 49478 59310 49530
rect 59310 49478 59356 49530
rect 59380 49478 59426 49530
rect 59426 49478 59436 49530
rect 59460 49478 59490 49530
rect 59490 49478 59516 49530
rect 59220 49476 59276 49478
rect 59300 49476 59356 49478
rect 59380 49476 59436 49478
rect 59460 49476 59516 49478
rect 59220 48442 59276 48444
rect 59300 48442 59356 48444
rect 59380 48442 59436 48444
rect 59460 48442 59516 48444
rect 59220 48390 59246 48442
rect 59246 48390 59276 48442
rect 59300 48390 59310 48442
rect 59310 48390 59356 48442
rect 59380 48390 59426 48442
rect 59426 48390 59436 48442
rect 59460 48390 59490 48442
rect 59490 48390 59516 48442
rect 59220 48388 59276 48390
rect 59300 48388 59356 48390
rect 59380 48388 59436 48390
rect 59460 48388 59516 48390
rect 59220 47354 59276 47356
rect 59300 47354 59356 47356
rect 59380 47354 59436 47356
rect 59460 47354 59516 47356
rect 59220 47302 59246 47354
rect 59246 47302 59276 47354
rect 59300 47302 59310 47354
rect 59310 47302 59356 47354
rect 59380 47302 59426 47354
rect 59426 47302 59436 47354
rect 59460 47302 59490 47354
rect 59490 47302 59516 47354
rect 59220 47300 59276 47302
rect 59300 47300 59356 47302
rect 59380 47300 59436 47302
rect 59460 47300 59516 47302
rect 59220 46266 59276 46268
rect 59300 46266 59356 46268
rect 59380 46266 59436 46268
rect 59460 46266 59516 46268
rect 59220 46214 59246 46266
rect 59246 46214 59276 46266
rect 59300 46214 59310 46266
rect 59310 46214 59356 46266
rect 59380 46214 59426 46266
rect 59426 46214 59436 46266
rect 59460 46214 59490 46266
rect 59490 46214 59516 46266
rect 59220 46212 59276 46214
rect 59300 46212 59356 46214
rect 59380 46212 59436 46214
rect 59460 46212 59516 46214
rect 59220 45178 59276 45180
rect 59300 45178 59356 45180
rect 59380 45178 59436 45180
rect 59460 45178 59516 45180
rect 59220 45126 59246 45178
rect 59246 45126 59276 45178
rect 59300 45126 59310 45178
rect 59310 45126 59356 45178
rect 59380 45126 59426 45178
rect 59426 45126 59436 45178
rect 59460 45126 59490 45178
rect 59490 45126 59516 45178
rect 59220 45124 59276 45126
rect 59300 45124 59356 45126
rect 59380 45124 59436 45126
rect 59460 45124 59516 45126
rect 59220 44090 59276 44092
rect 59300 44090 59356 44092
rect 59380 44090 59436 44092
rect 59460 44090 59516 44092
rect 59220 44038 59246 44090
rect 59246 44038 59276 44090
rect 59300 44038 59310 44090
rect 59310 44038 59356 44090
rect 59380 44038 59426 44090
rect 59426 44038 59436 44090
rect 59460 44038 59490 44090
rect 59490 44038 59516 44090
rect 59220 44036 59276 44038
rect 59300 44036 59356 44038
rect 59380 44036 59436 44038
rect 59460 44036 59516 44038
rect 59220 43002 59276 43004
rect 59300 43002 59356 43004
rect 59380 43002 59436 43004
rect 59460 43002 59516 43004
rect 59220 42950 59246 43002
rect 59246 42950 59276 43002
rect 59300 42950 59310 43002
rect 59310 42950 59356 43002
rect 59380 42950 59426 43002
rect 59426 42950 59436 43002
rect 59460 42950 59490 43002
rect 59490 42950 59516 43002
rect 59220 42948 59276 42950
rect 59300 42948 59356 42950
rect 59380 42948 59436 42950
rect 59460 42948 59516 42950
rect 59220 41914 59276 41916
rect 59300 41914 59356 41916
rect 59380 41914 59436 41916
rect 59460 41914 59516 41916
rect 59220 41862 59246 41914
rect 59246 41862 59276 41914
rect 59300 41862 59310 41914
rect 59310 41862 59356 41914
rect 59380 41862 59426 41914
rect 59426 41862 59436 41914
rect 59460 41862 59490 41914
rect 59490 41862 59516 41914
rect 59220 41860 59276 41862
rect 59300 41860 59356 41862
rect 59380 41860 59436 41862
rect 59460 41860 59516 41862
rect 59220 40826 59276 40828
rect 59300 40826 59356 40828
rect 59380 40826 59436 40828
rect 59460 40826 59516 40828
rect 59220 40774 59246 40826
rect 59246 40774 59276 40826
rect 59300 40774 59310 40826
rect 59310 40774 59356 40826
rect 59380 40774 59426 40826
rect 59426 40774 59436 40826
rect 59460 40774 59490 40826
rect 59490 40774 59516 40826
rect 59220 40772 59276 40774
rect 59300 40772 59356 40774
rect 59380 40772 59436 40774
rect 59460 40772 59516 40774
rect 59220 39738 59276 39740
rect 59300 39738 59356 39740
rect 59380 39738 59436 39740
rect 59460 39738 59516 39740
rect 59220 39686 59246 39738
rect 59246 39686 59276 39738
rect 59300 39686 59310 39738
rect 59310 39686 59356 39738
rect 59380 39686 59426 39738
rect 59426 39686 59436 39738
rect 59460 39686 59490 39738
rect 59490 39686 59516 39738
rect 59220 39684 59276 39686
rect 59300 39684 59356 39686
rect 59380 39684 59436 39686
rect 59460 39684 59516 39686
rect 59220 38650 59276 38652
rect 59300 38650 59356 38652
rect 59380 38650 59436 38652
rect 59460 38650 59516 38652
rect 59220 38598 59246 38650
rect 59246 38598 59276 38650
rect 59300 38598 59310 38650
rect 59310 38598 59356 38650
rect 59380 38598 59426 38650
rect 59426 38598 59436 38650
rect 59460 38598 59490 38650
rect 59490 38598 59516 38650
rect 59220 38596 59276 38598
rect 59300 38596 59356 38598
rect 59380 38596 59436 38598
rect 59460 38596 59516 38598
rect 59220 37562 59276 37564
rect 59300 37562 59356 37564
rect 59380 37562 59436 37564
rect 59460 37562 59516 37564
rect 59220 37510 59246 37562
rect 59246 37510 59276 37562
rect 59300 37510 59310 37562
rect 59310 37510 59356 37562
rect 59380 37510 59426 37562
rect 59426 37510 59436 37562
rect 59460 37510 59490 37562
rect 59490 37510 59516 37562
rect 59220 37508 59276 37510
rect 59300 37508 59356 37510
rect 59380 37508 59436 37510
rect 59460 37508 59516 37510
rect 59220 36474 59276 36476
rect 59300 36474 59356 36476
rect 59380 36474 59436 36476
rect 59460 36474 59516 36476
rect 59220 36422 59246 36474
rect 59246 36422 59276 36474
rect 59300 36422 59310 36474
rect 59310 36422 59356 36474
rect 59380 36422 59426 36474
rect 59426 36422 59436 36474
rect 59460 36422 59490 36474
rect 59490 36422 59516 36474
rect 59220 36420 59276 36422
rect 59300 36420 59356 36422
rect 59380 36420 59436 36422
rect 59460 36420 59516 36422
rect 59220 35386 59276 35388
rect 59300 35386 59356 35388
rect 59380 35386 59436 35388
rect 59460 35386 59516 35388
rect 59220 35334 59246 35386
rect 59246 35334 59276 35386
rect 59300 35334 59310 35386
rect 59310 35334 59356 35386
rect 59380 35334 59426 35386
rect 59426 35334 59436 35386
rect 59460 35334 59490 35386
rect 59490 35334 59516 35386
rect 59220 35332 59276 35334
rect 59300 35332 59356 35334
rect 59380 35332 59436 35334
rect 59460 35332 59516 35334
rect 59220 34298 59276 34300
rect 59300 34298 59356 34300
rect 59380 34298 59436 34300
rect 59460 34298 59516 34300
rect 59220 34246 59246 34298
rect 59246 34246 59276 34298
rect 59300 34246 59310 34298
rect 59310 34246 59356 34298
rect 59380 34246 59426 34298
rect 59426 34246 59436 34298
rect 59460 34246 59490 34298
rect 59490 34246 59516 34298
rect 59220 34244 59276 34246
rect 59300 34244 59356 34246
rect 59380 34244 59436 34246
rect 59460 34244 59516 34246
rect 59220 33210 59276 33212
rect 59300 33210 59356 33212
rect 59380 33210 59436 33212
rect 59460 33210 59516 33212
rect 59220 33158 59246 33210
rect 59246 33158 59276 33210
rect 59300 33158 59310 33210
rect 59310 33158 59356 33210
rect 59380 33158 59426 33210
rect 59426 33158 59436 33210
rect 59460 33158 59490 33210
rect 59490 33158 59516 33210
rect 59220 33156 59276 33158
rect 59300 33156 59356 33158
rect 59380 33156 59436 33158
rect 59460 33156 59516 33158
rect 59220 32122 59276 32124
rect 59300 32122 59356 32124
rect 59380 32122 59436 32124
rect 59460 32122 59516 32124
rect 59220 32070 59246 32122
rect 59246 32070 59276 32122
rect 59300 32070 59310 32122
rect 59310 32070 59356 32122
rect 59380 32070 59426 32122
rect 59426 32070 59436 32122
rect 59460 32070 59490 32122
rect 59490 32070 59516 32122
rect 59220 32068 59276 32070
rect 59300 32068 59356 32070
rect 59380 32068 59436 32070
rect 59460 32068 59516 32070
rect 59220 31034 59276 31036
rect 59300 31034 59356 31036
rect 59380 31034 59436 31036
rect 59460 31034 59516 31036
rect 59220 30982 59246 31034
rect 59246 30982 59276 31034
rect 59300 30982 59310 31034
rect 59310 30982 59356 31034
rect 59380 30982 59426 31034
rect 59426 30982 59436 31034
rect 59460 30982 59490 31034
rect 59490 30982 59516 31034
rect 59220 30980 59276 30982
rect 59300 30980 59356 30982
rect 59380 30980 59436 30982
rect 59460 30980 59516 30982
rect 59220 29946 59276 29948
rect 59300 29946 59356 29948
rect 59380 29946 59436 29948
rect 59460 29946 59516 29948
rect 59220 29894 59246 29946
rect 59246 29894 59276 29946
rect 59300 29894 59310 29946
rect 59310 29894 59356 29946
rect 59380 29894 59426 29946
rect 59426 29894 59436 29946
rect 59460 29894 59490 29946
rect 59490 29894 59516 29946
rect 59220 29892 59276 29894
rect 59300 29892 59356 29894
rect 59380 29892 59436 29894
rect 59460 29892 59516 29894
rect 59220 28858 59276 28860
rect 59300 28858 59356 28860
rect 59380 28858 59436 28860
rect 59460 28858 59516 28860
rect 59220 28806 59246 28858
rect 59246 28806 59276 28858
rect 59300 28806 59310 28858
rect 59310 28806 59356 28858
rect 59380 28806 59426 28858
rect 59426 28806 59436 28858
rect 59460 28806 59490 28858
rect 59490 28806 59516 28858
rect 59220 28804 59276 28806
rect 59300 28804 59356 28806
rect 59380 28804 59436 28806
rect 59460 28804 59516 28806
rect 59220 27770 59276 27772
rect 59300 27770 59356 27772
rect 59380 27770 59436 27772
rect 59460 27770 59516 27772
rect 59220 27718 59246 27770
rect 59246 27718 59276 27770
rect 59300 27718 59310 27770
rect 59310 27718 59356 27770
rect 59380 27718 59426 27770
rect 59426 27718 59436 27770
rect 59460 27718 59490 27770
rect 59490 27718 59516 27770
rect 59220 27716 59276 27718
rect 59300 27716 59356 27718
rect 59380 27716 59436 27718
rect 59460 27716 59516 27718
rect 59220 26682 59276 26684
rect 59300 26682 59356 26684
rect 59380 26682 59436 26684
rect 59460 26682 59516 26684
rect 59220 26630 59246 26682
rect 59246 26630 59276 26682
rect 59300 26630 59310 26682
rect 59310 26630 59356 26682
rect 59380 26630 59426 26682
rect 59426 26630 59436 26682
rect 59460 26630 59490 26682
rect 59490 26630 59516 26682
rect 59220 26628 59276 26630
rect 59300 26628 59356 26630
rect 59380 26628 59436 26630
rect 59460 26628 59516 26630
rect 59220 25594 59276 25596
rect 59300 25594 59356 25596
rect 59380 25594 59436 25596
rect 59460 25594 59516 25596
rect 59220 25542 59246 25594
rect 59246 25542 59276 25594
rect 59300 25542 59310 25594
rect 59310 25542 59356 25594
rect 59380 25542 59426 25594
rect 59426 25542 59436 25594
rect 59460 25542 59490 25594
rect 59490 25542 59516 25594
rect 59220 25540 59276 25542
rect 59300 25540 59356 25542
rect 59380 25540 59436 25542
rect 59460 25540 59516 25542
rect 59220 24506 59276 24508
rect 59300 24506 59356 24508
rect 59380 24506 59436 24508
rect 59460 24506 59516 24508
rect 59220 24454 59246 24506
rect 59246 24454 59276 24506
rect 59300 24454 59310 24506
rect 59310 24454 59356 24506
rect 59380 24454 59426 24506
rect 59426 24454 59436 24506
rect 59460 24454 59490 24506
rect 59490 24454 59516 24506
rect 59220 24452 59276 24454
rect 59300 24452 59356 24454
rect 59380 24452 59436 24454
rect 59460 24452 59516 24454
rect 59220 23418 59276 23420
rect 59300 23418 59356 23420
rect 59380 23418 59436 23420
rect 59460 23418 59516 23420
rect 59220 23366 59246 23418
rect 59246 23366 59276 23418
rect 59300 23366 59310 23418
rect 59310 23366 59356 23418
rect 59380 23366 59426 23418
rect 59426 23366 59436 23418
rect 59460 23366 59490 23418
rect 59490 23366 59516 23418
rect 59220 23364 59276 23366
rect 59300 23364 59356 23366
rect 59380 23364 59436 23366
rect 59460 23364 59516 23366
rect 59220 22330 59276 22332
rect 59300 22330 59356 22332
rect 59380 22330 59436 22332
rect 59460 22330 59516 22332
rect 59220 22278 59246 22330
rect 59246 22278 59276 22330
rect 59300 22278 59310 22330
rect 59310 22278 59356 22330
rect 59380 22278 59426 22330
rect 59426 22278 59436 22330
rect 59460 22278 59490 22330
rect 59490 22278 59516 22330
rect 59220 22276 59276 22278
rect 59300 22276 59356 22278
rect 59380 22276 59436 22278
rect 59460 22276 59516 22278
rect 59220 21242 59276 21244
rect 59300 21242 59356 21244
rect 59380 21242 59436 21244
rect 59460 21242 59516 21244
rect 59220 21190 59246 21242
rect 59246 21190 59276 21242
rect 59300 21190 59310 21242
rect 59310 21190 59356 21242
rect 59380 21190 59426 21242
rect 59426 21190 59436 21242
rect 59460 21190 59490 21242
rect 59490 21190 59516 21242
rect 59220 21188 59276 21190
rect 59300 21188 59356 21190
rect 59380 21188 59436 21190
rect 59460 21188 59516 21190
rect 59220 20154 59276 20156
rect 59300 20154 59356 20156
rect 59380 20154 59436 20156
rect 59460 20154 59516 20156
rect 59220 20102 59246 20154
rect 59246 20102 59276 20154
rect 59300 20102 59310 20154
rect 59310 20102 59356 20154
rect 59380 20102 59426 20154
rect 59426 20102 59436 20154
rect 59460 20102 59490 20154
rect 59490 20102 59516 20154
rect 59220 20100 59276 20102
rect 59300 20100 59356 20102
rect 59380 20100 59436 20102
rect 59460 20100 59516 20102
rect 59220 19066 59276 19068
rect 59300 19066 59356 19068
rect 59380 19066 59436 19068
rect 59460 19066 59516 19068
rect 59220 19014 59246 19066
rect 59246 19014 59276 19066
rect 59300 19014 59310 19066
rect 59310 19014 59356 19066
rect 59380 19014 59426 19066
rect 59426 19014 59436 19066
rect 59460 19014 59490 19066
rect 59490 19014 59516 19066
rect 59220 19012 59276 19014
rect 59300 19012 59356 19014
rect 59380 19012 59436 19014
rect 59460 19012 59516 19014
rect 59220 17978 59276 17980
rect 59300 17978 59356 17980
rect 59380 17978 59436 17980
rect 59460 17978 59516 17980
rect 59220 17926 59246 17978
rect 59246 17926 59276 17978
rect 59300 17926 59310 17978
rect 59310 17926 59356 17978
rect 59380 17926 59426 17978
rect 59426 17926 59436 17978
rect 59460 17926 59490 17978
rect 59490 17926 59516 17978
rect 59220 17924 59276 17926
rect 59300 17924 59356 17926
rect 59380 17924 59436 17926
rect 59460 17924 59516 17926
rect 59220 16890 59276 16892
rect 59300 16890 59356 16892
rect 59380 16890 59436 16892
rect 59460 16890 59516 16892
rect 59220 16838 59246 16890
rect 59246 16838 59276 16890
rect 59300 16838 59310 16890
rect 59310 16838 59356 16890
rect 59380 16838 59426 16890
rect 59426 16838 59436 16890
rect 59460 16838 59490 16890
rect 59490 16838 59516 16890
rect 59220 16836 59276 16838
rect 59300 16836 59356 16838
rect 59380 16836 59436 16838
rect 59460 16836 59516 16838
rect 59220 15802 59276 15804
rect 59300 15802 59356 15804
rect 59380 15802 59436 15804
rect 59460 15802 59516 15804
rect 59220 15750 59246 15802
rect 59246 15750 59276 15802
rect 59300 15750 59310 15802
rect 59310 15750 59356 15802
rect 59380 15750 59426 15802
rect 59426 15750 59436 15802
rect 59460 15750 59490 15802
rect 59490 15750 59516 15802
rect 59220 15748 59276 15750
rect 59300 15748 59356 15750
rect 59380 15748 59436 15750
rect 59460 15748 59516 15750
rect 59220 14714 59276 14716
rect 59300 14714 59356 14716
rect 59380 14714 59436 14716
rect 59460 14714 59516 14716
rect 59220 14662 59246 14714
rect 59246 14662 59276 14714
rect 59300 14662 59310 14714
rect 59310 14662 59356 14714
rect 59380 14662 59426 14714
rect 59426 14662 59436 14714
rect 59460 14662 59490 14714
rect 59490 14662 59516 14714
rect 59220 14660 59276 14662
rect 59300 14660 59356 14662
rect 59380 14660 59436 14662
rect 59460 14660 59516 14662
rect 59220 13626 59276 13628
rect 59300 13626 59356 13628
rect 59380 13626 59436 13628
rect 59460 13626 59516 13628
rect 59220 13574 59246 13626
rect 59246 13574 59276 13626
rect 59300 13574 59310 13626
rect 59310 13574 59356 13626
rect 59380 13574 59426 13626
rect 59426 13574 59436 13626
rect 59460 13574 59490 13626
rect 59490 13574 59516 13626
rect 59220 13572 59276 13574
rect 59300 13572 59356 13574
rect 59380 13572 59436 13574
rect 59460 13572 59516 13574
rect 59220 12538 59276 12540
rect 59300 12538 59356 12540
rect 59380 12538 59436 12540
rect 59460 12538 59516 12540
rect 59220 12486 59246 12538
rect 59246 12486 59276 12538
rect 59300 12486 59310 12538
rect 59310 12486 59356 12538
rect 59380 12486 59426 12538
rect 59426 12486 59436 12538
rect 59460 12486 59490 12538
rect 59490 12486 59516 12538
rect 59220 12484 59276 12486
rect 59300 12484 59356 12486
rect 59380 12484 59436 12486
rect 59460 12484 59516 12486
rect 59220 11450 59276 11452
rect 59300 11450 59356 11452
rect 59380 11450 59436 11452
rect 59460 11450 59516 11452
rect 59220 11398 59246 11450
rect 59246 11398 59276 11450
rect 59300 11398 59310 11450
rect 59310 11398 59356 11450
rect 59380 11398 59426 11450
rect 59426 11398 59436 11450
rect 59460 11398 59490 11450
rect 59490 11398 59516 11450
rect 59220 11396 59276 11398
rect 59300 11396 59356 11398
rect 59380 11396 59436 11398
rect 59460 11396 59516 11398
rect 59220 10362 59276 10364
rect 59300 10362 59356 10364
rect 59380 10362 59436 10364
rect 59460 10362 59516 10364
rect 59220 10310 59246 10362
rect 59246 10310 59276 10362
rect 59300 10310 59310 10362
rect 59310 10310 59356 10362
rect 59380 10310 59426 10362
rect 59426 10310 59436 10362
rect 59460 10310 59490 10362
rect 59490 10310 59516 10362
rect 59220 10308 59276 10310
rect 59300 10308 59356 10310
rect 59380 10308 59436 10310
rect 59460 10308 59516 10310
rect 59220 9274 59276 9276
rect 59300 9274 59356 9276
rect 59380 9274 59436 9276
rect 59460 9274 59516 9276
rect 59220 9222 59246 9274
rect 59246 9222 59276 9274
rect 59300 9222 59310 9274
rect 59310 9222 59356 9274
rect 59380 9222 59426 9274
rect 59426 9222 59436 9274
rect 59460 9222 59490 9274
rect 59490 9222 59516 9274
rect 59220 9220 59276 9222
rect 59300 9220 59356 9222
rect 59380 9220 59436 9222
rect 59460 9220 59516 9222
rect 59220 8186 59276 8188
rect 59300 8186 59356 8188
rect 59380 8186 59436 8188
rect 59460 8186 59516 8188
rect 59220 8134 59246 8186
rect 59246 8134 59276 8186
rect 59300 8134 59310 8186
rect 59310 8134 59356 8186
rect 59380 8134 59426 8186
rect 59426 8134 59436 8186
rect 59460 8134 59490 8186
rect 59490 8134 59516 8186
rect 59220 8132 59276 8134
rect 59300 8132 59356 8134
rect 59380 8132 59436 8134
rect 59460 8132 59516 8134
rect 59220 7098 59276 7100
rect 59300 7098 59356 7100
rect 59380 7098 59436 7100
rect 59460 7098 59516 7100
rect 59220 7046 59246 7098
rect 59246 7046 59276 7098
rect 59300 7046 59310 7098
rect 59310 7046 59356 7098
rect 59380 7046 59426 7098
rect 59426 7046 59436 7098
rect 59460 7046 59490 7098
rect 59490 7046 59516 7098
rect 59220 7044 59276 7046
rect 59300 7044 59356 7046
rect 59380 7044 59436 7046
rect 59460 7044 59516 7046
rect 59220 6010 59276 6012
rect 59300 6010 59356 6012
rect 59380 6010 59436 6012
rect 59460 6010 59516 6012
rect 59220 5958 59246 6010
rect 59246 5958 59276 6010
rect 59300 5958 59310 6010
rect 59310 5958 59356 6010
rect 59380 5958 59426 6010
rect 59426 5958 59436 6010
rect 59460 5958 59490 6010
rect 59490 5958 59516 6010
rect 59220 5956 59276 5958
rect 59300 5956 59356 5958
rect 59380 5956 59436 5958
rect 59460 5956 59516 5958
rect 64220 65306 64276 65308
rect 64300 65306 64356 65308
rect 64380 65306 64436 65308
rect 64460 65306 64516 65308
rect 64220 65254 64246 65306
rect 64246 65254 64276 65306
rect 64300 65254 64310 65306
rect 64310 65254 64356 65306
rect 64380 65254 64426 65306
rect 64426 65254 64436 65306
rect 64460 65254 64490 65306
rect 64490 65254 64516 65306
rect 64220 65252 64276 65254
rect 64300 65252 64356 65254
rect 64380 65252 64436 65254
rect 64460 65252 64516 65254
rect 64220 64218 64276 64220
rect 64300 64218 64356 64220
rect 64380 64218 64436 64220
rect 64460 64218 64516 64220
rect 64220 64166 64246 64218
rect 64246 64166 64276 64218
rect 64300 64166 64310 64218
rect 64310 64166 64356 64218
rect 64380 64166 64426 64218
rect 64426 64166 64436 64218
rect 64460 64166 64490 64218
rect 64490 64166 64516 64218
rect 64220 64164 64276 64166
rect 64300 64164 64356 64166
rect 64380 64164 64436 64166
rect 64460 64164 64516 64166
rect 64220 63130 64276 63132
rect 64300 63130 64356 63132
rect 64380 63130 64436 63132
rect 64460 63130 64516 63132
rect 64220 63078 64246 63130
rect 64246 63078 64276 63130
rect 64300 63078 64310 63130
rect 64310 63078 64356 63130
rect 64380 63078 64426 63130
rect 64426 63078 64436 63130
rect 64460 63078 64490 63130
rect 64490 63078 64516 63130
rect 64220 63076 64276 63078
rect 64300 63076 64356 63078
rect 64380 63076 64436 63078
rect 64460 63076 64516 63078
rect 64220 62042 64276 62044
rect 64300 62042 64356 62044
rect 64380 62042 64436 62044
rect 64460 62042 64516 62044
rect 64220 61990 64246 62042
rect 64246 61990 64276 62042
rect 64300 61990 64310 62042
rect 64310 61990 64356 62042
rect 64380 61990 64426 62042
rect 64426 61990 64436 62042
rect 64460 61990 64490 62042
rect 64490 61990 64516 62042
rect 64220 61988 64276 61990
rect 64300 61988 64356 61990
rect 64380 61988 64436 61990
rect 64460 61988 64516 61990
rect 64220 60954 64276 60956
rect 64300 60954 64356 60956
rect 64380 60954 64436 60956
rect 64460 60954 64516 60956
rect 64220 60902 64246 60954
rect 64246 60902 64276 60954
rect 64300 60902 64310 60954
rect 64310 60902 64356 60954
rect 64380 60902 64426 60954
rect 64426 60902 64436 60954
rect 64460 60902 64490 60954
rect 64490 60902 64516 60954
rect 64220 60900 64276 60902
rect 64300 60900 64356 60902
rect 64380 60900 64436 60902
rect 64460 60900 64516 60902
rect 64220 59866 64276 59868
rect 64300 59866 64356 59868
rect 64380 59866 64436 59868
rect 64460 59866 64516 59868
rect 64220 59814 64246 59866
rect 64246 59814 64276 59866
rect 64300 59814 64310 59866
rect 64310 59814 64356 59866
rect 64380 59814 64426 59866
rect 64426 59814 64436 59866
rect 64460 59814 64490 59866
rect 64490 59814 64516 59866
rect 64220 59812 64276 59814
rect 64300 59812 64356 59814
rect 64380 59812 64436 59814
rect 64460 59812 64516 59814
rect 59542 5616 59598 5672
rect 59220 4922 59276 4924
rect 59300 4922 59356 4924
rect 59380 4922 59436 4924
rect 59460 4922 59516 4924
rect 59220 4870 59246 4922
rect 59246 4870 59276 4922
rect 59300 4870 59310 4922
rect 59310 4870 59356 4922
rect 59380 4870 59426 4922
rect 59426 4870 59436 4922
rect 59460 4870 59490 4922
rect 59490 4870 59516 4922
rect 59220 4868 59276 4870
rect 59300 4868 59356 4870
rect 59380 4868 59436 4870
rect 59460 4868 59516 4870
rect 59220 3834 59276 3836
rect 59300 3834 59356 3836
rect 59380 3834 59436 3836
rect 59460 3834 59516 3836
rect 59220 3782 59246 3834
rect 59246 3782 59276 3834
rect 59300 3782 59310 3834
rect 59310 3782 59356 3834
rect 59380 3782 59426 3834
rect 59426 3782 59436 3834
rect 59460 3782 59490 3834
rect 59490 3782 59516 3834
rect 59220 3780 59276 3782
rect 59300 3780 59356 3782
rect 59380 3780 59436 3782
rect 59460 3780 59516 3782
rect 59220 2746 59276 2748
rect 59300 2746 59356 2748
rect 59380 2746 59436 2748
rect 59460 2746 59516 2748
rect 59220 2694 59246 2746
rect 59246 2694 59276 2746
rect 59300 2694 59310 2746
rect 59310 2694 59356 2746
rect 59380 2694 59426 2746
rect 59426 2694 59436 2746
rect 59460 2694 59490 2746
rect 59490 2694 59516 2746
rect 59220 2692 59276 2694
rect 59300 2692 59356 2694
rect 59380 2692 59436 2694
rect 59460 2692 59516 2694
rect 60646 5616 60702 5672
rect 64220 58778 64276 58780
rect 64300 58778 64356 58780
rect 64380 58778 64436 58780
rect 64460 58778 64516 58780
rect 64220 58726 64246 58778
rect 64246 58726 64276 58778
rect 64300 58726 64310 58778
rect 64310 58726 64356 58778
rect 64380 58726 64426 58778
rect 64426 58726 64436 58778
rect 64460 58726 64490 58778
rect 64490 58726 64516 58778
rect 64220 58724 64276 58726
rect 64300 58724 64356 58726
rect 64380 58724 64436 58726
rect 64460 58724 64516 58726
rect 64220 57690 64276 57692
rect 64300 57690 64356 57692
rect 64380 57690 64436 57692
rect 64460 57690 64516 57692
rect 64220 57638 64246 57690
rect 64246 57638 64276 57690
rect 64300 57638 64310 57690
rect 64310 57638 64356 57690
rect 64380 57638 64426 57690
rect 64426 57638 64436 57690
rect 64460 57638 64490 57690
rect 64490 57638 64516 57690
rect 64220 57636 64276 57638
rect 64300 57636 64356 57638
rect 64380 57636 64436 57638
rect 64460 57636 64516 57638
rect 64220 56602 64276 56604
rect 64300 56602 64356 56604
rect 64380 56602 64436 56604
rect 64460 56602 64516 56604
rect 64220 56550 64246 56602
rect 64246 56550 64276 56602
rect 64300 56550 64310 56602
rect 64310 56550 64356 56602
rect 64380 56550 64426 56602
rect 64426 56550 64436 56602
rect 64460 56550 64490 56602
rect 64490 56550 64516 56602
rect 64220 56548 64276 56550
rect 64300 56548 64356 56550
rect 64380 56548 64436 56550
rect 64460 56548 64516 56550
rect 64220 55514 64276 55516
rect 64300 55514 64356 55516
rect 64380 55514 64436 55516
rect 64460 55514 64516 55516
rect 64220 55462 64246 55514
rect 64246 55462 64276 55514
rect 64300 55462 64310 55514
rect 64310 55462 64356 55514
rect 64380 55462 64426 55514
rect 64426 55462 64436 55514
rect 64460 55462 64490 55514
rect 64490 55462 64516 55514
rect 64220 55460 64276 55462
rect 64300 55460 64356 55462
rect 64380 55460 64436 55462
rect 64460 55460 64516 55462
rect 64220 54426 64276 54428
rect 64300 54426 64356 54428
rect 64380 54426 64436 54428
rect 64460 54426 64516 54428
rect 64220 54374 64246 54426
rect 64246 54374 64276 54426
rect 64300 54374 64310 54426
rect 64310 54374 64356 54426
rect 64380 54374 64426 54426
rect 64426 54374 64436 54426
rect 64460 54374 64490 54426
rect 64490 54374 64516 54426
rect 64220 54372 64276 54374
rect 64300 54372 64356 54374
rect 64380 54372 64436 54374
rect 64460 54372 64516 54374
rect 64220 53338 64276 53340
rect 64300 53338 64356 53340
rect 64380 53338 64436 53340
rect 64460 53338 64516 53340
rect 64220 53286 64246 53338
rect 64246 53286 64276 53338
rect 64300 53286 64310 53338
rect 64310 53286 64356 53338
rect 64380 53286 64426 53338
rect 64426 53286 64436 53338
rect 64460 53286 64490 53338
rect 64490 53286 64516 53338
rect 64220 53284 64276 53286
rect 64300 53284 64356 53286
rect 64380 53284 64436 53286
rect 64460 53284 64516 53286
rect 64220 52250 64276 52252
rect 64300 52250 64356 52252
rect 64380 52250 64436 52252
rect 64460 52250 64516 52252
rect 64220 52198 64246 52250
rect 64246 52198 64276 52250
rect 64300 52198 64310 52250
rect 64310 52198 64356 52250
rect 64380 52198 64426 52250
rect 64426 52198 64436 52250
rect 64460 52198 64490 52250
rect 64490 52198 64516 52250
rect 64220 52196 64276 52198
rect 64300 52196 64356 52198
rect 64380 52196 64436 52198
rect 64460 52196 64516 52198
rect 64220 51162 64276 51164
rect 64300 51162 64356 51164
rect 64380 51162 64436 51164
rect 64460 51162 64516 51164
rect 64220 51110 64246 51162
rect 64246 51110 64276 51162
rect 64300 51110 64310 51162
rect 64310 51110 64356 51162
rect 64380 51110 64426 51162
rect 64426 51110 64436 51162
rect 64460 51110 64490 51162
rect 64490 51110 64516 51162
rect 64220 51108 64276 51110
rect 64300 51108 64356 51110
rect 64380 51108 64436 51110
rect 64460 51108 64516 51110
rect 64220 50074 64276 50076
rect 64300 50074 64356 50076
rect 64380 50074 64436 50076
rect 64460 50074 64516 50076
rect 64220 50022 64246 50074
rect 64246 50022 64276 50074
rect 64300 50022 64310 50074
rect 64310 50022 64356 50074
rect 64380 50022 64426 50074
rect 64426 50022 64436 50074
rect 64460 50022 64490 50074
rect 64490 50022 64516 50074
rect 64220 50020 64276 50022
rect 64300 50020 64356 50022
rect 64380 50020 64436 50022
rect 64460 50020 64516 50022
rect 64220 48986 64276 48988
rect 64300 48986 64356 48988
rect 64380 48986 64436 48988
rect 64460 48986 64516 48988
rect 64220 48934 64246 48986
rect 64246 48934 64276 48986
rect 64300 48934 64310 48986
rect 64310 48934 64356 48986
rect 64380 48934 64426 48986
rect 64426 48934 64436 48986
rect 64460 48934 64490 48986
rect 64490 48934 64516 48986
rect 64220 48932 64276 48934
rect 64300 48932 64356 48934
rect 64380 48932 64436 48934
rect 64460 48932 64516 48934
rect 64220 47898 64276 47900
rect 64300 47898 64356 47900
rect 64380 47898 64436 47900
rect 64460 47898 64516 47900
rect 64220 47846 64246 47898
rect 64246 47846 64276 47898
rect 64300 47846 64310 47898
rect 64310 47846 64356 47898
rect 64380 47846 64426 47898
rect 64426 47846 64436 47898
rect 64460 47846 64490 47898
rect 64490 47846 64516 47898
rect 64220 47844 64276 47846
rect 64300 47844 64356 47846
rect 64380 47844 64436 47846
rect 64460 47844 64516 47846
rect 64220 46810 64276 46812
rect 64300 46810 64356 46812
rect 64380 46810 64436 46812
rect 64460 46810 64516 46812
rect 64220 46758 64246 46810
rect 64246 46758 64276 46810
rect 64300 46758 64310 46810
rect 64310 46758 64356 46810
rect 64380 46758 64426 46810
rect 64426 46758 64436 46810
rect 64460 46758 64490 46810
rect 64490 46758 64516 46810
rect 64220 46756 64276 46758
rect 64300 46756 64356 46758
rect 64380 46756 64436 46758
rect 64460 46756 64516 46758
rect 64220 45722 64276 45724
rect 64300 45722 64356 45724
rect 64380 45722 64436 45724
rect 64460 45722 64516 45724
rect 64220 45670 64246 45722
rect 64246 45670 64276 45722
rect 64300 45670 64310 45722
rect 64310 45670 64356 45722
rect 64380 45670 64426 45722
rect 64426 45670 64436 45722
rect 64460 45670 64490 45722
rect 64490 45670 64516 45722
rect 64220 45668 64276 45670
rect 64300 45668 64356 45670
rect 64380 45668 64436 45670
rect 64460 45668 64516 45670
rect 64220 44634 64276 44636
rect 64300 44634 64356 44636
rect 64380 44634 64436 44636
rect 64460 44634 64516 44636
rect 64220 44582 64246 44634
rect 64246 44582 64276 44634
rect 64300 44582 64310 44634
rect 64310 44582 64356 44634
rect 64380 44582 64426 44634
rect 64426 44582 64436 44634
rect 64460 44582 64490 44634
rect 64490 44582 64516 44634
rect 64220 44580 64276 44582
rect 64300 44580 64356 44582
rect 64380 44580 64436 44582
rect 64460 44580 64516 44582
rect 64220 43546 64276 43548
rect 64300 43546 64356 43548
rect 64380 43546 64436 43548
rect 64460 43546 64516 43548
rect 64220 43494 64246 43546
rect 64246 43494 64276 43546
rect 64300 43494 64310 43546
rect 64310 43494 64356 43546
rect 64380 43494 64426 43546
rect 64426 43494 64436 43546
rect 64460 43494 64490 43546
rect 64490 43494 64516 43546
rect 64220 43492 64276 43494
rect 64300 43492 64356 43494
rect 64380 43492 64436 43494
rect 64460 43492 64516 43494
rect 64220 42458 64276 42460
rect 64300 42458 64356 42460
rect 64380 42458 64436 42460
rect 64460 42458 64516 42460
rect 64220 42406 64246 42458
rect 64246 42406 64276 42458
rect 64300 42406 64310 42458
rect 64310 42406 64356 42458
rect 64380 42406 64426 42458
rect 64426 42406 64436 42458
rect 64460 42406 64490 42458
rect 64490 42406 64516 42458
rect 64220 42404 64276 42406
rect 64300 42404 64356 42406
rect 64380 42404 64436 42406
rect 64460 42404 64516 42406
rect 64220 41370 64276 41372
rect 64300 41370 64356 41372
rect 64380 41370 64436 41372
rect 64460 41370 64516 41372
rect 64220 41318 64246 41370
rect 64246 41318 64276 41370
rect 64300 41318 64310 41370
rect 64310 41318 64356 41370
rect 64380 41318 64426 41370
rect 64426 41318 64436 41370
rect 64460 41318 64490 41370
rect 64490 41318 64516 41370
rect 64220 41316 64276 41318
rect 64300 41316 64356 41318
rect 64380 41316 64436 41318
rect 64460 41316 64516 41318
rect 64220 40282 64276 40284
rect 64300 40282 64356 40284
rect 64380 40282 64436 40284
rect 64460 40282 64516 40284
rect 64220 40230 64246 40282
rect 64246 40230 64276 40282
rect 64300 40230 64310 40282
rect 64310 40230 64356 40282
rect 64380 40230 64426 40282
rect 64426 40230 64436 40282
rect 64460 40230 64490 40282
rect 64490 40230 64516 40282
rect 64220 40228 64276 40230
rect 64300 40228 64356 40230
rect 64380 40228 64436 40230
rect 64460 40228 64516 40230
rect 64220 39194 64276 39196
rect 64300 39194 64356 39196
rect 64380 39194 64436 39196
rect 64460 39194 64516 39196
rect 64220 39142 64246 39194
rect 64246 39142 64276 39194
rect 64300 39142 64310 39194
rect 64310 39142 64356 39194
rect 64380 39142 64426 39194
rect 64426 39142 64436 39194
rect 64460 39142 64490 39194
rect 64490 39142 64516 39194
rect 64220 39140 64276 39142
rect 64300 39140 64356 39142
rect 64380 39140 64436 39142
rect 64460 39140 64516 39142
rect 64220 38106 64276 38108
rect 64300 38106 64356 38108
rect 64380 38106 64436 38108
rect 64460 38106 64516 38108
rect 64220 38054 64246 38106
rect 64246 38054 64276 38106
rect 64300 38054 64310 38106
rect 64310 38054 64356 38106
rect 64380 38054 64426 38106
rect 64426 38054 64436 38106
rect 64460 38054 64490 38106
rect 64490 38054 64516 38106
rect 64220 38052 64276 38054
rect 64300 38052 64356 38054
rect 64380 38052 64436 38054
rect 64460 38052 64516 38054
rect 64220 37018 64276 37020
rect 64300 37018 64356 37020
rect 64380 37018 64436 37020
rect 64460 37018 64516 37020
rect 64220 36966 64246 37018
rect 64246 36966 64276 37018
rect 64300 36966 64310 37018
rect 64310 36966 64356 37018
rect 64380 36966 64426 37018
rect 64426 36966 64436 37018
rect 64460 36966 64490 37018
rect 64490 36966 64516 37018
rect 64220 36964 64276 36966
rect 64300 36964 64356 36966
rect 64380 36964 64436 36966
rect 64460 36964 64516 36966
rect 64220 35930 64276 35932
rect 64300 35930 64356 35932
rect 64380 35930 64436 35932
rect 64460 35930 64516 35932
rect 64220 35878 64246 35930
rect 64246 35878 64276 35930
rect 64300 35878 64310 35930
rect 64310 35878 64356 35930
rect 64380 35878 64426 35930
rect 64426 35878 64436 35930
rect 64460 35878 64490 35930
rect 64490 35878 64516 35930
rect 64220 35876 64276 35878
rect 64300 35876 64356 35878
rect 64380 35876 64436 35878
rect 64460 35876 64516 35878
rect 64220 34842 64276 34844
rect 64300 34842 64356 34844
rect 64380 34842 64436 34844
rect 64460 34842 64516 34844
rect 64220 34790 64246 34842
rect 64246 34790 64276 34842
rect 64300 34790 64310 34842
rect 64310 34790 64356 34842
rect 64380 34790 64426 34842
rect 64426 34790 64436 34842
rect 64460 34790 64490 34842
rect 64490 34790 64516 34842
rect 64220 34788 64276 34790
rect 64300 34788 64356 34790
rect 64380 34788 64436 34790
rect 64460 34788 64516 34790
rect 64220 33754 64276 33756
rect 64300 33754 64356 33756
rect 64380 33754 64436 33756
rect 64460 33754 64516 33756
rect 64220 33702 64246 33754
rect 64246 33702 64276 33754
rect 64300 33702 64310 33754
rect 64310 33702 64356 33754
rect 64380 33702 64426 33754
rect 64426 33702 64436 33754
rect 64460 33702 64490 33754
rect 64490 33702 64516 33754
rect 64220 33700 64276 33702
rect 64300 33700 64356 33702
rect 64380 33700 64436 33702
rect 64460 33700 64516 33702
rect 64220 32666 64276 32668
rect 64300 32666 64356 32668
rect 64380 32666 64436 32668
rect 64460 32666 64516 32668
rect 64220 32614 64246 32666
rect 64246 32614 64276 32666
rect 64300 32614 64310 32666
rect 64310 32614 64356 32666
rect 64380 32614 64426 32666
rect 64426 32614 64436 32666
rect 64460 32614 64490 32666
rect 64490 32614 64516 32666
rect 64220 32612 64276 32614
rect 64300 32612 64356 32614
rect 64380 32612 64436 32614
rect 64460 32612 64516 32614
rect 64220 31578 64276 31580
rect 64300 31578 64356 31580
rect 64380 31578 64436 31580
rect 64460 31578 64516 31580
rect 64220 31526 64246 31578
rect 64246 31526 64276 31578
rect 64300 31526 64310 31578
rect 64310 31526 64356 31578
rect 64380 31526 64426 31578
rect 64426 31526 64436 31578
rect 64460 31526 64490 31578
rect 64490 31526 64516 31578
rect 64220 31524 64276 31526
rect 64300 31524 64356 31526
rect 64380 31524 64436 31526
rect 64460 31524 64516 31526
rect 64220 30490 64276 30492
rect 64300 30490 64356 30492
rect 64380 30490 64436 30492
rect 64460 30490 64516 30492
rect 64220 30438 64246 30490
rect 64246 30438 64276 30490
rect 64300 30438 64310 30490
rect 64310 30438 64356 30490
rect 64380 30438 64426 30490
rect 64426 30438 64436 30490
rect 64460 30438 64490 30490
rect 64490 30438 64516 30490
rect 64220 30436 64276 30438
rect 64300 30436 64356 30438
rect 64380 30436 64436 30438
rect 64460 30436 64516 30438
rect 64220 29402 64276 29404
rect 64300 29402 64356 29404
rect 64380 29402 64436 29404
rect 64460 29402 64516 29404
rect 64220 29350 64246 29402
rect 64246 29350 64276 29402
rect 64300 29350 64310 29402
rect 64310 29350 64356 29402
rect 64380 29350 64426 29402
rect 64426 29350 64436 29402
rect 64460 29350 64490 29402
rect 64490 29350 64516 29402
rect 64220 29348 64276 29350
rect 64300 29348 64356 29350
rect 64380 29348 64436 29350
rect 64460 29348 64516 29350
rect 64220 28314 64276 28316
rect 64300 28314 64356 28316
rect 64380 28314 64436 28316
rect 64460 28314 64516 28316
rect 64220 28262 64246 28314
rect 64246 28262 64276 28314
rect 64300 28262 64310 28314
rect 64310 28262 64356 28314
rect 64380 28262 64426 28314
rect 64426 28262 64436 28314
rect 64460 28262 64490 28314
rect 64490 28262 64516 28314
rect 64220 28260 64276 28262
rect 64300 28260 64356 28262
rect 64380 28260 64436 28262
rect 64460 28260 64516 28262
rect 64220 27226 64276 27228
rect 64300 27226 64356 27228
rect 64380 27226 64436 27228
rect 64460 27226 64516 27228
rect 64220 27174 64246 27226
rect 64246 27174 64276 27226
rect 64300 27174 64310 27226
rect 64310 27174 64356 27226
rect 64380 27174 64426 27226
rect 64426 27174 64436 27226
rect 64460 27174 64490 27226
rect 64490 27174 64516 27226
rect 64220 27172 64276 27174
rect 64300 27172 64356 27174
rect 64380 27172 64436 27174
rect 64460 27172 64516 27174
rect 64220 26138 64276 26140
rect 64300 26138 64356 26140
rect 64380 26138 64436 26140
rect 64460 26138 64516 26140
rect 64220 26086 64246 26138
rect 64246 26086 64276 26138
rect 64300 26086 64310 26138
rect 64310 26086 64356 26138
rect 64380 26086 64426 26138
rect 64426 26086 64436 26138
rect 64460 26086 64490 26138
rect 64490 26086 64516 26138
rect 64220 26084 64276 26086
rect 64300 26084 64356 26086
rect 64380 26084 64436 26086
rect 64460 26084 64516 26086
rect 64220 25050 64276 25052
rect 64300 25050 64356 25052
rect 64380 25050 64436 25052
rect 64460 25050 64516 25052
rect 64220 24998 64246 25050
rect 64246 24998 64276 25050
rect 64300 24998 64310 25050
rect 64310 24998 64356 25050
rect 64380 24998 64426 25050
rect 64426 24998 64436 25050
rect 64460 24998 64490 25050
rect 64490 24998 64516 25050
rect 64220 24996 64276 24998
rect 64300 24996 64356 24998
rect 64380 24996 64436 24998
rect 64460 24996 64516 24998
rect 64220 23962 64276 23964
rect 64300 23962 64356 23964
rect 64380 23962 64436 23964
rect 64460 23962 64516 23964
rect 64220 23910 64246 23962
rect 64246 23910 64276 23962
rect 64300 23910 64310 23962
rect 64310 23910 64356 23962
rect 64380 23910 64426 23962
rect 64426 23910 64436 23962
rect 64460 23910 64490 23962
rect 64490 23910 64516 23962
rect 64220 23908 64276 23910
rect 64300 23908 64356 23910
rect 64380 23908 64436 23910
rect 64460 23908 64516 23910
rect 64220 22874 64276 22876
rect 64300 22874 64356 22876
rect 64380 22874 64436 22876
rect 64460 22874 64516 22876
rect 64220 22822 64246 22874
rect 64246 22822 64276 22874
rect 64300 22822 64310 22874
rect 64310 22822 64356 22874
rect 64380 22822 64426 22874
rect 64426 22822 64436 22874
rect 64460 22822 64490 22874
rect 64490 22822 64516 22874
rect 64220 22820 64276 22822
rect 64300 22820 64356 22822
rect 64380 22820 64436 22822
rect 64460 22820 64516 22822
rect 64220 21786 64276 21788
rect 64300 21786 64356 21788
rect 64380 21786 64436 21788
rect 64460 21786 64516 21788
rect 64220 21734 64246 21786
rect 64246 21734 64276 21786
rect 64300 21734 64310 21786
rect 64310 21734 64356 21786
rect 64380 21734 64426 21786
rect 64426 21734 64436 21786
rect 64460 21734 64490 21786
rect 64490 21734 64516 21786
rect 64220 21732 64276 21734
rect 64300 21732 64356 21734
rect 64380 21732 64436 21734
rect 64460 21732 64516 21734
rect 64220 20698 64276 20700
rect 64300 20698 64356 20700
rect 64380 20698 64436 20700
rect 64460 20698 64516 20700
rect 64220 20646 64246 20698
rect 64246 20646 64276 20698
rect 64300 20646 64310 20698
rect 64310 20646 64356 20698
rect 64380 20646 64426 20698
rect 64426 20646 64436 20698
rect 64460 20646 64490 20698
rect 64490 20646 64516 20698
rect 64220 20644 64276 20646
rect 64300 20644 64356 20646
rect 64380 20644 64436 20646
rect 64460 20644 64516 20646
rect 64220 19610 64276 19612
rect 64300 19610 64356 19612
rect 64380 19610 64436 19612
rect 64460 19610 64516 19612
rect 64220 19558 64246 19610
rect 64246 19558 64276 19610
rect 64300 19558 64310 19610
rect 64310 19558 64356 19610
rect 64380 19558 64426 19610
rect 64426 19558 64436 19610
rect 64460 19558 64490 19610
rect 64490 19558 64516 19610
rect 64220 19556 64276 19558
rect 64300 19556 64356 19558
rect 64380 19556 64436 19558
rect 64460 19556 64516 19558
rect 64220 18522 64276 18524
rect 64300 18522 64356 18524
rect 64380 18522 64436 18524
rect 64460 18522 64516 18524
rect 64220 18470 64246 18522
rect 64246 18470 64276 18522
rect 64300 18470 64310 18522
rect 64310 18470 64356 18522
rect 64380 18470 64426 18522
rect 64426 18470 64436 18522
rect 64460 18470 64490 18522
rect 64490 18470 64516 18522
rect 64220 18468 64276 18470
rect 64300 18468 64356 18470
rect 64380 18468 64436 18470
rect 64460 18468 64516 18470
rect 64220 17434 64276 17436
rect 64300 17434 64356 17436
rect 64380 17434 64436 17436
rect 64460 17434 64516 17436
rect 64220 17382 64246 17434
rect 64246 17382 64276 17434
rect 64300 17382 64310 17434
rect 64310 17382 64356 17434
rect 64380 17382 64426 17434
rect 64426 17382 64436 17434
rect 64460 17382 64490 17434
rect 64490 17382 64516 17434
rect 64220 17380 64276 17382
rect 64300 17380 64356 17382
rect 64380 17380 64436 17382
rect 64460 17380 64516 17382
rect 64220 16346 64276 16348
rect 64300 16346 64356 16348
rect 64380 16346 64436 16348
rect 64460 16346 64516 16348
rect 64220 16294 64246 16346
rect 64246 16294 64276 16346
rect 64300 16294 64310 16346
rect 64310 16294 64356 16346
rect 64380 16294 64426 16346
rect 64426 16294 64436 16346
rect 64460 16294 64490 16346
rect 64490 16294 64516 16346
rect 64220 16292 64276 16294
rect 64300 16292 64356 16294
rect 64380 16292 64436 16294
rect 64460 16292 64516 16294
rect 64220 15258 64276 15260
rect 64300 15258 64356 15260
rect 64380 15258 64436 15260
rect 64460 15258 64516 15260
rect 64220 15206 64246 15258
rect 64246 15206 64276 15258
rect 64300 15206 64310 15258
rect 64310 15206 64356 15258
rect 64380 15206 64426 15258
rect 64426 15206 64436 15258
rect 64460 15206 64490 15258
rect 64490 15206 64516 15258
rect 64220 15204 64276 15206
rect 64300 15204 64356 15206
rect 64380 15204 64436 15206
rect 64460 15204 64516 15206
rect 64220 14170 64276 14172
rect 64300 14170 64356 14172
rect 64380 14170 64436 14172
rect 64460 14170 64516 14172
rect 64220 14118 64246 14170
rect 64246 14118 64276 14170
rect 64300 14118 64310 14170
rect 64310 14118 64356 14170
rect 64380 14118 64426 14170
rect 64426 14118 64436 14170
rect 64460 14118 64490 14170
rect 64490 14118 64516 14170
rect 64220 14116 64276 14118
rect 64300 14116 64356 14118
rect 64380 14116 64436 14118
rect 64460 14116 64516 14118
rect 64220 13082 64276 13084
rect 64300 13082 64356 13084
rect 64380 13082 64436 13084
rect 64460 13082 64516 13084
rect 64220 13030 64246 13082
rect 64246 13030 64276 13082
rect 64300 13030 64310 13082
rect 64310 13030 64356 13082
rect 64380 13030 64426 13082
rect 64426 13030 64436 13082
rect 64460 13030 64490 13082
rect 64490 13030 64516 13082
rect 64220 13028 64276 13030
rect 64300 13028 64356 13030
rect 64380 13028 64436 13030
rect 64460 13028 64516 13030
rect 64220 11994 64276 11996
rect 64300 11994 64356 11996
rect 64380 11994 64436 11996
rect 64460 11994 64516 11996
rect 64220 11942 64246 11994
rect 64246 11942 64276 11994
rect 64300 11942 64310 11994
rect 64310 11942 64356 11994
rect 64380 11942 64426 11994
rect 64426 11942 64436 11994
rect 64460 11942 64490 11994
rect 64490 11942 64516 11994
rect 64220 11940 64276 11942
rect 64300 11940 64356 11942
rect 64380 11940 64436 11942
rect 64460 11940 64516 11942
rect 64220 10906 64276 10908
rect 64300 10906 64356 10908
rect 64380 10906 64436 10908
rect 64460 10906 64516 10908
rect 64220 10854 64246 10906
rect 64246 10854 64276 10906
rect 64300 10854 64310 10906
rect 64310 10854 64356 10906
rect 64380 10854 64426 10906
rect 64426 10854 64436 10906
rect 64460 10854 64490 10906
rect 64490 10854 64516 10906
rect 64220 10852 64276 10854
rect 64300 10852 64356 10854
rect 64380 10852 64436 10854
rect 64460 10852 64516 10854
rect 65154 33496 65210 33552
rect 64220 9818 64276 9820
rect 64300 9818 64356 9820
rect 64380 9818 64436 9820
rect 64460 9818 64516 9820
rect 64220 9766 64246 9818
rect 64246 9766 64276 9818
rect 64300 9766 64310 9818
rect 64310 9766 64356 9818
rect 64380 9766 64426 9818
rect 64426 9766 64436 9818
rect 64460 9766 64490 9818
rect 64490 9766 64516 9818
rect 64220 9764 64276 9766
rect 64300 9764 64356 9766
rect 64380 9764 64436 9766
rect 64460 9764 64516 9766
rect 64220 8730 64276 8732
rect 64300 8730 64356 8732
rect 64380 8730 64436 8732
rect 64460 8730 64516 8732
rect 64220 8678 64246 8730
rect 64246 8678 64276 8730
rect 64300 8678 64310 8730
rect 64310 8678 64356 8730
rect 64380 8678 64426 8730
rect 64426 8678 64436 8730
rect 64460 8678 64490 8730
rect 64490 8678 64516 8730
rect 64220 8676 64276 8678
rect 64300 8676 64356 8678
rect 64380 8676 64436 8678
rect 64460 8676 64516 8678
rect 64220 7642 64276 7644
rect 64300 7642 64356 7644
rect 64380 7642 64436 7644
rect 64460 7642 64516 7644
rect 64220 7590 64246 7642
rect 64246 7590 64276 7642
rect 64300 7590 64310 7642
rect 64310 7590 64356 7642
rect 64380 7590 64426 7642
rect 64426 7590 64436 7642
rect 64460 7590 64490 7642
rect 64490 7590 64516 7642
rect 64220 7588 64276 7590
rect 64300 7588 64356 7590
rect 64380 7588 64436 7590
rect 64460 7588 64516 7590
rect 64220 6554 64276 6556
rect 64300 6554 64356 6556
rect 64380 6554 64436 6556
rect 64460 6554 64516 6556
rect 64220 6502 64246 6554
rect 64246 6502 64276 6554
rect 64300 6502 64310 6554
rect 64310 6502 64356 6554
rect 64380 6502 64426 6554
rect 64426 6502 64436 6554
rect 64460 6502 64490 6554
rect 64490 6502 64516 6554
rect 64220 6500 64276 6502
rect 64300 6500 64356 6502
rect 64380 6500 64436 6502
rect 64460 6500 64516 6502
rect 64220 5466 64276 5468
rect 64300 5466 64356 5468
rect 64380 5466 64436 5468
rect 64460 5466 64516 5468
rect 64220 5414 64246 5466
rect 64246 5414 64276 5466
rect 64300 5414 64310 5466
rect 64310 5414 64356 5466
rect 64380 5414 64426 5466
rect 64426 5414 64436 5466
rect 64460 5414 64490 5466
rect 64490 5414 64516 5466
rect 64220 5412 64276 5414
rect 64300 5412 64356 5414
rect 64380 5412 64436 5414
rect 64460 5412 64516 5414
rect 64220 4378 64276 4380
rect 64300 4378 64356 4380
rect 64380 4378 64436 4380
rect 64460 4378 64516 4380
rect 64220 4326 64246 4378
rect 64246 4326 64276 4378
rect 64300 4326 64310 4378
rect 64310 4326 64356 4378
rect 64380 4326 64426 4378
rect 64426 4326 64436 4378
rect 64460 4326 64490 4378
rect 64490 4326 64516 4378
rect 64220 4324 64276 4326
rect 64300 4324 64356 4326
rect 64380 4324 64436 4326
rect 64460 4324 64516 4326
rect 64220 3290 64276 3292
rect 64300 3290 64356 3292
rect 64380 3290 64436 3292
rect 64460 3290 64516 3292
rect 64220 3238 64246 3290
rect 64246 3238 64276 3290
rect 64300 3238 64310 3290
rect 64310 3238 64356 3290
rect 64380 3238 64426 3290
rect 64426 3238 64436 3290
rect 64460 3238 64490 3290
rect 64490 3238 64516 3290
rect 64220 3236 64276 3238
rect 64300 3236 64356 3238
rect 64380 3236 64436 3238
rect 64460 3236 64516 3238
rect 64220 2202 64276 2204
rect 64300 2202 64356 2204
rect 64380 2202 64436 2204
rect 64460 2202 64516 2204
rect 64220 2150 64246 2202
rect 64246 2150 64276 2202
rect 64300 2150 64310 2202
rect 64310 2150 64356 2202
rect 64380 2150 64426 2202
rect 64426 2150 64436 2202
rect 64460 2150 64490 2202
rect 64490 2150 64516 2202
rect 64220 2148 64276 2150
rect 64300 2148 64356 2150
rect 64380 2148 64436 2150
rect 64460 2148 64516 2150
rect 64326 1944 64382 2000
rect 64694 4528 64750 4584
rect 68098 66544 68154 66600
rect 65246 6840 65302 6896
rect 65246 6160 65302 6216
rect 65154 3848 65210 3904
rect 65522 3440 65578 3496
rect 66166 28328 66222 28384
rect 65798 6840 65854 6896
rect 2870 584 2926 640
rect 68098 63980 68154 64016
rect 68098 63960 68100 63980
rect 68100 63960 68152 63980
rect 68152 63960 68154 63980
rect 68098 62600 68154 62656
rect 68098 61260 68154 61296
rect 68098 61240 68100 61260
rect 68100 61240 68152 61260
rect 68152 61240 68154 61260
rect 68098 58656 68154 58712
rect 68098 57316 68154 57352
rect 68098 57296 68100 57316
rect 68100 57296 68152 57316
rect 68152 57296 68154 57316
rect 68098 56072 68154 56128
rect 68098 53352 68154 53408
rect 68098 52012 68154 52048
rect 68098 51992 68100 52012
rect 68100 51992 68152 52012
rect 68152 51992 68154 52012
rect 68098 50804 68100 50824
rect 68100 50804 68152 50824
rect 68152 50804 68154 50824
rect 68098 50768 68154 50804
rect 68098 48068 68154 48104
rect 68098 48048 68100 48068
rect 68100 48048 68152 48068
rect 68152 48048 68154 48068
rect 68098 46824 68154 46880
rect 68098 45464 68154 45520
rect 68098 42764 68154 42800
rect 68098 42744 68100 42764
rect 68100 42744 68152 42764
rect 68152 42744 68154 42764
rect 68098 41540 68154 41576
rect 68098 41520 68100 41540
rect 68100 41520 68152 41540
rect 68152 41520 68154 41540
rect 68098 40160 68154 40216
rect 68098 37576 68154 37632
rect 68098 36236 68154 36272
rect 68098 36216 68100 36236
rect 68100 36216 68152 36236
rect 68152 36216 68154 36236
rect 68926 34892 68928 34912
rect 68928 34892 68980 34912
rect 68980 34892 68982 34912
rect 68926 34856 68982 34892
rect 68098 32292 68154 32328
rect 68098 32272 68100 32292
rect 68100 32272 68152 32292
rect 68152 32272 68154 32292
rect 68098 30912 68154 30968
rect 68098 29552 68154 29608
rect 68098 26988 68154 27024
rect 68098 26968 68100 26988
rect 68100 26968 68152 26988
rect 68152 26968 68154 26988
rect 68098 25608 68154 25664
rect 68098 24248 68154 24304
rect 68098 23044 68154 23080
rect 68098 23024 68100 23044
rect 68100 23024 68152 23044
rect 68152 23024 68154 23044
rect 68098 21664 68154 21720
rect 68098 20340 68100 20360
rect 68100 20340 68152 20360
rect 68152 20340 68154 20360
rect 68098 20304 68154 20340
rect 68098 19080 68154 19136
rect 68098 17740 68154 17776
rect 68098 17720 68100 17740
rect 68100 17720 68152 17740
rect 68152 17720 68154 17740
rect 68098 16360 68154 16416
rect 68098 15020 68154 15056
rect 68098 15000 68100 15020
rect 68100 15000 68152 15020
rect 68152 15000 68154 15020
rect 68098 13812 68100 13832
rect 68100 13812 68152 13832
rect 68152 13812 68154 13832
rect 68098 13776 68154 13812
rect 68098 12416 68154 12472
rect 67546 4528 67602 4584
rect 67454 3576 67510 3632
rect 67454 3168 67510 3224
rect 68098 11076 68154 11112
rect 68098 11056 68100 11076
rect 68100 11056 68152 11076
rect 68152 11056 68154 11076
rect 68098 9832 68154 9888
rect 68098 8472 68154 8528
rect 68098 7112 68154 7168
rect 68098 5772 68154 5808
rect 68098 5752 68100 5772
rect 68100 5752 68152 5772
rect 68152 5752 68154 5772
rect 68282 5072 68338 5128
rect 68098 3168 68154 3224
rect 68190 1808 68246 1864
rect 66074 584 66130 640
<< metal3 >>
rect 0 69232 800 69352
rect 67357 69322 67423 69325
rect 69200 69322 70000 69352
rect 67357 69320 70000 69322
rect 67357 69264 67362 69320
rect 67418 69264 70000 69320
rect 67357 69262 70000 69264
rect 67357 69259 67423 69262
rect 69200 69232 70000 69262
rect 0 67962 800 67992
rect 2773 67962 2839 67965
rect 0 67960 2839 67962
rect 0 67904 2778 67960
rect 2834 67904 2839 67960
rect 0 67902 2839 67904
rect 0 67872 800 67902
rect 2773 67899 2839 67902
rect 67541 67962 67607 67965
rect 69200 67962 70000 67992
rect 67541 67960 70000 67962
rect 67541 67904 67546 67960
rect 67602 67904 70000 67960
rect 67541 67902 70000 67904
rect 67541 67899 67607 67902
rect 69200 67872 70000 67902
rect 4208 67488 4528 67489
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 14208 67488 14528 67489
rect 14208 67424 14216 67488
rect 14280 67424 14296 67488
rect 14360 67424 14376 67488
rect 14440 67424 14456 67488
rect 14520 67424 14528 67488
rect 14208 67423 14528 67424
rect 24208 67488 24528 67489
rect 24208 67424 24216 67488
rect 24280 67424 24296 67488
rect 24360 67424 24376 67488
rect 24440 67424 24456 67488
rect 24520 67424 24528 67488
rect 24208 67423 24528 67424
rect 34208 67488 34528 67489
rect 34208 67424 34216 67488
rect 34280 67424 34296 67488
rect 34360 67424 34376 67488
rect 34440 67424 34456 67488
rect 34520 67424 34528 67488
rect 34208 67423 34528 67424
rect 44208 67488 44528 67489
rect 44208 67424 44216 67488
rect 44280 67424 44296 67488
rect 44360 67424 44376 67488
rect 44440 67424 44456 67488
rect 44520 67424 44528 67488
rect 44208 67423 44528 67424
rect 54208 67488 54528 67489
rect 54208 67424 54216 67488
rect 54280 67424 54296 67488
rect 54360 67424 54376 67488
rect 54440 67424 54456 67488
rect 54520 67424 54528 67488
rect 54208 67423 54528 67424
rect 64208 67488 64528 67489
rect 64208 67424 64216 67488
rect 64280 67424 64296 67488
rect 64360 67424 64376 67488
rect 64440 67424 64456 67488
rect 64520 67424 64528 67488
rect 64208 67423 64528 67424
rect 9208 66944 9528 66945
rect 9208 66880 9216 66944
rect 9280 66880 9296 66944
rect 9360 66880 9376 66944
rect 9440 66880 9456 66944
rect 9520 66880 9528 66944
rect 9208 66879 9528 66880
rect 19208 66944 19528 66945
rect 19208 66880 19216 66944
rect 19280 66880 19296 66944
rect 19360 66880 19376 66944
rect 19440 66880 19456 66944
rect 19520 66880 19528 66944
rect 19208 66879 19528 66880
rect 29208 66944 29528 66945
rect 29208 66880 29216 66944
rect 29280 66880 29296 66944
rect 29360 66880 29376 66944
rect 29440 66880 29456 66944
rect 29520 66880 29528 66944
rect 29208 66879 29528 66880
rect 39208 66944 39528 66945
rect 39208 66880 39216 66944
rect 39280 66880 39296 66944
rect 39360 66880 39376 66944
rect 39440 66880 39456 66944
rect 39520 66880 39528 66944
rect 39208 66879 39528 66880
rect 49208 66944 49528 66945
rect 49208 66880 49216 66944
rect 49280 66880 49296 66944
rect 49360 66880 49376 66944
rect 49440 66880 49456 66944
rect 49520 66880 49528 66944
rect 49208 66879 49528 66880
rect 59208 66944 59528 66945
rect 59208 66880 59216 66944
rect 59280 66880 59296 66944
rect 59360 66880 59376 66944
rect 59440 66880 59456 66944
rect 59520 66880 59528 66944
rect 59208 66879 59528 66880
rect 0 66738 800 66768
rect 1761 66738 1827 66741
rect 0 66736 1827 66738
rect 0 66680 1766 66736
rect 1822 66680 1827 66736
rect 0 66678 1827 66680
rect 0 66648 800 66678
rect 1761 66675 1827 66678
rect 68093 66602 68159 66605
rect 69200 66602 70000 66632
rect 68093 66600 70000 66602
rect 68093 66544 68098 66600
rect 68154 66544 70000 66600
rect 68093 66542 70000 66544
rect 68093 66539 68159 66542
rect 69200 66512 70000 66542
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 14208 66400 14528 66401
rect 14208 66336 14216 66400
rect 14280 66336 14296 66400
rect 14360 66336 14376 66400
rect 14440 66336 14456 66400
rect 14520 66336 14528 66400
rect 14208 66335 14528 66336
rect 24208 66400 24528 66401
rect 24208 66336 24216 66400
rect 24280 66336 24296 66400
rect 24360 66336 24376 66400
rect 24440 66336 24456 66400
rect 24520 66336 24528 66400
rect 24208 66335 24528 66336
rect 34208 66400 34528 66401
rect 34208 66336 34216 66400
rect 34280 66336 34296 66400
rect 34360 66336 34376 66400
rect 34440 66336 34456 66400
rect 34520 66336 34528 66400
rect 34208 66335 34528 66336
rect 44208 66400 44528 66401
rect 44208 66336 44216 66400
rect 44280 66336 44296 66400
rect 44360 66336 44376 66400
rect 44440 66336 44456 66400
rect 44520 66336 44528 66400
rect 44208 66335 44528 66336
rect 54208 66400 54528 66401
rect 54208 66336 54216 66400
rect 54280 66336 54296 66400
rect 54360 66336 54376 66400
rect 54440 66336 54456 66400
rect 54520 66336 54528 66400
rect 54208 66335 54528 66336
rect 64208 66400 64528 66401
rect 64208 66336 64216 66400
rect 64280 66336 64296 66400
rect 64360 66336 64376 66400
rect 64440 66336 64456 66400
rect 64520 66336 64528 66400
rect 64208 66335 64528 66336
rect 9208 65856 9528 65857
rect 9208 65792 9216 65856
rect 9280 65792 9296 65856
rect 9360 65792 9376 65856
rect 9440 65792 9456 65856
rect 9520 65792 9528 65856
rect 9208 65791 9528 65792
rect 19208 65856 19528 65857
rect 19208 65792 19216 65856
rect 19280 65792 19296 65856
rect 19360 65792 19376 65856
rect 19440 65792 19456 65856
rect 19520 65792 19528 65856
rect 19208 65791 19528 65792
rect 29208 65856 29528 65857
rect 29208 65792 29216 65856
rect 29280 65792 29296 65856
rect 29360 65792 29376 65856
rect 29440 65792 29456 65856
rect 29520 65792 29528 65856
rect 29208 65791 29528 65792
rect 39208 65856 39528 65857
rect 39208 65792 39216 65856
rect 39280 65792 39296 65856
rect 39360 65792 39376 65856
rect 39440 65792 39456 65856
rect 39520 65792 39528 65856
rect 39208 65791 39528 65792
rect 49208 65856 49528 65857
rect 49208 65792 49216 65856
rect 49280 65792 49296 65856
rect 49360 65792 49376 65856
rect 49440 65792 49456 65856
rect 49520 65792 49528 65856
rect 49208 65791 49528 65792
rect 59208 65856 59528 65857
rect 59208 65792 59216 65856
rect 59280 65792 59296 65856
rect 59360 65792 59376 65856
rect 59440 65792 59456 65856
rect 59520 65792 59528 65856
rect 59208 65791 59528 65792
rect 0 65378 800 65408
rect 1853 65378 1919 65381
rect 0 65376 1919 65378
rect 0 65320 1858 65376
rect 1914 65320 1919 65376
rect 0 65318 1919 65320
rect 0 65288 800 65318
rect 1853 65315 1919 65318
rect 4208 65312 4528 65313
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 14208 65312 14528 65313
rect 14208 65248 14216 65312
rect 14280 65248 14296 65312
rect 14360 65248 14376 65312
rect 14440 65248 14456 65312
rect 14520 65248 14528 65312
rect 14208 65247 14528 65248
rect 24208 65312 24528 65313
rect 24208 65248 24216 65312
rect 24280 65248 24296 65312
rect 24360 65248 24376 65312
rect 24440 65248 24456 65312
rect 24520 65248 24528 65312
rect 24208 65247 24528 65248
rect 34208 65312 34528 65313
rect 34208 65248 34216 65312
rect 34280 65248 34296 65312
rect 34360 65248 34376 65312
rect 34440 65248 34456 65312
rect 34520 65248 34528 65312
rect 34208 65247 34528 65248
rect 44208 65312 44528 65313
rect 44208 65248 44216 65312
rect 44280 65248 44296 65312
rect 44360 65248 44376 65312
rect 44440 65248 44456 65312
rect 44520 65248 44528 65312
rect 44208 65247 44528 65248
rect 54208 65312 54528 65313
rect 54208 65248 54216 65312
rect 54280 65248 54296 65312
rect 54360 65248 54376 65312
rect 54440 65248 54456 65312
rect 54520 65248 54528 65312
rect 54208 65247 54528 65248
rect 64208 65312 64528 65313
rect 64208 65248 64216 65312
rect 64280 65248 64296 65312
rect 64360 65248 64376 65312
rect 64440 65248 64456 65312
rect 64520 65248 64528 65312
rect 69200 65288 70000 65408
rect 64208 65247 64528 65248
rect 9208 64768 9528 64769
rect 9208 64704 9216 64768
rect 9280 64704 9296 64768
rect 9360 64704 9376 64768
rect 9440 64704 9456 64768
rect 9520 64704 9528 64768
rect 9208 64703 9528 64704
rect 19208 64768 19528 64769
rect 19208 64704 19216 64768
rect 19280 64704 19296 64768
rect 19360 64704 19376 64768
rect 19440 64704 19456 64768
rect 19520 64704 19528 64768
rect 19208 64703 19528 64704
rect 29208 64768 29528 64769
rect 29208 64704 29216 64768
rect 29280 64704 29296 64768
rect 29360 64704 29376 64768
rect 29440 64704 29456 64768
rect 29520 64704 29528 64768
rect 29208 64703 29528 64704
rect 39208 64768 39528 64769
rect 39208 64704 39216 64768
rect 39280 64704 39296 64768
rect 39360 64704 39376 64768
rect 39440 64704 39456 64768
rect 39520 64704 39528 64768
rect 39208 64703 39528 64704
rect 49208 64768 49528 64769
rect 49208 64704 49216 64768
rect 49280 64704 49296 64768
rect 49360 64704 49376 64768
rect 49440 64704 49456 64768
rect 49520 64704 49528 64768
rect 49208 64703 49528 64704
rect 59208 64768 59528 64769
rect 59208 64704 59216 64768
rect 59280 64704 59296 64768
rect 59360 64704 59376 64768
rect 59440 64704 59456 64768
rect 59520 64704 59528 64768
rect 59208 64703 59528 64704
rect 4208 64224 4528 64225
rect 0 64064 800 64184
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 14208 64224 14528 64225
rect 14208 64160 14216 64224
rect 14280 64160 14296 64224
rect 14360 64160 14376 64224
rect 14440 64160 14456 64224
rect 14520 64160 14528 64224
rect 14208 64159 14528 64160
rect 24208 64224 24528 64225
rect 24208 64160 24216 64224
rect 24280 64160 24296 64224
rect 24360 64160 24376 64224
rect 24440 64160 24456 64224
rect 24520 64160 24528 64224
rect 24208 64159 24528 64160
rect 34208 64224 34528 64225
rect 34208 64160 34216 64224
rect 34280 64160 34296 64224
rect 34360 64160 34376 64224
rect 34440 64160 34456 64224
rect 34520 64160 34528 64224
rect 34208 64159 34528 64160
rect 44208 64224 44528 64225
rect 44208 64160 44216 64224
rect 44280 64160 44296 64224
rect 44360 64160 44376 64224
rect 44440 64160 44456 64224
rect 44520 64160 44528 64224
rect 44208 64159 44528 64160
rect 54208 64224 54528 64225
rect 54208 64160 54216 64224
rect 54280 64160 54296 64224
rect 54360 64160 54376 64224
rect 54440 64160 54456 64224
rect 54520 64160 54528 64224
rect 54208 64159 54528 64160
rect 64208 64224 64528 64225
rect 64208 64160 64216 64224
rect 64280 64160 64296 64224
rect 64360 64160 64376 64224
rect 64440 64160 64456 64224
rect 64520 64160 64528 64224
rect 64208 64159 64528 64160
rect 68093 64018 68159 64021
rect 69200 64018 70000 64048
rect 68093 64016 70000 64018
rect 68093 63960 68098 64016
rect 68154 63960 70000 64016
rect 68093 63958 70000 63960
rect 68093 63955 68159 63958
rect 69200 63928 70000 63958
rect 9208 63680 9528 63681
rect 9208 63616 9216 63680
rect 9280 63616 9296 63680
rect 9360 63616 9376 63680
rect 9440 63616 9456 63680
rect 9520 63616 9528 63680
rect 9208 63615 9528 63616
rect 19208 63680 19528 63681
rect 19208 63616 19216 63680
rect 19280 63616 19296 63680
rect 19360 63616 19376 63680
rect 19440 63616 19456 63680
rect 19520 63616 19528 63680
rect 19208 63615 19528 63616
rect 29208 63680 29528 63681
rect 29208 63616 29216 63680
rect 29280 63616 29296 63680
rect 29360 63616 29376 63680
rect 29440 63616 29456 63680
rect 29520 63616 29528 63680
rect 29208 63615 29528 63616
rect 39208 63680 39528 63681
rect 39208 63616 39216 63680
rect 39280 63616 39296 63680
rect 39360 63616 39376 63680
rect 39440 63616 39456 63680
rect 39520 63616 39528 63680
rect 39208 63615 39528 63616
rect 49208 63680 49528 63681
rect 49208 63616 49216 63680
rect 49280 63616 49296 63680
rect 49360 63616 49376 63680
rect 49440 63616 49456 63680
rect 49520 63616 49528 63680
rect 49208 63615 49528 63616
rect 59208 63680 59528 63681
rect 59208 63616 59216 63680
rect 59280 63616 59296 63680
rect 59360 63616 59376 63680
rect 59440 63616 59456 63680
rect 59520 63616 59528 63680
rect 59208 63615 59528 63616
rect 4208 63136 4528 63137
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 14208 63136 14528 63137
rect 14208 63072 14216 63136
rect 14280 63072 14296 63136
rect 14360 63072 14376 63136
rect 14440 63072 14456 63136
rect 14520 63072 14528 63136
rect 14208 63071 14528 63072
rect 24208 63136 24528 63137
rect 24208 63072 24216 63136
rect 24280 63072 24296 63136
rect 24360 63072 24376 63136
rect 24440 63072 24456 63136
rect 24520 63072 24528 63136
rect 24208 63071 24528 63072
rect 34208 63136 34528 63137
rect 34208 63072 34216 63136
rect 34280 63072 34296 63136
rect 34360 63072 34376 63136
rect 34440 63072 34456 63136
rect 34520 63072 34528 63136
rect 34208 63071 34528 63072
rect 44208 63136 44528 63137
rect 44208 63072 44216 63136
rect 44280 63072 44296 63136
rect 44360 63072 44376 63136
rect 44440 63072 44456 63136
rect 44520 63072 44528 63136
rect 44208 63071 44528 63072
rect 54208 63136 54528 63137
rect 54208 63072 54216 63136
rect 54280 63072 54296 63136
rect 54360 63072 54376 63136
rect 54440 63072 54456 63136
rect 54520 63072 54528 63136
rect 54208 63071 54528 63072
rect 64208 63136 64528 63137
rect 64208 63072 64216 63136
rect 64280 63072 64296 63136
rect 64360 63072 64376 63136
rect 64440 63072 64456 63136
rect 64520 63072 64528 63136
rect 64208 63071 64528 63072
rect 0 62794 800 62824
rect 1577 62794 1643 62797
rect 0 62792 1643 62794
rect 0 62736 1582 62792
rect 1638 62736 1643 62792
rect 0 62734 1643 62736
rect 0 62704 800 62734
rect 1577 62731 1643 62734
rect 68093 62658 68159 62661
rect 69200 62658 70000 62688
rect 68093 62656 70000 62658
rect 68093 62600 68098 62656
rect 68154 62600 70000 62656
rect 68093 62598 70000 62600
rect 68093 62595 68159 62598
rect 9208 62592 9528 62593
rect 9208 62528 9216 62592
rect 9280 62528 9296 62592
rect 9360 62528 9376 62592
rect 9440 62528 9456 62592
rect 9520 62528 9528 62592
rect 9208 62527 9528 62528
rect 19208 62592 19528 62593
rect 19208 62528 19216 62592
rect 19280 62528 19296 62592
rect 19360 62528 19376 62592
rect 19440 62528 19456 62592
rect 19520 62528 19528 62592
rect 19208 62527 19528 62528
rect 29208 62592 29528 62593
rect 29208 62528 29216 62592
rect 29280 62528 29296 62592
rect 29360 62528 29376 62592
rect 29440 62528 29456 62592
rect 29520 62528 29528 62592
rect 29208 62527 29528 62528
rect 39208 62592 39528 62593
rect 39208 62528 39216 62592
rect 39280 62528 39296 62592
rect 39360 62528 39376 62592
rect 39440 62528 39456 62592
rect 39520 62528 39528 62592
rect 39208 62527 39528 62528
rect 49208 62592 49528 62593
rect 49208 62528 49216 62592
rect 49280 62528 49296 62592
rect 49360 62528 49376 62592
rect 49440 62528 49456 62592
rect 49520 62528 49528 62592
rect 49208 62527 49528 62528
rect 59208 62592 59528 62593
rect 59208 62528 59216 62592
rect 59280 62528 59296 62592
rect 59360 62528 59376 62592
rect 59440 62528 59456 62592
rect 59520 62528 59528 62592
rect 69200 62568 70000 62598
rect 59208 62527 59528 62528
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 14208 62048 14528 62049
rect 14208 61984 14216 62048
rect 14280 61984 14296 62048
rect 14360 61984 14376 62048
rect 14440 61984 14456 62048
rect 14520 61984 14528 62048
rect 14208 61983 14528 61984
rect 24208 62048 24528 62049
rect 24208 61984 24216 62048
rect 24280 61984 24296 62048
rect 24360 61984 24376 62048
rect 24440 61984 24456 62048
rect 24520 61984 24528 62048
rect 24208 61983 24528 61984
rect 34208 62048 34528 62049
rect 34208 61984 34216 62048
rect 34280 61984 34296 62048
rect 34360 61984 34376 62048
rect 34440 61984 34456 62048
rect 34520 61984 34528 62048
rect 34208 61983 34528 61984
rect 44208 62048 44528 62049
rect 44208 61984 44216 62048
rect 44280 61984 44296 62048
rect 44360 61984 44376 62048
rect 44440 61984 44456 62048
rect 44520 61984 44528 62048
rect 44208 61983 44528 61984
rect 54208 62048 54528 62049
rect 54208 61984 54216 62048
rect 54280 61984 54296 62048
rect 54360 61984 54376 62048
rect 54440 61984 54456 62048
rect 54520 61984 54528 62048
rect 54208 61983 54528 61984
rect 64208 62048 64528 62049
rect 64208 61984 64216 62048
rect 64280 61984 64296 62048
rect 64360 61984 64376 62048
rect 64440 61984 64456 62048
rect 64520 61984 64528 62048
rect 64208 61983 64528 61984
rect 0 61570 800 61600
rect 1853 61570 1919 61573
rect 0 61568 1919 61570
rect 0 61512 1858 61568
rect 1914 61512 1919 61568
rect 0 61510 1919 61512
rect 0 61480 800 61510
rect 1853 61507 1919 61510
rect 9208 61504 9528 61505
rect 9208 61440 9216 61504
rect 9280 61440 9296 61504
rect 9360 61440 9376 61504
rect 9440 61440 9456 61504
rect 9520 61440 9528 61504
rect 9208 61439 9528 61440
rect 19208 61504 19528 61505
rect 19208 61440 19216 61504
rect 19280 61440 19296 61504
rect 19360 61440 19376 61504
rect 19440 61440 19456 61504
rect 19520 61440 19528 61504
rect 19208 61439 19528 61440
rect 29208 61504 29528 61505
rect 29208 61440 29216 61504
rect 29280 61440 29296 61504
rect 29360 61440 29376 61504
rect 29440 61440 29456 61504
rect 29520 61440 29528 61504
rect 29208 61439 29528 61440
rect 39208 61504 39528 61505
rect 39208 61440 39216 61504
rect 39280 61440 39296 61504
rect 39360 61440 39376 61504
rect 39440 61440 39456 61504
rect 39520 61440 39528 61504
rect 39208 61439 39528 61440
rect 49208 61504 49528 61505
rect 49208 61440 49216 61504
rect 49280 61440 49296 61504
rect 49360 61440 49376 61504
rect 49440 61440 49456 61504
rect 49520 61440 49528 61504
rect 49208 61439 49528 61440
rect 59208 61504 59528 61505
rect 59208 61440 59216 61504
rect 59280 61440 59296 61504
rect 59360 61440 59376 61504
rect 59440 61440 59456 61504
rect 59520 61440 59528 61504
rect 59208 61439 59528 61440
rect 68093 61298 68159 61301
rect 69200 61298 70000 61328
rect 68093 61296 70000 61298
rect 68093 61240 68098 61296
rect 68154 61240 70000 61296
rect 68093 61238 70000 61240
rect 68093 61235 68159 61238
rect 69200 61208 70000 61238
rect 4208 60960 4528 60961
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 14208 60960 14528 60961
rect 14208 60896 14216 60960
rect 14280 60896 14296 60960
rect 14360 60896 14376 60960
rect 14440 60896 14456 60960
rect 14520 60896 14528 60960
rect 14208 60895 14528 60896
rect 24208 60960 24528 60961
rect 24208 60896 24216 60960
rect 24280 60896 24296 60960
rect 24360 60896 24376 60960
rect 24440 60896 24456 60960
rect 24520 60896 24528 60960
rect 24208 60895 24528 60896
rect 34208 60960 34528 60961
rect 34208 60896 34216 60960
rect 34280 60896 34296 60960
rect 34360 60896 34376 60960
rect 34440 60896 34456 60960
rect 34520 60896 34528 60960
rect 34208 60895 34528 60896
rect 44208 60960 44528 60961
rect 44208 60896 44216 60960
rect 44280 60896 44296 60960
rect 44360 60896 44376 60960
rect 44440 60896 44456 60960
rect 44520 60896 44528 60960
rect 44208 60895 44528 60896
rect 54208 60960 54528 60961
rect 54208 60896 54216 60960
rect 54280 60896 54296 60960
rect 54360 60896 54376 60960
rect 54440 60896 54456 60960
rect 54520 60896 54528 60960
rect 54208 60895 54528 60896
rect 64208 60960 64528 60961
rect 64208 60896 64216 60960
rect 64280 60896 64296 60960
rect 64360 60896 64376 60960
rect 64440 60896 64456 60960
rect 64520 60896 64528 60960
rect 64208 60895 64528 60896
rect 9208 60416 9528 60417
rect 9208 60352 9216 60416
rect 9280 60352 9296 60416
rect 9360 60352 9376 60416
rect 9440 60352 9456 60416
rect 9520 60352 9528 60416
rect 9208 60351 9528 60352
rect 19208 60416 19528 60417
rect 19208 60352 19216 60416
rect 19280 60352 19296 60416
rect 19360 60352 19376 60416
rect 19440 60352 19456 60416
rect 19520 60352 19528 60416
rect 19208 60351 19528 60352
rect 29208 60416 29528 60417
rect 29208 60352 29216 60416
rect 29280 60352 29296 60416
rect 29360 60352 29376 60416
rect 29440 60352 29456 60416
rect 29520 60352 29528 60416
rect 29208 60351 29528 60352
rect 39208 60416 39528 60417
rect 39208 60352 39216 60416
rect 39280 60352 39296 60416
rect 39360 60352 39376 60416
rect 39440 60352 39456 60416
rect 39520 60352 39528 60416
rect 39208 60351 39528 60352
rect 49208 60416 49528 60417
rect 49208 60352 49216 60416
rect 49280 60352 49296 60416
rect 49360 60352 49376 60416
rect 49440 60352 49456 60416
rect 49520 60352 49528 60416
rect 49208 60351 49528 60352
rect 59208 60416 59528 60417
rect 59208 60352 59216 60416
rect 59280 60352 59296 60416
rect 59360 60352 59376 60416
rect 59440 60352 59456 60416
rect 59520 60352 59528 60416
rect 59208 60351 59528 60352
rect 0 60210 800 60240
rect 1761 60210 1827 60213
rect 0 60208 1827 60210
rect 0 60152 1766 60208
rect 1822 60152 1827 60208
rect 0 60150 1827 60152
rect 0 60120 800 60150
rect 1761 60147 1827 60150
rect 69200 59984 70000 60104
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 14208 59872 14528 59873
rect 14208 59808 14216 59872
rect 14280 59808 14296 59872
rect 14360 59808 14376 59872
rect 14440 59808 14456 59872
rect 14520 59808 14528 59872
rect 14208 59807 14528 59808
rect 24208 59872 24528 59873
rect 24208 59808 24216 59872
rect 24280 59808 24296 59872
rect 24360 59808 24376 59872
rect 24440 59808 24456 59872
rect 24520 59808 24528 59872
rect 24208 59807 24528 59808
rect 34208 59872 34528 59873
rect 34208 59808 34216 59872
rect 34280 59808 34296 59872
rect 34360 59808 34376 59872
rect 34440 59808 34456 59872
rect 34520 59808 34528 59872
rect 34208 59807 34528 59808
rect 44208 59872 44528 59873
rect 44208 59808 44216 59872
rect 44280 59808 44296 59872
rect 44360 59808 44376 59872
rect 44440 59808 44456 59872
rect 44520 59808 44528 59872
rect 44208 59807 44528 59808
rect 54208 59872 54528 59873
rect 54208 59808 54216 59872
rect 54280 59808 54296 59872
rect 54360 59808 54376 59872
rect 54440 59808 54456 59872
rect 54520 59808 54528 59872
rect 54208 59807 54528 59808
rect 64208 59872 64528 59873
rect 64208 59808 64216 59872
rect 64280 59808 64296 59872
rect 64360 59808 64376 59872
rect 64440 59808 64456 59872
rect 64520 59808 64528 59872
rect 64208 59807 64528 59808
rect 9208 59328 9528 59329
rect 9208 59264 9216 59328
rect 9280 59264 9296 59328
rect 9360 59264 9376 59328
rect 9440 59264 9456 59328
rect 9520 59264 9528 59328
rect 9208 59263 9528 59264
rect 19208 59328 19528 59329
rect 19208 59264 19216 59328
rect 19280 59264 19296 59328
rect 19360 59264 19376 59328
rect 19440 59264 19456 59328
rect 19520 59264 19528 59328
rect 19208 59263 19528 59264
rect 29208 59328 29528 59329
rect 29208 59264 29216 59328
rect 29280 59264 29296 59328
rect 29360 59264 29376 59328
rect 29440 59264 29456 59328
rect 29520 59264 29528 59328
rect 29208 59263 29528 59264
rect 39208 59328 39528 59329
rect 39208 59264 39216 59328
rect 39280 59264 39296 59328
rect 39360 59264 39376 59328
rect 39440 59264 39456 59328
rect 39520 59264 39528 59328
rect 39208 59263 39528 59264
rect 49208 59328 49528 59329
rect 49208 59264 49216 59328
rect 49280 59264 49296 59328
rect 49360 59264 49376 59328
rect 49440 59264 49456 59328
rect 49520 59264 49528 59328
rect 49208 59263 49528 59264
rect 59208 59328 59528 59329
rect 59208 59264 59216 59328
rect 59280 59264 59296 59328
rect 59360 59264 59376 59328
rect 59440 59264 59456 59328
rect 59520 59264 59528 59328
rect 59208 59263 59528 59264
rect 0 58896 800 59016
rect 4208 58784 4528 58785
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 14208 58784 14528 58785
rect 14208 58720 14216 58784
rect 14280 58720 14296 58784
rect 14360 58720 14376 58784
rect 14440 58720 14456 58784
rect 14520 58720 14528 58784
rect 14208 58719 14528 58720
rect 24208 58784 24528 58785
rect 24208 58720 24216 58784
rect 24280 58720 24296 58784
rect 24360 58720 24376 58784
rect 24440 58720 24456 58784
rect 24520 58720 24528 58784
rect 24208 58719 24528 58720
rect 34208 58784 34528 58785
rect 34208 58720 34216 58784
rect 34280 58720 34296 58784
rect 34360 58720 34376 58784
rect 34440 58720 34456 58784
rect 34520 58720 34528 58784
rect 34208 58719 34528 58720
rect 44208 58784 44528 58785
rect 44208 58720 44216 58784
rect 44280 58720 44296 58784
rect 44360 58720 44376 58784
rect 44440 58720 44456 58784
rect 44520 58720 44528 58784
rect 44208 58719 44528 58720
rect 54208 58784 54528 58785
rect 54208 58720 54216 58784
rect 54280 58720 54296 58784
rect 54360 58720 54376 58784
rect 54440 58720 54456 58784
rect 54520 58720 54528 58784
rect 54208 58719 54528 58720
rect 64208 58784 64528 58785
rect 64208 58720 64216 58784
rect 64280 58720 64296 58784
rect 64360 58720 64376 58784
rect 64440 58720 64456 58784
rect 64520 58720 64528 58784
rect 64208 58719 64528 58720
rect 68093 58714 68159 58717
rect 69200 58714 70000 58744
rect 68093 58712 70000 58714
rect 68093 58656 68098 58712
rect 68154 58656 70000 58712
rect 68093 58654 70000 58656
rect 68093 58651 68159 58654
rect 69200 58624 70000 58654
rect 9208 58240 9528 58241
rect 9208 58176 9216 58240
rect 9280 58176 9296 58240
rect 9360 58176 9376 58240
rect 9440 58176 9456 58240
rect 9520 58176 9528 58240
rect 9208 58175 9528 58176
rect 19208 58240 19528 58241
rect 19208 58176 19216 58240
rect 19280 58176 19296 58240
rect 19360 58176 19376 58240
rect 19440 58176 19456 58240
rect 19520 58176 19528 58240
rect 19208 58175 19528 58176
rect 29208 58240 29528 58241
rect 29208 58176 29216 58240
rect 29280 58176 29296 58240
rect 29360 58176 29376 58240
rect 29440 58176 29456 58240
rect 29520 58176 29528 58240
rect 29208 58175 29528 58176
rect 39208 58240 39528 58241
rect 39208 58176 39216 58240
rect 39280 58176 39296 58240
rect 39360 58176 39376 58240
rect 39440 58176 39456 58240
rect 39520 58176 39528 58240
rect 39208 58175 39528 58176
rect 49208 58240 49528 58241
rect 49208 58176 49216 58240
rect 49280 58176 49296 58240
rect 49360 58176 49376 58240
rect 49440 58176 49456 58240
rect 49520 58176 49528 58240
rect 49208 58175 49528 58176
rect 59208 58240 59528 58241
rect 59208 58176 59216 58240
rect 59280 58176 59296 58240
rect 59360 58176 59376 58240
rect 59440 58176 59456 58240
rect 59520 58176 59528 58240
rect 59208 58175 59528 58176
rect 4208 57696 4528 57697
rect 0 57626 800 57656
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 14208 57696 14528 57697
rect 14208 57632 14216 57696
rect 14280 57632 14296 57696
rect 14360 57632 14376 57696
rect 14440 57632 14456 57696
rect 14520 57632 14528 57696
rect 14208 57631 14528 57632
rect 24208 57696 24528 57697
rect 24208 57632 24216 57696
rect 24280 57632 24296 57696
rect 24360 57632 24376 57696
rect 24440 57632 24456 57696
rect 24520 57632 24528 57696
rect 24208 57631 24528 57632
rect 34208 57696 34528 57697
rect 34208 57632 34216 57696
rect 34280 57632 34296 57696
rect 34360 57632 34376 57696
rect 34440 57632 34456 57696
rect 34520 57632 34528 57696
rect 34208 57631 34528 57632
rect 44208 57696 44528 57697
rect 44208 57632 44216 57696
rect 44280 57632 44296 57696
rect 44360 57632 44376 57696
rect 44440 57632 44456 57696
rect 44520 57632 44528 57696
rect 44208 57631 44528 57632
rect 54208 57696 54528 57697
rect 54208 57632 54216 57696
rect 54280 57632 54296 57696
rect 54360 57632 54376 57696
rect 54440 57632 54456 57696
rect 54520 57632 54528 57696
rect 54208 57631 54528 57632
rect 64208 57696 64528 57697
rect 64208 57632 64216 57696
rect 64280 57632 64296 57696
rect 64360 57632 64376 57696
rect 64440 57632 64456 57696
rect 64520 57632 64528 57696
rect 64208 57631 64528 57632
rect 1577 57626 1643 57629
rect 0 57624 1643 57626
rect 0 57568 1582 57624
rect 1638 57568 1643 57624
rect 0 57566 1643 57568
rect 0 57536 800 57566
rect 1577 57563 1643 57566
rect 68093 57354 68159 57357
rect 69200 57354 70000 57384
rect 68093 57352 70000 57354
rect 68093 57296 68098 57352
rect 68154 57296 70000 57352
rect 68093 57294 70000 57296
rect 68093 57291 68159 57294
rect 69200 57264 70000 57294
rect 9208 57152 9528 57153
rect 9208 57088 9216 57152
rect 9280 57088 9296 57152
rect 9360 57088 9376 57152
rect 9440 57088 9456 57152
rect 9520 57088 9528 57152
rect 9208 57087 9528 57088
rect 19208 57152 19528 57153
rect 19208 57088 19216 57152
rect 19280 57088 19296 57152
rect 19360 57088 19376 57152
rect 19440 57088 19456 57152
rect 19520 57088 19528 57152
rect 19208 57087 19528 57088
rect 29208 57152 29528 57153
rect 29208 57088 29216 57152
rect 29280 57088 29296 57152
rect 29360 57088 29376 57152
rect 29440 57088 29456 57152
rect 29520 57088 29528 57152
rect 29208 57087 29528 57088
rect 39208 57152 39528 57153
rect 39208 57088 39216 57152
rect 39280 57088 39296 57152
rect 39360 57088 39376 57152
rect 39440 57088 39456 57152
rect 39520 57088 39528 57152
rect 39208 57087 39528 57088
rect 49208 57152 49528 57153
rect 49208 57088 49216 57152
rect 49280 57088 49296 57152
rect 49360 57088 49376 57152
rect 49440 57088 49456 57152
rect 49520 57088 49528 57152
rect 49208 57087 49528 57088
rect 59208 57152 59528 57153
rect 59208 57088 59216 57152
rect 59280 57088 59296 57152
rect 59360 57088 59376 57152
rect 59440 57088 59456 57152
rect 59520 57088 59528 57152
rect 59208 57087 59528 57088
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 14208 56608 14528 56609
rect 14208 56544 14216 56608
rect 14280 56544 14296 56608
rect 14360 56544 14376 56608
rect 14440 56544 14456 56608
rect 14520 56544 14528 56608
rect 14208 56543 14528 56544
rect 24208 56608 24528 56609
rect 24208 56544 24216 56608
rect 24280 56544 24296 56608
rect 24360 56544 24376 56608
rect 24440 56544 24456 56608
rect 24520 56544 24528 56608
rect 24208 56543 24528 56544
rect 34208 56608 34528 56609
rect 34208 56544 34216 56608
rect 34280 56544 34296 56608
rect 34360 56544 34376 56608
rect 34440 56544 34456 56608
rect 34520 56544 34528 56608
rect 34208 56543 34528 56544
rect 44208 56608 44528 56609
rect 44208 56544 44216 56608
rect 44280 56544 44296 56608
rect 44360 56544 44376 56608
rect 44440 56544 44456 56608
rect 44520 56544 44528 56608
rect 44208 56543 44528 56544
rect 54208 56608 54528 56609
rect 54208 56544 54216 56608
rect 54280 56544 54296 56608
rect 54360 56544 54376 56608
rect 54440 56544 54456 56608
rect 54520 56544 54528 56608
rect 54208 56543 54528 56544
rect 64208 56608 64528 56609
rect 64208 56544 64216 56608
rect 64280 56544 64296 56608
rect 64360 56544 64376 56608
rect 64440 56544 64456 56608
rect 64520 56544 64528 56608
rect 64208 56543 64528 56544
rect 0 56402 800 56432
rect 1761 56402 1827 56405
rect 0 56400 1827 56402
rect 0 56344 1766 56400
rect 1822 56344 1827 56400
rect 0 56342 1827 56344
rect 0 56312 800 56342
rect 1761 56339 1827 56342
rect 68093 56130 68159 56133
rect 69200 56130 70000 56160
rect 68093 56128 70000 56130
rect 68093 56072 68098 56128
rect 68154 56072 70000 56128
rect 68093 56070 70000 56072
rect 68093 56067 68159 56070
rect 9208 56064 9528 56065
rect 9208 56000 9216 56064
rect 9280 56000 9296 56064
rect 9360 56000 9376 56064
rect 9440 56000 9456 56064
rect 9520 56000 9528 56064
rect 9208 55999 9528 56000
rect 19208 56064 19528 56065
rect 19208 56000 19216 56064
rect 19280 56000 19296 56064
rect 19360 56000 19376 56064
rect 19440 56000 19456 56064
rect 19520 56000 19528 56064
rect 19208 55999 19528 56000
rect 29208 56064 29528 56065
rect 29208 56000 29216 56064
rect 29280 56000 29296 56064
rect 29360 56000 29376 56064
rect 29440 56000 29456 56064
rect 29520 56000 29528 56064
rect 29208 55999 29528 56000
rect 39208 56064 39528 56065
rect 39208 56000 39216 56064
rect 39280 56000 39296 56064
rect 39360 56000 39376 56064
rect 39440 56000 39456 56064
rect 39520 56000 39528 56064
rect 39208 55999 39528 56000
rect 49208 56064 49528 56065
rect 49208 56000 49216 56064
rect 49280 56000 49296 56064
rect 49360 56000 49376 56064
rect 49440 56000 49456 56064
rect 49520 56000 49528 56064
rect 49208 55999 49528 56000
rect 59208 56064 59528 56065
rect 59208 56000 59216 56064
rect 59280 56000 59296 56064
rect 59360 56000 59376 56064
rect 59440 56000 59456 56064
rect 59520 56000 59528 56064
rect 69200 56040 70000 56070
rect 59208 55999 59528 56000
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 14208 55520 14528 55521
rect 14208 55456 14216 55520
rect 14280 55456 14296 55520
rect 14360 55456 14376 55520
rect 14440 55456 14456 55520
rect 14520 55456 14528 55520
rect 14208 55455 14528 55456
rect 24208 55520 24528 55521
rect 24208 55456 24216 55520
rect 24280 55456 24296 55520
rect 24360 55456 24376 55520
rect 24440 55456 24456 55520
rect 24520 55456 24528 55520
rect 24208 55455 24528 55456
rect 34208 55520 34528 55521
rect 34208 55456 34216 55520
rect 34280 55456 34296 55520
rect 34360 55456 34376 55520
rect 34440 55456 34456 55520
rect 34520 55456 34528 55520
rect 34208 55455 34528 55456
rect 44208 55520 44528 55521
rect 44208 55456 44216 55520
rect 44280 55456 44296 55520
rect 44360 55456 44376 55520
rect 44440 55456 44456 55520
rect 44520 55456 44528 55520
rect 44208 55455 44528 55456
rect 54208 55520 54528 55521
rect 54208 55456 54216 55520
rect 54280 55456 54296 55520
rect 54360 55456 54376 55520
rect 54440 55456 54456 55520
rect 54520 55456 54528 55520
rect 54208 55455 54528 55456
rect 64208 55520 64528 55521
rect 64208 55456 64216 55520
rect 64280 55456 64296 55520
rect 64360 55456 64376 55520
rect 64440 55456 64456 55520
rect 64520 55456 64528 55520
rect 64208 55455 64528 55456
rect 0 55042 800 55072
rect 1853 55042 1919 55045
rect 0 55040 1919 55042
rect 0 54984 1858 55040
rect 1914 54984 1919 55040
rect 0 54982 1919 54984
rect 0 54952 800 54982
rect 1853 54979 1919 54982
rect 9208 54976 9528 54977
rect 9208 54912 9216 54976
rect 9280 54912 9296 54976
rect 9360 54912 9376 54976
rect 9440 54912 9456 54976
rect 9520 54912 9528 54976
rect 9208 54911 9528 54912
rect 19208 54976 19528 54977
rect 19208 54912 19216 54976
rect 19280 54912 19296 54976
rect 19360 54912 19376 54976
rect 19440 54912 19456 54976
rect 19520 54912 19528 54976
rect 19208 54911 19528 54912
rect 29208 54976 29528 54977
rect 29208 54912 29216 54976
rect 29280 54912 29296 54976
rect 29360 54912 29376 54976
rect 29440 54912 29456 54976
rect 29520 54912 29528 54976
rect 29208 54911 29528 54912
rect 39208 54976 39528 54977
rect 39208 54912 39216 54976
rect 39280 54912 39296 54976
rect 39360 54912 39376 54976
rect 39440 54912 39456 54976
rect 39520 54912 39528 54976
rect 39208 54911 39528 54912
rect 49208 54976 49528 54977
rect 49208 54912 49216 54976
rect 49280 54912 49296 54976
rect 49360 54912 49376 54976
rect 49440 54912 49456 54976
rect 49520 54912 49528 54976
rect 49208 54911 49528 54912
rect 59208 54976 59528 54977
rect 59208 54912 59216 54976
rect 59280 54912 59296 54976
rect 59360 54912 59376 54976
rect 59440 54912 59456 54976
rect 59520 54912 59528 54976
rect 59208 54911 59528 54912
rect 69200 54680 70000 54800
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 14208 54432 14528 54433
rect 14208 54368 14216 54432
rect 14280 54368 14296 54432
rect 14360 54368 14376 54432
rect 14440 54368 14456 54432
rect 14520 54368 14528 54432
rect 14208 54367 14528 54368
rect 24208 54432 24528 54433
rect 24208 54368 24216 54432
rect 24280 54368 24296 54432
rect 24360 54368 24376 54432
rect 24440 54368 24456 54432
rect 24520 54368 24528 54432
rect 24208 54367 24528 54368
rect 34208 54432 34528 54433
rect 34208 54368 34216 54432
rect 34280 54368 34296 54432
rect 34360 54368 34376 54432
rect 34440 54368 34456 54432
rect 34520 54368 34528 54432
rect 34208 54367 34528 54368
rect 44208 54432 44528 54433
rect 44208 54368 44216 54432
rect 44280 54368 44296 54432
rect 44360 54368 44376 54432
rect 44440 54368 44456 54432
rect 44520 54368 44528 54432
rect 44208 54367 44528 54368
rect 54208 54432 54528 54433
rect 54208 54368 54216 54432
rect 54280 54368 54296 54432
rect 54360 54368 54376 54432
rect 54440 54368 54456 54432
rect 54520 54368 54528 54432
rect 54208 54367 54528 54368
rect 64208 54432 64528 54433
rect 64208 54368 64216 54432
rect 64280 54368 64296 54432
rect 64360 54368 64376 54432
rect 64440 54368 64456 54432
rect 64520 54368 64528 54432
rect 64208 54367 64528 54368
rect 9208 53888 9528 53889
rect 0 53728 800 53848
rect 9208 53824 9216 53888
rect 9280 53824 9296 53888
rect 9360 53824 9376 53888
rect 9440 53824 9456 53888
rect 9520 53824 9528 53888
rect 9208 53823 9528 53824
rect 19208 53888 19528 53889
rect 19208 53824 19216 53888
rect 19280 53824 19296 53888
rect 19360 53824 19376 53888
rect 19440 53824 19456 53888
rect 19520 53824 19528 53888
rect 19208 53823 19528 53824
rect 29208 53888 29528 53889
rect 29208 53824 29216 53888
rect 29280 53824 29296 53888
rect 29360 53824 29376 53888
rect 29440 53824 29456 53888
rect 29520 53824 29528 53888
rect 29208 53823 29528 53824
rect 39208 53888 39528 53889
rect 39208 53824 39216 53888
rect 39280 53824 39296 53888
rect 39360 53824 39376 53888
rect 39440 53824 39456 53888
rect 39520 53824 39528 53888
rect 39208 53823 39528 53824
rect 49208 53888 49528 53889
rect 49208 53824 49216 53888
rect 49280 53824 49296 53888
rect 49360 53824 49376 53888
rect 49440 53824 49456 53888
rect 49520 53824 49528 53888
rect 49208 53823 49528 53824
rect 59208 53888 59528 53889
rect 59208 53824 59216 53888
rect 59280 53824 59296 53888
rect 59360 53824 59376 53888
rect 59440 53824 59456 53888
rect 59520 53824 59528 53888
rect 59208 53823 59528 53824
rect 68093 53410 68159 53413
rect 69200 53410 70000 53440
rect 68093 53408 70000 53410
rect 68093 53352 68098 53408
rect 68154 53352 70000 53408
rect 68093 53350 70000 53352
rect 68093 53347 68159 53350
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 14208 53344 14528 53345
rect 14208 53280 14216 53344
rect 14280 53280 14296 53344
rect 14360 53280 14376 53344
rect 14440 53280 14456 53344
rect 14520 53280 14528 53344
rect 14208 53279 14528 53280
rect 24208 53344 24528 53345
rect 24208 53280 24216 53344
rect 24280 53280 24296 53344
rect 24360 53280 24376 53344
rect 24440 53280 24456 53344
rect 24520 53280 24528 53344
rect 24208 53279 24528 53280
rect 34208 53344 34528 53345
rect 34208 53280 34216 53344
rect 34280 53280 34296 53344
rect 34360 53280 34376 53344
rect 34440 53280 34456 53344
rect 34520 53280 34528 53344
rect 34208 53279 34528 53280
rect 44208 53344 44528 53345
rect 44208 53280 44216 53344
rect 44280 53280 44296 53344
rect 44360 53280 44376 53344
rect 44440 53280 44456 53344
rect 44520 53280 44528 53344
rect 44208 53279 44528 53280
rect 54208 53344 54528 53345
rect 54208 53280 54216 53344
rect 54280 53280 54296 53344
rect 54360 53280 54376 53344
rect 54440 53280 54456 53344
rect 54520 53280 54528 53344
rect 54208 53279 54528 53280
rect 64208 53344 64528 53345
rect 64208 53280 64216 53344
rect 64280 53280 64296 53344
rect 64360 53280 64376 53344
rect 64440 53280 64456 53344
rect 64520 53280 64528 53344
rect 69200 53320 70000 53350
rect 64208 53279 64528 53280
rect 9208 52800 9528 52801
rect 9208 52736 9216 52800
rect 9280 52736 9296 52800
rect 9360 52736 9376 52800
rect 9440 52736 9456 52800
rect 9520 52736 9528 52800
rect 9208 52735 9528 52736
rect 19208 52800 19528 52801
rect 19208 52736 19216 52800
rect 19280 52736 19296 52800
rect 19360 52736 19376 52800
rect 19440 52736 19456 52800
rect 19520 52736 19528 52800
rect 19208 52735 19528 52736
rect 29208 52800 29528 52801
rect 29208 52736 29216 52800
rect 29280 52736 29296 52800
rect 29360 52736 29376 52800
rect 29440 52736 29456 52800
rect 29520 52736 29528 52800
rect 29208 52735 29528 52736
rect 39208 52800 39528 52801
rect 39208 52736 39216 52800
rect 39280 52736 39296 52800
rect 39360 52736 39376 52800
rect 39440 52736 39456 52800
rect 39520 52736 39528 52800
rect 39208 52735 39528 52736
rect 49208 52800 49528 52801
rect 49208 52736 49216 52800
rect 49280 52736 49296 52800
rect 49360 52736 49376 52800
rect 49440 52736 49456 52800
rect 49520 52736 49528 52800
rect 49208 52735 49528 52736
rect 59208 52800 59528 52801
rect 59208 52736 59216 52800
rect 59280 52736 59296 52800
rect 59360 52736 59376 52800
rect 59440 52736 59456 52800
rect 59520 52736 59528 52800
rect 59208 52735 59528 52736
rect 0 52458 800 52488
rect 1577 52458 1643 52461
rect 0 52456 1643 52458
rect 0 52400 1582 52456
rect 1638 52400 1643 52456
rect 0 52398 1643 52400
rect 0 52368 800 52398
rect 1577 52395 1643 52398
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 14208 52256 14528 52257
rect 14208 52192 14216 52256
rect 14280 52192 14296 52256
rect 14360 52192 14376 52256
rect 14440 52192 14456 52256
rect 14520 52192 14528 52256
rect 14208 52191 14528 52192
rect 24208 52256 24528 52257
rect 24208 52192 24216 52256
rect 24280 52192 24296 52256
rect 24360 52192 24376 52256
rect 24440 52192 24456 52256
rect 24520 52192 24528 52256
rect 24208 52191 24528 52192
rect 34208 52256 34528 52257
rect 34208 52192 34216 52256
rect 34280 52192 34296 52256
rect 34360 52192 34376 52256
rect 34440 52192 34456 52256
rect 34520 52192 34528 52256
rect 34208 52191 34528 52192
rect 44208 52256 44528 52257
rect 44208 52192 44216 52256
rect 44280 52192 44296 52256
rect 44360 52192 44376 52256
rect 44440 52192 44456 52256
rect 44520 52192 44528 52256
rect 44208 52191 44528 52192
rect 54208 52256 54528 52257
rect 54208 52192 54216 52256
rect 54280 52192 54296 52256
rect 54360 52192 54376 52256
rect 54440 52192 54456 52256
rect 54520 52192 54528 52256
rect 54208 52191 54528 52192
rect 64208 52256 64528 52257
rect 64208 52192 64216 52256
rect 64280 52192 64296 52256
rect 64360 52192 64376 52256
rect 64440 52192 64456 52256
rect 64520 52192 64528 52256
rect 64208 52191 64528 52192
rect 68093 52050 68159 52053
rect 69200 52050 70000 52080
rect 68093 52048 70000 52050
rect 68093 51992 68098 52048
rect 68154 51992 70000 52048
rect 68093 51990 70000 51992
rect 68093 51987 68159 51990
rect 69200 51960 70000 51990
rect 9208 51712 9528 51713
rect 9208 51648 9216 51712
rect 9280 51648 9296 51712
rect 9360 51648 9376 51712
rect 9440 51648 9456 51712
rect 9520 51648 9528 51712
rect 9208 51647 9528 51648
rect 19208 51712 19528 51713
rect 19208 51648 19216 51712
rect 19280 51648 19296 51712
rect 19360 51648 19376 51712
rect 19440 51648 19456 51712
rect 19520 51648 19528 51712
rect 19208 51647 19528 51648
rect 29208 51712 29528 51713
rect 29208 51648 29216 51712
rect 29280 51648 29296 51712
rect 29360 51648 29376 51712
rect 29440 51648 29456 51712
rect 29520 51648 29528 51712
rect 29208 51647 29528 51648
rect 39208 51712 39528 51713
rect 39208 51648 39216 51712
rect 39280 51648 39296 51712
rect 39360 51648 39376 51712
rect 39440 51648 39456 51712
rect 39520 51648 39528 51712
rect 39208 51647 39528 51648
rect 49208 51712 49528 51713
rect 49208 51648 49216 51712
rect 49280 51648 49296 51712
rect 49360 51648 49376 51712
rect 49440 51648 49456 51712
rect 49520 51648 49528 51712
rect 49208 51647 49528 51648
rect 59208 51712 59528 51713
rect 59208 51648 59216 51712
rect 59280 51648 59296 51712
rect 59360 51648 59376 51712
rect 59440 51648 59456 51712
rect 59520 51648 59528 51712
rect 59208 51647 59528 51648
rect 4208 51168 4528 51169
rect 0 51098 800 51128
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 14208 51168 14528 51169
rect 14208 51104 14216 51168
rect 14280 51104 14296 51168
rect 14360 51104 14376 51168
rect 14440 51104 14456 51168
rect 14520 51104 14528 51168
rect 14208 51103 14528 51104
rect 24208 51168 24528 51169
rect 24208 51104 24216 51168
rect 24280 51104 24296 51168
rect 24360 51104 24376 51168
rect 24440 51104 24456 51168
rect 24520 51104 24528 51168
rect 24208 51103 24528 51104
rect 34208 51168 34528 51169
rect 34208 51104 34216 51168
rect 34280 51104 34296 51168
rect 34360 51104 34376 51168
rect 34440 51104 34456 51168
rect 34520 51104 34528 51168
rect 34208 51103 34528 51104
rect 44208 51168 44528 51169
rect 44208 51104 44216 51168
rect 44280 51104 44296 51168
rect 44360 51104 44376 51168
rect 44440 51104 44456 51168
rect 44520 51104 44528 51168
rect 44208 51103 44528 51104
rect 54208 51168 54528 51169
rect 54208 51104 54216 51168
rect 54280 51104 54296 51168
rect 54360 51104 54376 51168
rect 54440 51104 54456 51168
rect 54520 51104 54528 51168
rect 54208 51103 54528 51104
rect 64208 51168 64528 51169
rect 64208 51104 64216 51168
rect 64280 51104 64296 51168
rect 64360 51104 64376 51168
rect 64440 51104 64456 51168
rect 64520 51104 64528 51168
rect 64208 51103 64528 51104
rect 1853 51098 1919 51101
rect 0 51096 1919 51098
rect 0 51040 1858 51096
rect 1914 51040 1919 51096
rect 0 51038 1919 51040
rect 0 51008 800 51038
rect 1853 51035 1919 51038
rect 68093 50826 68159 50829
rect 69200 50826 70000 50856
rect 68093 50824 70000 50826
rect 68093 50768 68098 50824
rect 68154 50768 70000 50824
rect 68093 50766 70000 50768
rect 68093 50763 68159 50766
rect 69200 50736 70000 50766
rect 9208 50624 9528 50625
rect 9208 50560 9216 50624
rect 9280 50560 9296 50624
rect 9360 50560 9376 50624
rect 9440 50560 9456 50624
rect 9520 50560 9528 50624
rect 9208 50559 9528 50560
rect 19208 50624 19528 50625
rect 19208 50560 19216 50624
rect 19280 50560 19296 50624
rect 19360 50560 19376 50624
rect 19440 50560 19456 50624
rect 19520 50560 19528 50624
rect 19208 50559 19528 50560
rect 29208 50624 29528 50625
rect 29208 50560 29216 50624
rect 29280 50560 29296 50624
rect 29360 50560 29376 50624
rect 29440 50560 29456 50624
rect 29520 50560 29528 50624
rect 29208 50559 29528 50560
rect 39208 50624 39528 50625
rect 39208 50560 39216 50624
rect 39280 50560 39296 50624
rect 39360 50560 39376 50624
rect 39440 50560 39456 50624
rect 39520 50560 39528 50624
rect 39208 50559 39528 50560
rect 49208 50624 49528 50625
rect 49208 50560 49216 50624
rect 49280 50560 49296 50624
rect 49360 50560 49376 50624
rect 49440 50560 49456 50624
rect 49520 50560 49528 50624
rect 49208 50559 49528 50560
rect 59208 50624 59528 50625
rect 59208 50560 59216 50624
rect 59280 50560 59296 50624
rect 59360 50560 59376 50624
rect 59440 50560 59456 50624
rect 59520 50560 59528 50624
rect 59208 50559 59528 50560
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 14208 50080 14528 50081
rect 14208 50016 14216 50080
rect 14280 50016 14296 50080
rect 14360 50016 14376 50080
rect 14440 50016 14456 50080
rect 14520 50016 14528 50080
rect 14208 50015 14528 50016
rect 24208 50080 24528 50081
rect 24208 50016 24216 50080
rect 24280 50016 24296 50080
rect 24360 50016 24376 50080
rect 24440 50016 24456 50080
rect 24520 50016 24528 50080
rect 24208 50015 24528 50016
rect 34208 50080 34528 50081
rect 34208 50016 34216 50080
rect 34280 50016 34296 50080
rect 34360 50016 34376 50080
rect 34440 50016 34456 50080
rect 34520 50016 34528 50080
rect 34208 50015 34528 50016
rect 44208 50080 44528 50081
rect 44208 50016 44216 50080
rect 44280 50016 44296 50080
rect 44360 50016 44376 50080
rect 44440 50016 44456 50080
rect 44520 50016 44528 50080
rect 44208 50015 44528 50016
rect 54208 50080 54528 50081
rect 54208 50016 54216 50080
rect 54280 50016 54296 50080
rect 54360 50016 54376 50080
rect 54440 50016 54456 50080
rect 54520 50016 54528 50080
rect 54208 50015 54528 50016
rect 64208 50080 64528 50081
rect 64208 50016 64216 50080
rect 64280 50016 64296 50080
rect 64360 50016 64376 50080
rect 64440 50016 64456 50080
rect 64520 50016 64528 50080
rect 64208 50015 64528 50016
rect 0 49874 800 49904
rect 1761 49874 1827 49877
rect 0 49872 1827 49874
rect 0 49816 1766 49872
rect 1822 49816 1827 49872
rect 0 49814 1827 49816
rect 0 49784 800 49814
rect 1761 49811 1827 49814
rect 9208 49536 9528 49537
rect 9208 49472 9216 49536
rect 9280 49472 9296 49536
rect 9360 49472 9376 49536
rect 9440 49472 9456 49536
rect 9520 49472 9528 49536
rect 9208 49471 9528 49472
rect 19208 49536 19528 49537
rect 19208 49472 19216 49536
rect 19280 49472 19296 49536
rect 19360 49472 19376 49536
rect 19440 49472 19456 49536
rect 19520 49472 19528 49536
rect 19208 49471 19528 49472
rect 29208 49536 29528 49537
rect 29208 49472 29216 49536
rect 29280 49472 29296 49536
rect 29360 49472 29376 49536
rect 29440 49472 29456 49536
rect 29520 49472 29528 49536
rect 29208 49471 29528 49472
rect 39208 49536 39528 49537
rect 39208 49472 39216 49536
rect 39280 49472 39296 49536
rect 39360 49472 39376 49536
rect 39440 49472 39456 49536
rect 39520 49472 39528 49536
rect 39208 49471 39528 49472
rect 49208 49536 49528 49537
rect 49208 49472 49216 49536
rect 49280 49472 49296 49536
rect 49360 49472 49376 49536
rect 49440 49472 49456 49536
rect 49520 49472 49528 49536
rect 49208 49471 49528 49472
rect 59208 49536 59528 49537
rect 59208 49472 59216 49536
rect 59280 49472 59296 49536
rect 59360 49472 59376 49536
rect 59440 49472 59456 49536
rect 59520 49472 59528 49536
rect 59208 49471 59528 49472
rect 69200 49376 70000 49496
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 14208 48992 14528 48993
rect 14208 48928 14216 48992
rect 14280 48928 14296 48992
rect 14360 48928 14376 48992
rect 14440 48928 14456 48992
rect 14520 48928 14528 48992
rect 14208 48927 14528 48928
rect 24208 48992 24528 48993
rect 24208 48928 24216 48992
rect 24280 48928 24296 48992
rect 24360 48928 24376 48992
rect 24440 48928 24456 48992
rect 24520 48928 24528 48992
rect 24208 48927 24528 48928
rect 34208 48992 34528 48993
rect 34208 48928 34216 48992
rect 34280 48928 34296 48992
rect 34360 48928 34376 48992
rect 34440 48928 34456 48992
rect 34520 48928 34528 48992
rect 34208 48927 34528 48928
rect 44208 48992 44528 48993
rect 44208 48928 44216 48992
rect 44280 48928 44296 48992
rect 44360 48928 44376 48992
rect 44440 48928 44456 48992
rect 44520 48928 44528 48992
rect 44208 48927 44528 48928
rect 54208 48992 54528 48993
rect 54208 48928 54216 48992
rect 54280 48928 54296 48992
rect 54360 48928 54376 48992
rect 54440 48928 54456 48992
rect 54520 48928 54528 48992
rect 54208 48927 54528 48928
rect 64208 48992 64528 48993
rect 64208 48928 64216 48992
rect 64280 48928 64296 48992
rect 64360 48928 64376 48992
rect 64440 48928 64456 48992
rect 64520 48928 64528 48992
rect 64208 48927 64528 48928
rect 0 48424 800 48544
rect 9208 48448 9528 48449
rect 9208 48384 9216 48448
rect 9280 48384 9296 48448
rect 9360 48384 9376 48448
rect 9440 48384 9456 48448
rect 9520 48384 9528 48448
rect 9208 48383 9528 48384
rect 19208 48448 19528 48449
rect 19208 48384 19216 48448
rect 19280 48384 19296 48448
rect 19360 48384 19376 48448
rect 19440 48384 19456 48448
rect 19520 48384 19528 48448
rect 19208 48383 19528 48384
rect 29208 48448 29528 48449
rect 29208 48384 29216 48448
rect 29280 48384 29296 48448
rect 29360 48384 29376 48448
rect 29440 48384 29456 48448
rect 29520 48384 29528 48448
rect 29208 48383 29528 48384
rect 39208 48448 39528 48449
rect 39208 48384 39216 48448
rect 39280 48384 39296 48448
rect 39360 48384 39376 48448
rect 39440 48384 39456 48448
rect 39520 48384 39528 48448
rect 39208 48383 39528 48384
rect 49208 48448 49528 48449
rect 49208 48384 49216 48448
rect 49280 48384 49296 48448
rect 49360 48384 49376 48448
rect 49440 48384 49456 48448
rect 49520 48384 49528 48448
rect 49208 48383 49528 48384
rect 59208 48448 59528 48449
rect 59208 48384 59216 48448
rect 59280 48384 59296 48448
rect 59360 48384 59376 48448
rect 59440 48384 59456 48448
rect 59520 48384 59528 48448
rect 59208 48383 59528 48384
rect 68093 48106 68159 48109
rect 69200 48106 70000 48136
rect 68093 48104 70000 48106
rect 68093 48048 68098 48104
rect 68154 48048 70000 48104
rect 68093 48046 70000 48048
rect 68093 48043 68159 48046
rect 69200 48016 70000 48046
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 14208 47904 14528 47905
rect 14208 47840 14216 47904
rect 14280 47840 14296 47904
rect 14360 47840 14376 47904
rect 14440 47840 14456 47904
rect 14520 47840 14528 47904
rect 14208 47839 14528 47840
rect 24208 47904 24528 47905
rect 24208 47840 24216 47904
rect 24280 47840 24296 47904
rect 24360 47840 24376 47904
rect 24440 47840 24456 47904
rect 24520 47840 24528 47904
rect 24208 47839 24528 47840
rect 34208 47904 34528 47905
rect 34208 47840 34216 47904
rect 34280 47840 34296 47904
rect 34360 47840 34376 47904
rect 34440 47840 34456 47904
rect 34520 47840 34528 47904
rect 34208 47839 34528 47840
rect 44208 47904 44528 47905
rect 44208 47840 44216 47904
rect 44280 47840 44296 47904
rect 44360 47840 44376 47904
rect 44440 47840 44456 47904
rect 44520 47840 44528 47904
rect 44208 47839 44528 47840
rect 54208 47904 54528 47905
rect 54208 47840 54216 47904
rect 54280 47840 54296 47904
rect 54360 47840 54376 47904
rect 54440 47840 54456 47904
rect 54520 47840 54528 47904
rect 54208 47839 54528 47840
rect 64208 47904 64528 47905
rect 64208 47840 64216 47904
rect 64280 47840 64296 47904
rect 64360 47840 64376 47904
rect 64440 47840 64456 47904
rect 64520 47840 64528 47904
rect 64208 47839 64528 47840
rect 9208 47360 9528 47361
rect 0 47290 800 47320
rect 9208 47296 9216 47360
rect 9280 47296 9296 47360
rect 9360 47296 9376 47360
rect 9440 47296 9456 47360
rect 9520 47296 9528 47360
rect 9208 47295 9528 47296
rect 19208 47360 19528 47361
rect 19208 47296 19216 47360
rect 19280 47296 19296 47360
rect 19360 47296 19376 47360
rect 19440 47296 19456 47360
rect 19520 47296 19528 47360
rect 19208 47295 19528 47296
rect 29208 47360 29528 47361
rect 29208 47296 29216 47360
rect 29280 47296 29296 47360
rect 29360 47296 29376 47360
rect 29440 47296 29456 47360
rect 29520 47296 29528 47360
rect 29208 47295 29528 47296
rect 39208 47360 39528 47361
rect 39208 47296 39216 47360
rect 39280 47296 39296 47360
rect 39360 47296 39376 47360
rect 39440 47296 39456 47360
rect 39520 47296 39528 47360
rect 39208 47295 39528 47296
rect 49208 47360 49528 47361
rect 49208 47296 49216 47360
rect 49280 47296 49296 47360
rect 49360 47296 49376 47360
rect 49440 47296 49456 47360
rect 49520 47296 49528 47360
rect 49208 47295 49528 47296
rect 59208 47360 59528 47361
rect 59208 47296 59216 47360
rect 59280 47296 59296 47360
rect 59360 47296 59376 47360
rect 59440 47296 59456 47360
rect 59520 47296 59528 47360
rect 59208 47295 59528 47296
rect 1853 47290 1919 47293
rect 0 47288 1919 47290
rect 0 47232 1858 47288
rect 1914 47232 1919 47288
rect 0 47230 1919 47232
rect 0 47200 800 47230
rect 1853 47227 1919 47230
rect 68093 46882 68159 46885
rect 69200 46882 70000 46912
rect 68093 46880 70000 46882
rect 68093 46824 68098 46880
rect 68154 46824 70000 46880
rect 68093 46822 70000 46824
rect 68093 46819 68159 46822
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 14208 46816 14528 46817
rect 14208 46752 14216 46816
rect 14280 46752 14296 46816
rect 14360 46752 14376 46816
rect 14440 46752 14456 46816
rect 14520 46752 14528 46816
rect 14208 46751 14528 46752
rect 24208 46816 24528 46817
rect 24208 46752 24216 46816
rect 24280 46752 24296 46816
rect 24360 46752 24376 46816
rect 24440 46752 24456 46816
rect 24520 46752 24528 46816
rect 24208 46751 24528 46752
rect 34208 46816 34528 46817
rect 34208 46752 34216 46816
rect 34280 46752 34296 46816
rect 34360 46752 34376 46816
rect 34440 46752 34456 46816
rect 34520 46752 34528 46816
rect 34208 46751 34528 46752
rect 44208 46816 44528 46817
rect 44208 46752 44216 46816
rect 44280 46752 44296 46816
rect 44360 46752 44376 46816
rect 44440 46752 44456 46816
rect 44520 46752 44528 46816
rect 44208 46751 44528 46752
rect 54208 46816 54528 46817
rect 54208 46752 54216 46816
rect 54280 46752 54296 46816
rect 54360 46752 54376 46816
rect 54440 46752 54456 46816
rect 54520 46752 54528 46816
rect 54208 46751 54528 46752
rect 64208 46816 64528 46817
rect 64208 46752 64216 46816
rect 64280 46752 64296 46816
rect 64360 46752 64376 46816
rect 64440 46752 64456 46816
rect 64520 46752 64528 46816
rect 69200 46792 70000 46822
rect 64208 46751 64528 46752
rect 9208 46272 9528 46273
rect 9208 46208 9216 46272
rect 9280 46208 9296 46272
rect 9360 46208 9376 46272
rect 9440 46208 9456 46272
rect 9520 46208 9528 46272
rect 9208 46207 9528 46208
rect 19208 46272 19528 46273
rect 19208 46208 19216 46272
rect 19280 46208 19296 46272
rect 19360 46208 19376 46272
rect 19440 46208 19456 46272
rect 19520 46208 19528 46272
rect 19208 46207 19528 46208
rect 29208 46272 29528 46273
rect 29208 46208 29216 46272
rect 29280 46208 29296 46272
rect 29360 46208 29376 46272
rect 29440 46208 29456 46272
rect 29520 46208 29528 46272
rect 29208 46207 29528 46208
rect 39208 46272 39528 46273
rect 39208 46208 39216 46272
rect 39280 46208 39296 46272
rect 39360 46208 39376 46272
rect 39440 46208 39456 46272
rect 39520 46208 39528 46272
rect 39208 46207 39528 46208
rect 49208 46272 49528 46273
rect 49208 46208 49216 46272
rect 49280 46208 49296 46272
rect 49360 46208 49376 46272
rect 49440 46208 49456 46272
rect 49520 46208 49528 46272
rect 49208 46207 49528 46208
rect 59208 46272 59528 46273
rect 59208 46208 59216 46272
rect 59280 46208 59296 46272
rect 59360 46208 59376 46272
rect 59440 46208 59456 46272
rect 59520 46208 59528 46272
rect 59208 46207 59528 46208
rect 0 45930 800 45960
rect 1761 45930 1827 45933
rect 0 45928 1827 45930
rect 0 45872 1766 45928
rect 1822 45872 1827 45928
rect 0 45870 1827 45872
rect 0 45840 800 45870
rect 1761 45867 1827 45870
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 14208 45728 14528 45729
rect 14208 45664 14216 45728
rect 14280 45664 14296 45728
rect 14360 45664 14376 45728
rect 14440 45664 14456 45728
rect 14520 45664 14528 45728
rect 14208 45663 14528 45664
rect 24208 45728 24528 45729
rect 24208 45664 24216 45728
rect 24280 45664 24296 45728
rect 24360 45664 24376 45728
rect 24440 45664 24456 45728
rect 24520 45664 24528 45728
rect 24208 45663 24528 45664
rect 34208 45728 34528 45729
rect 34208 45664 34216 45728
rect 34280 45664 34296 45728
rect 34360 45664 34376 45728
rect 34440 45664 34456 45728
rect 34520 45664 34528 45728
rect 34208 45663 34528 45664
rect 44208 45728 44528 45729
rect 44208 45664 44216 45728
rect 44280 45664 44296 45728
rect 44360 45664 44376 45728
rect 44440 45664 44456 45728
rect 44520 45664 44528 45728
rect 44208 45663 44528 45664
rect 54208 45728 54528 45729
rect 54208 45664 54216 45728
rect 54280 45664 54296 45728
rect 54360 45664 54376 45728
rect 54440 45664 54456 45728
rect 54520 45664 54528 45728
rect 54208 45663 54528 45664
rect 64208 45728 64528 45729
rect 64208 45664 64216 45728
rect 64280 45664 64296 45728
rect 64360 45664 64376 45728
rect 64440 45664 64456 45728
rect 64520 45664 64528 45728
rect 64208 45663 64528 45664
rect 68093 45522 68159 45525
rect 69200 45522 70000 45552
rect 68093 45520 70000 45522
rect 68093 45464 68098 45520
rect 68154 45464 70000 45520
rect 68093 45462 70000 45464
rect 68093 45459 68159 45462
rect 69200 45432 70000 45462
rect 9208 45184 9528 45185
rect 9208 45120 9216 45184
rect 9280 45120 9296 45184
rect 9360 45120 9376 45184
rect 9440 45120 9456 45184
rect 9520 45120 9528 45184
rect 9208 45119 9528 45120
rect 19208 45184 19528 45185
rect 19208 45120 19216 45184
rect 19280 45120 19296 45184
rect 19360 45120 19376 45184
rect 19440 45120 19456 45184
rect 19520 45120 19528 45184
rect 19208 45119 19528 45120
rect 29208 45184 29528 45185
rect 29208 45120 29216 45184
rect 29280 45120 29296 45184
rect 29360 45120 29376 45184
rect 29440 45120 29456 45184
rect 29520 45120 29528 45184
rect 29208 45119 29528 45120
rect 39208 45184 39528 45185
rect 39208 45120 39216 45184
rect 39280 45120 39296 45184
rect 39360 45120 39376 45184
rect 39440 45120 39456 45184
rect 39520 45120 39528 45184
rect 39208 45119 39528 45120
rect 49208 45184 49528 45185
rect 49208 45120 49216 45184
rect 49280 45120 49296 45184
rect 49360 45120 49376 45184
rect 49440 45120 49456 45184
rect 49520 45120 49528 45184
rect 49208 45119 49528 45120
rect 59208 45184 59528 45185
rect 59208 45120 59216 45184
rect 59280 45120 59296 45184
rect 59360 45120 59376 45184
rect 59440 45120 59456 45184
rect 59520 45120 59528 45184
rect 59208 45119 59528 45120
rect 0 44706 800 44736
rect 1853 44706 1919 44709
rect 0 44704 1919 44706
rect 0 44648 1858 44704
rect 1914 44648 1919 44704
rect 0 44646 1919 44648
rect 0 44616 800 44646
rect 1853 44643 1919 44646
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 14208 44640 14528 44641
rect 14208 44576 14216 44640
rect 14280 44576 14296 44640
rect 14360 44576 14376 44640
rect 14440 44576 14456 44640
rect 14520 44576 14528 44640
rect 14208 44575 14528 44576
rect 24208 44640 24528 44641
rect 24208 44576 24216 44640
rect 24280 44576 24296 44640
rect 24360 44576 24376 44640
rect 24440 44576 24456 44640
rect 24520 44576 24528 44640
rect 24208 44575 24528 44576
rect 34208 44640 34528 44641
rect 34208 44576 34216 44640
rect 34280 44576 34296 44640
rect 34360 44576 34376 44640
rect 34440 44576 34456 44640
rect 34520 44576 34528 44640
rect 34208 44575 34528 44576
rect 44208 44640 44528 44641
rect 44208 44576 44216 44640
rect 44280 44576 44296 44640
rect 44360 44576 44376 44640
rect 44440 44576 44456 44640
rect 44520 44576 44528 44640
rect 44208 44575 44528 44576
rect 54208 44640 54528 44641
rect 54208 44576 54216 44640
rect 54280 44576 54296 44640
rect 54360 44576 54376 44640
rect 54440 44576 54456 44640
rect 54520 44576 54528 44640
rect 54208 44575 54528 44576
rect 64208 44640 64528 44641
rect 64208 44576 64216 44640
rect 64280 44576 64296 44640
rect 64360 44576 64376 44640
rect 64440 44576 64456 44640
rect 64520 44576 64528 44640
rect 64208 44575 64528 44576
rect 9208 44096 9528 44097
rect 9208 44032 9216 44096
rect 9280 44032 9296 44096
rect 9360 44032 9376 44096
rect 9440 44032 9456 44096
rect 9520 44032 9528 44096
rect 9208 44031 9528 44032
rect 19208 44096 19528 44097
rect 19208 44032 19216 44096
rect 19280 44032 19296 44096
rect 19360 44032 19376 44096
rect 19440 44032 19456 44096
rect 19520 44032 19528 44096
rect 19208 44031 19528 44032
rect 29208 44096 29528 44097
rect 29208 44032 29216 44096
rect 29280 44032 29296 44096
rect 29360 44032 29376 44096
rect 29440 44032 29456 44096
rect 29520 44032 29528 44096
rect 29208 44031 29528 44032
rect 39208 44096 39528 44097
rect 39208 44032 39216 44096
rect 39280 44032 39296 44096
rect 39360 44032 39376 44096
rect 39440 44032 39456 44096
rect 39520 44032 39528 44096
rect 39208 44031 39528 44032
rect 49208 44096 49528 44097
rect 49208 44032 49216 44096
rect 49280 44032 49296 44096
rect 49360 44032 49376 44096
rect 49440 44032 49456 44096
rect 49520 44032 49528 44096
rect 49208 44031 49528 44032
rect 59208 44096 59528 44097
rect 59208 44032 59216 44096
rect 59280 44032 59296 44096
rect 59360 44032 59376 44096
rect 59440 44032 59456 44096
rect 59520 44032 59528 44096
rect 69200 44072 70000 44192
rect 59208 44031 59528 44032
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 14208 43552 14528 43553
rect 14208 43488 14216 43552
rect 14280 43488 14296 43552
rect 14360 43488 14376 43552
rect 14440 43488 14456 43552
rect 14520 43488 14528 43552
rect 14208 43487 14528 43488
rect 24208 43552 24528 43553
rect 24208 43488 24216 43552
rect 24280 43488 24296 43552
rect 24360 43488 24376 43552
rect 24440 43488 24456 43552
rect 24520 43488 24528 43552
rect 24208 43487 24528 43488
rect 34208 43552 34528 43553
rect 34208 43488 34216 43552
rect 34280 43488 34296 43552
rect 34360 43488 34376 43552
rect 34440 43488 34456 43552
rect 34520 43488 34528 43552
rect 34208 43487 34528 43488
rect 44208 43552 44528 43553
rect 44208 43488 44216 43552
rect 44280 43488 44296 43552
rect 44360 43488 44376 43552
rect 44440 43488 44456 43552
rect 44520 43488 44528 43552
rect 44208 43487 44528 43488
rect 54208 43552 54528 43553
rect 54208 43488 54216 43552
rect 54280 43488 54296 43552
rect 54360 43488 54376 43552
rect 54440 43488 54456 43552
rect 54520 43488 54528 43552
rect 54208 43487 54528 43488
rect 64208 43552 64528 43553
rect 64208 43488 64216 43552
rect 64280 43488 64296 43552
rect 64360 43488 64376 43552
rect 64440 43488 64456 43552
rect 64520 43488 64528 43552
rect 64208 43487 64528 43488
rect 0 43256 800 43376
rect 9208 43008 9528 43009
rect 9208 42944 9216 43008
rect 9280 42944 9296 43008
rect 9360 42944 9376 43008
rect 9440 42944 9456 43008
rect 9520 42944 9528 43008
rect 9208 42943 9528 42944
rect 19208 43008 19528 43009
rect 19208 42944 19216 43008
rect 19280 42944 19296 43008
rect 19360 42944 19376 43008
rect 19440 42944 19456 43008
rect 19520 42944 19528 43008
rect 19208 42943 19528 42944
rect 29208 43008 29528 43009
rect 29208 42944 29216 43008
rect 29280 42944 29296 43008
rect 29360 42944 29376 43008
rect 29440 42944 29456 43008
rect 29520 42944 29528 43008
rect 29208 42943 29528 42944
rect 39208 43008 39528 43009
rect 39208 42944 39216 43008
rect 39280 42944 39296 43008
rect 39360 42944 39376 43008
rect 39440 42944 39456 43008
rect 39520 42944 39528 43008
rect 39208 42943 39528 42944
rect 49208 43008 49528 43009
rect 49208 42944 49216 43008
rect 49280 42944 49296 43008
rect 49360 42944 49376 43008
rect 49440 42944 49456 43008
rect 49520 42944 49528 43008
rect 49208 42943 49528 42944
rect 59208 43008 59528 43009
rect 59208 42944 59216 43008
rect 59280 42944 59296 43008
rect 59360 42944 59376 43008
rect 59440 42944 59456 43008
rect 59520 42944 59528 43008
rect 59208 42943 59528 42944
rect 68093 42802 68159 42805
rect 69200 42802 70000 42832
rect 68093 42800 70000 42802
rect 68093 42744 68098 42800
rect 68154 42744 70000 42800
rect 68093 42742 70000 42744
rect 68093 42739 68159 42742
rect 69200 42712 70000 42742
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 14208 42464 14528 42465
rect 14208 42400 14216 42464
rect 14280 42400 14296 42464
rect 14360 42400 14376 42464
rect 14440 42400 14456 42464
rect 14520 42400 14528 42464
rect 14208 42399 14528 42400
rect 24208 42464 24528 42465
rect 24208 42400 24216 42464
rect 24280 42400 24296 42464
rect 24360 42400 24376 42464
rect 24440 42400 24456 42464
rect 24520 42400 24528 42464
rect 24208 42399 24528 42400
rect 34208 42464 34528 42465
rect 34208 42400 34216 42464
rect 34280 42400 34296 42464
rect 34360 42400 34376 42464
rect 34440 42400 34456 42464
rect 34520 42400 34528 42464
rect 34208 42399 34528 42400
rect 44208 42464 44528 42465
rect 44208 42400 44216 42464
rect 44280 42400 44296 42464
rect 44360 42400 44376 42464
rect 44440 42400 44456 42464
rect 44520 42400 44528 42464
rect 44208 42399 44528 42400
rect 54208 42464 54528 42465
rect 54208 42400 54216 42464
rect 54280 42400 54296 42464
rect 54360 42400 54376 42464
rect 54440 42400 54456 42464
rect 54520 42400 54528 42464
rect 54208 42399 54528 42400
rect 64208 42464 64528 42465
rect 64208 42400 64216 42464
rect 64280 42400 64296 42464
rect 64360 42400 64376 42464
rect 64440 42400 64456 42464
rect 64520 42400 64528 42464
rect 64208 42399 64528 42400
rect 0 42122 800 42152
rect 1577 42122 1643 42125
rect 0 42120 1643 42122
rect 0 42064 1582 42120
rect 1638 42064 1643 42120
rect 0 42062 1643 42064
rect 0 42032 800 42062
rect 1577 42059 1643 42062
rect 9208 41920 9528 41921
rect 9208 41856 9216 41920
rect 9280 41856 9296 41920
rect 9360 41856 9376 41920
rect 9440 41856 9456 41920
rect 9520 41856 9528 41920
rect 9208 41855 9528 41856
rect 19208 41920 19528 41921
rect 19208 41856 19216 41920
rect 19280 41856 19296 41920
rect 19360 41856 19376 41920
rect 19440 41856 19456 41920
rect 19520 41856 19528 41920
rect 19208 41855 19528 41856
rect 29208 41920 29528 41921
rect 29208 41856 29216 41920
rect 29280 41856 29296 41920
rect 29360 41856 29376 41920
rect 29440 41856 29456 41920
rect 29520 41856 29528 41920
rect 29208 41855 29528 41856
rect 39208 41920 39528 41921
rect 39208 41856 39216 41920
rect 39280 41856 39296 41920
rect 39360 41856 39376 41920
rect 39440 41856 39456 41920
rect 39520 41856 39528 41920
rect 39208 41855 39528 41856
rect 49208 41920 49528 41921
rect 49208 41856 49216 41920
rect 49280 41856 49296 41920
rect 49360 41856 49376 41920
rect 49440 41856 49456 41920
rect 49520 41856 49528 41920
rect 49208 41855 49528 41856
rect 59208 41920 59528 41921
rect 59208 41856 59216 41920
rect 59280 41856 59296 41920
rect 59360 41856 59376 41920
rect 59440 41856 59456 41920
rect 59520 41856 59528 41920
rect 59208 41855 59528 41856
rect 68093 41578 68159 41581
rect 69200 41578 70000 41608
rect 68093 41576 70000 41578
rect 68093 41520 68098 41576
rect 68154 41520 70000 41576
rect 68093 41518 70000 41520
rect 68093 41515 68159 41518
rect 69200 41488 70000 41518
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 14208 41376 14528 41377
rect 14208 41312 14216 41376
rect 14280 41312 14296 41376
rect 14360 41312 14376 41376
rect 14440 41312 14456 41376
rect 14520 41312 14528 41376
rect 14208 41311 14528 41312
rect 24208 41376 24528 41377
rect 24208 41312 24216 41376
rect 24280 41312 24296 41376
rect 24360 41312 24376 41376
rect 24440 41312 24456 41376
rect 24520 41312 24528 41376
rect 24208 41311 24528 41312
rect 34208 41376 34528 41377
rect 34208 41312 34216 41376
rect 34280 41312 34296 41376
rect 34360 41312 34376 41376
rect 34440 41312 34456 41376
rect 34520 41312 34528 41376
rect 34208 41311 34528 41312
rect 44208 41376 44528 41377
rect 44208 41312 44216 41376
rect 44280 41312 44296 41376
rect 44360 41312 44376 41376
rect 44440 41312 44456 41376
rect 44520 41312 44528 41376
rect 44208 41311 44528 41312
rect 54208 41376 54528 41377
rect 54208 41312 54216 41376
rect 54280 41312 54296 41376
rect 54360 41312 54376 41376
rect 54440 41312 54456 41376
rect 54520 41312 54528 41376
rect 54208 41311 54528 41312
rect 64208 41376 64528 41377
rect 64208 41312 64216 41376
rect 64280 41312 64296 41376
rect 64360 41312 64376 41376
rect 64440 41312 64456 41376
rect 64520 41312 64528 41376
rect 64208 41311 64528 41312
rect 9208 40832 9528 40833
rect 0 40762 800 40792
rect 9208 40768 9216 40832
rect 9280 40768 9296 40832
rect 9360 40768 9376 40832
rect 9440 40768 9456 40832
rect 9520 40768 9528 40832
rect 9208 40767 9528 40768
rect 19208 40832 19528 40833
rect 19208 40768 19216 40832
rect 19280 40768 19296 40832
rect 19360 40768 19376 40832
rect 19440 40768 19456 40832
rect 19520 40768 19528 40832
rect 19208 40767 19528 40768
rect 29208 40832 29528 40833
rect 29208 40768 29216 40832
rect 29280 40768 29296 40832
rect 29360 40768 29376 40832
rect 29440 40768 29456 40832
rect 29520 40768 29528 40832
rect 29208 40767 29528 40768
rect 39208 40832 39528 40833
rect 39208 40768 39216 40832
rect 39280 40768 39296 40832
rect 39360 40768 39376 40832
rect 39440 40768 39456 40832
rect 39520 40768 39528 40832
rect 39208 40767 39528 40768
rect 49208 40832 49528 40833
rect 49208 40768 49216 40832
rect 49280 40768 49296 40832
rect 49360 40768 49376 40832
rect 49440 40768 49456 40832
rect 49520 40768 49528 40832
rect 49208 40767 49528 40768
rect 59208 40832 59528 40833
rect 59208 40768 59216 40832
rect 59280 40768 59296 40832
rect 59360 40768 59376 40832
rect 59440 40768 59456 40832
rect 59520 40768 59528 40832
rect 59208 40767 59528 40768
rect 1853 40762 1919 40765
rect 0 40760 1919 40762
rect 0 40704 1858 40760
rect 1914 40704 1919 40760
rect 0 40702 1919 40704
rect 0 40672 800 40702
rect 1853 40699 1919 40702
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 14208 40288 14528 40289
rect 14208 40224 14216 40288
rect 14280 40224 14296 40288
rect 14360 40224 14376 40288
rect 14440 40224 14456 40288
rect 14520 40224 14528 40288
rect 14208 40223 14528 40224
rect 24208 40288 24528 40289
rect 24208 40224 24216 40288
rect 24280 40224 24296 40288
rect 24360 40224 24376 40288
rect 24440 40224 24456 40288
rect 24520 40224 24528 40288
rect 24208 40223 24528 40224
rect 34208 40288 34528 40289
rect 34208 40224 34216 40288
rect 34280 40224 34296 40288
rect 34360 40224 34376 40288
rect 34440 40224 34456 40288
rect 34520 40224 34528 40288
rect 34208 40223 34528 40224
rect 44208 40288 44528 40289
rect 44208 40224 44216 40288
rect 44280 40224 44296 40288
rect 44360 40224 44376 40288
rect 44440 40224 44456 40288
rect 44520 40224 44528 40288
rect 44208 40223 44528 40224
rect 54208 40288 54528 40289
rect 54208 40224 54216 40288
rect 54280 40224 54296 40288
rect 54360 40224 54376 40288
rect 54440 40224 54456 40288
rect 54520 40224 54528 40288
rect 54208 40223 54528 40224
rect 64208 40288 64528 40289
rect 64208 40224 64216 40288
rect 64280 40224 64296 40288
rect 64360 40224 64376 40288
rect 64440 40224 64456 40288
rect 64520 40224 64528 40288
rect 64208 40223 64528 40224
rect 68093 40218 68159 40221
rect 69200 40218 70000 40248
rect 68093 40216 70000 40218
rect 68093 40160 68098 40216
rect 68154 40160 70000 40216
rect 68093 40158 70000 40160
rect 68093 40155 68159 40158
rect 69200 40128 70000 40158
rect 9208 39744 9528 39745
rect 9208 39680 9216 39744
rect 9280 39680 9296 39744
rect 9360 39680 9376 39744
rect 9440 39680 9456 39744
rect 9520 39680 9528 39744
rect 9208 39679 9528 39680
rect 19208 39744 19528 39745
rect 19208 39680 19216 39744
rect 19280 39680 19296 39744
rect 19360 39680 19376 39744
rect 19440 39680 19456 39744
rect 19520 39680 19528 39744
rect 19208 39679 19528 39680
rect 29208 39744 29528 39745
rect 29208 39680 29216 39744
rect 29280 39680 29296 39744
rect 29360 39680 29376 39744
rect 29440 39680 29456 39744
rect 29520 39680 29528 39744
rect 29208 39679 29528 39680
rect 39208 39744 39528 39745
rect 39208 39680 39216 39744
rect 39280 39680 39296 39744
rect 39360 39680 39376 39744
rect 39440 39680 39456 39744
rect 39520 39680 39528 39744
rect 39208 39679 39528 39680
rect 49208 39744 49528 39745
rect 49208 39680 49216 39744
rect 49280 39680 49296 39744
rect 49360 39680 49376 39744
rect 49440 39680 49456 39744
rect 49520 39680 49528 39744
rect 49208 39679 49528 39680
rect 59208 39744 59528 39745
rect 59208 39680 59216 39744
rect 59280 39680 59296 39744
rect 59360 39680 59376 39744
rect 59440 39680 59456 39744
rect 59520 39680 59528 39744
rect 59208 39679 59528 39680
rect 0 39538 800 39568
rect 1761 39538 1827 39541
rect 0 39536 1827 39538
rect 0 39480 1766 39536
rect 1822 39480 1827 39536
rect 0 39478 1827 39480
rect 0 39448 800 39478
rect 1761 39475 1827 39478
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 14208 39200 14528 39201
rect 14208 39136 14216 39200
rect 14280 39136 14296 39200
rect 14360 39136 14376 39200
rect 14440 39136 14456 39200
rect 14520 39136 14528 39200
rect 14208 39135 14528 39136
rect 24208 39200 24528 39201
rect 24208 39136 24216 39200
rect 24280 39136 24296 39200
rect 24360 39136 24376 39200
rect 24440 39136 24456 39200
rect 24520 39136 24528 39200
rect 24208 39135 24528 39136
rect 34208 39200 34528 39201
rect 34208 39136 34216 39200
rect 34280 39136 34296 39200
rect 34360 39136 34376 39200
rect 34440 39136 34456 39200
rect 34520 39136 34528 39200
rect 34208 39135 34528 39136
rect 44208 39200 44528 39201
rect 44208 39136 44216 39200
rect 44280 39136 44296 39200
rect 44360 39136 44376 39200
rect 44440 39136 44456 39200
rect 44520 39136 44528 39200
rect 44208 39135 44528 39136
rect 54208 39200 54528 39201
rect 54208 39136 54216 39200
rect 54280 39136 54296 39200
rect 54360 39136 54376 39200
rect 54440 39136 54456 39200
rect 54520 39136 54528 39200
rect 54208 39135 54528 39136
rect 64208 39200 64528 39201
rect 64208 39136 64216 39200
rect 64280 39136 64296 39200
rect 64360 39136 64376 39200
rect 64440 39136 64456 39200
rect 64520 39136 64528 39200
rect 64208 39135 64528 39136
rect 69200 38768 70000 38888
rect 9208 38656 9528 38657
rect 9208 38592 9216 38656
rect 9280 38592 9296 38656
rect 9360 38592 9376 38656
rect 9440 38592 9456 38656
rect 9520 38592 9528 38656
rect 9208 38591 9528 38592
rect 19208 38656 19528 38657
rect 19208 38592 19216 38656
rect 19280 38592 19296 38656
rect 19360 38592 19376 38656
rect 19440 38592 19456 38656
rect 19520 38592 19528 38656
rect 19208 38591 19528 38592
rect 29208 38656 29528 38657
rect 29208 38592 29216 38656
rect 29280 38592 29296 38656
rect 29360 38592 29376 38656
rect 29440 38592 29456 38656
rect 29520 38592 29528 38656
rect 29208 38591 29528 38592
rect 39208 38656 39528 38657
rect 39208 38592 39216 38656
rect 39280 38592 39296 38656
rect 39360 38592 39376 38656
rect 39440 38592 39456 38656
rect 39520 38592 39528 38656
rect 39208 38591 39528 38592
rect 49208 38656 49528 38657
rect 49208 38592 49216 38656
rect 49280 38592 49296 38656
rect 49360 38592 49376 38656
rect 49440 38592 49456 38656
rect 49520 38592 49528 38656
rect 49208 38591 49528 38592
rect 59208 38656 59528 38657
rect 59208 38592 59216 38656
rect 59280 38592 59296 38656
rect 59360 38592 59376 38656
rect 59440 38592 59456 38656
rect 59520 38592 59528 38656
rect 59208 38591 59528 38592
rect 0 38088 800 38208
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 14208 38112 14528 38113
rect 14208 38048 14216 38112
rect 14280 38048 14296 38112
rect 14360 38048 14376 38112
rect 14440 38048 14456 38112
rect 14520 38048 14528 38112
rect 14208 38047 14528 38048
rect 24208 38112 24528 38113
rect 24208 38048 24216 38112
rect 24280 38048 24296 38112
rect 24360 38048 24376 38112
rect 24440 38048 24456 38112
rect 24520 38048 24528 38112
rect 24208 38047 24528 38048
rect 34208 38112 34528 38113
rect 34208 38048 34216 38112
rect 34280 38048 34296 38112
rect 34360 38048 34376 38112
rect 34440 38048 34456 38112
rect 34520 38048 34528 38112
rect 34208 38047 34528 38048
rect 44208 38112 44528 38113
rect 44208 38048 44216 38112
rect 44280 38048 44296 38112
rect 44360 38048 44376 38112
rect 44440 38048 44456 38112
rect 44520 38048 44528 38112
rect 44208 38047 44528 38048
rect 54208 38112 54528 38113
rect 54208 38048 54216 38112
rect 54280 38048 54296 38112
rect 54360 38048 54376 38112
rect 54440 38048 54456 38112
rect 54520 38048 54528 38112
rect 54208 38047 54528 38048
rect 64208 38112 64528 38113
rect 64208 38048 64216 38112
rect 64280 38048 64296 38112
rect 64360 38048 64376 38112
rect 64440 38048 64456 38112
rect 64520 38048 64528 38112
rect 64208 38047 64528 38048
rect 68093 37634 68159 37637
rect 69200 37634 70000 37664
rect 68093 37632 70000 37634
rect 68093 37576 68098 37632
rect 68154 37576 70000 37632
rect 68093 37574 70000 37576
rect 68093 37571 68159 37574
rect 9208 37568 9528 37569
rect 9208 37504 9216 37568
rect 9280 37504 9296 37568
rect 9360 37504 9376 37568
rect 9440 37504 9456 37568
rect 9520 37504 9528 37568
rect 9208 37503 9528 37504
rect 19208 37568 19528 37569
rect 19208 37504 19216 37568
rect 19280 37504 19296 37568
rect 19360 37504 19376 37568
rect 19440 37504 19456 37568
rect 19520 37504 19528 37568
rect 19208 37503 19528 37504
rect 29208 37568 29528 37569
rect 29208 37504 29216 37568
rect 29280 37504 29296 37568
rect 29360 37504 29376 37568
rect 29440 37504 29456 37568
rect 29520 37504 29528 37568
rect 29208 37503 29528 37504
rect 39208 37568 39528 37569
rect 39208 37504 39216 37568
rect 39280 37504 39296 37568
rect 39360 37504 39376 37568
rect 39440 37504 39456 37568
rect 39520 37504 39528 37568
rect 39208 37503 39528 37504
rect 49208 37568 49528 37569
rect 49208 37504 49216 37568
rect 49280 37504 49296 37568
rect 49360 37504 49376 37568
rect 49440 37504 49456 37568
rect 49520 37504 49528 37568
rect 49208 37503 49528 37504
rect 59208 37568 59528 37569
rect 59208 37504 59216 37568
rect 59280 37504 59296 37568
rect 59360 37504 59376 37568
rect 59440 37504 59456 37568
rect 59520 37504 59528 37568
rect 69200 37544 70000 37574
rect 59208 37503 59528 37504
rect 4208 37024 4528 37025
rect 0 36954 800 36984
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 14208 37024 14528 37025
rect 14208 36960 14216 37024
rect 14280 36960 14296 37024
rect 14360 36960 14376 37024
rect 14440 36960 14456 37024
rect 14520 36960 14528 37024
rect 14208 36959 14528 36960
rect 24208 37024 24528 37025
rect 24208 36960 24216 37024
rect 24280 36960 24296 37024
rect 24360 36960 24376 37024
rect 24440 36960 24456 37024
rect 24520 36960 24528 37024
rect 24208 36959 24528 36960
rect 34208 37024 34528 37025
rect 34208 36960 34216 37024
rect 34280 36960 34296 37024
rect 34360 36960 34376 37024
rect 34440 36960 34456 37024
rect 34520 36960 34528 37024
rect 34208 36959 34528 36960
rect 44208 37024 44528 37025
rect 44208 36960 44216 37024
rect 44280 36960 44296 37024
rect 44360 36960 44376 37024
rect 44440 36960 44456 37024
rect 44520 36960 44528 37024
rect 44208 36959 44528 36960
rect 54208 37024 54528 37025
rect 54208 36960 54216 37024
rect 54280 36960 54296 37024
rect 54360 36960 54376 37024
rect 54440 36960 54456 37024
rect 54520 36960 54528 37024
rect 54208 36959 54528 36960
rect 64208 37024 64528 37025
rect 64208 36960 64216 37024
rect 64280 36960 64296 37024
rect 64360 36960 64376 37024
rect 64440 36960 64456 37024
rect 64520 36960 64528 37024
rect 64208 36959 64528 36960
rect 1577 36954 1643 36957
rect 0 36952 1643 36954
rect 0 36896 1582 36952
rect 1638 36896 1643 36952
rect 0 36894 1643 36896
rect 0 36864 800 36894
rect 1577 36891 1643 36894
rect 9208 36480 9528 36481
rect 9208 36416 9216 36480
rect 9280 36416 9296 36480
rect 9360 36416 9376 36480
rect 9440 36416 9456 36480
rect 9520 36416 9528 36480
rect 9208 36415 9528 36416
rect 19208 36480 19528 36481
rect 19208 36416 19216 36480
rect 19280 36416 19296 36480
rect 19360 36416 19376 36480
rect 19440 36416 19456 36480
rect 19520 36416 19528 36480
rect 19208 36415 19528 36416
rect 29208 36480 29528 36481
rect 29208 36416 29216 36480
rect 29280 36416 29296 36480
rect 29360 36416 29376 36480
rect 29440 36416 29456 36480
rect 29520 36416 29528 36480
rect 29208 36415 29528 36416
rect 39208 36480 39528 36481
rect 39208 36416 39216 36480
rect 39280 36416 39296 36480
rect 39360 36416 39376 36480
rect 39440 36416 39456 36480
rect 39520 36416 39528 36480
rect 39208 36415 39528 36416
rect 49208 36480 49528 36481
rect 49208 36416 49216 36480
rect 49280 36416 49296 36480
rect 49360 36416 49376 36480
rect 49440 36416 49456 36480
rect 49520 36416 49528 36480
rect 49208 36415 49528 36416
rect 59208 36480 59528 36481
rect 59208 36416 59216 36480
rect 59280 36416 59296 36480
rect 59360 36416 59376 36480
rect 59440 36416 59456 36480
rect 59520 36416 59528 36480
rect 59208 36415 59528 36416
rect 68093 36274 68159 36277
rect 69200 36274 70000 36304
rect 68093 36272 70000 36274
rect 68093 36216 68098 36272
rect 68154 36216 70000 36272
rect 68093 36214 70000 36216
rect 68093 36211 68159 36214
rect 69200 36184 70000 36214
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 14208 35936 14528 35937
rect 14208 35872 14216 35936
rect 14280 35872 14296 35936
rect 14360 35872 14376 35936
rect 14440 35872 14456 35936
rect 14520 35872 14528 35936
rect 14208 35871 14528 35872
rect 24208 35936 24528 35937
rect 24208 35872 24216 35936
rect 24280 35872 24296 35936
rect 24360 35872 24376 35936
rect 24440 35872 24456 35936
rect 24520 35872 24528 35936
rect 24208 35871 24528 35872
rect 34208 35936 34528 35937
rect 34208 35872 34216 35936
rect 34280 35872 34296 35936
rect 34360 35872 34376 35936
rect 34440 35872 34456 35936
rect 34520 35872 34528 35936
rect 34208 35871 34528 35872
rect 44208 35936 44528 35937
rect 44208 35872 44216 35936
rect 44280 35872 44296 35936
rect 44360 35872 44376 35936
rect 44440 35872 44456 35936
rect 44520 35872 44528 35936
rect 44208 35871 44528 35872
rect 54208 35936 54528 35937
rect 54208 35872 54216 35936
rect 54280 35872 54296 35936
rect 54360 35872 54376 35936
rect 54440 35872 54456 35936
rect 54520 35872 54528 35936
rect 54208 35871 54528 35872
rect 64208 35936 64528 35937
rect 64208 35872 64216 35936
rect 64280 35872 64296 35936
rect 64360 35872 64376 35936
rect 64440 35872 64456 35936
rect 64520 35872 64528 35936
rect 64208 35871 64528 35872
rect 0 35594 800 35624
rect 1761 35594 1827 35597
rect 0 35592 1827 35594
rect 0 35536 1766 35592
rect 1822 35536 1827 35592
rect 0 35534 1827 35536
rect 0 35504 800 35534
rect 1761 35531 1827 35534
rect 9208 35392 9528 35393
rect 9208 35328 9216 35392
rect 9280 35328 9296 35392
rect 9360 35328 9376 35392
rect 9440 35328 9456 35392
rect 9520 35328 9528 35392
rect 9208 35327 9528 35328
rect 19208 35392 19528 35393
rect 19208 35328 19216 35392
rect 19280 35328 19296 35392
rect 19360 35328 19376 35392
rect 19440 35328 19456 35392
rect 19520 35328 19528 35392
rect 19208 35327 19528 35328
rect 29208 35392 29528 35393
rect 29208 35328 29216 35392
rect 29280 35328 29296 35392
rect 29360 35328 29376 35392
rect 29440 35328 29456 35392
rect 29520 35328 29528 35392
rect 29208 35327 29528 35328
rect 39208 35392 39528 35393
rect 39208 35328 39216 35392
rect 39280 35328 39296 35392
rect 39360 35328 39376 35392
rect 39440 35328 39456 35392
rect 39520 35328 39528 35392
rect 39208 35327 39528 35328
rect 49208 35392 49528 35393
rect 49208 35328 49216 35392
rect 49280 35328 49296 35392
rect 49360 35328 49376 35392
rect 49440 35328 49456 35392
rect 49520 35328 49528 35392
rect 49208 35327 49528 35328
rect 59208 35392 59528 35393
rect 59208 35328 59216 35392
rect 59280 35328 59296 35392
rect 59360 35328 59376 35392
rect 59440 35328 59456 35392
rect 59520 35328 59528 35392
rect 59208 35327 59528 35328
rect 68921 34914 68987 34917
rect 69200 34914 70000 34944
rect 68921 34912 70000 34914
rect 68921 34856 68926 34912
rect 68982 34856 70000 34912
rect 68921 34854 70000 34856
rect 68921 34851 68987 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 14208 34848 14528 34849
rect 14208 34784 14216 34848
rect 14280 34784 14296 34848
rect 14360 34784 14376 34848
rect 14440 34784 14456 34848
rect 14520 34784 14528 34848
rect 14208 34783 14528 34784
rect 24208 34848 24528 34849
rect 24208 34784 24216 34848
rect 24280 34784 24296 34848
rect 24360 34784 24376 34848
rect 24440 34784 24456 34848
rect 24520 34784 24528 34848
rect 24208 34783 24528 34784
rect 34208 34848 34528 34849
rect 34208 34784 34216 34848
rect 34280 34784 34296 34848
rect 34360 34784 34376 34848
rect 34440 34784 34456 34848
rect 34520 34784 34528 34848
rect 34208 34783 34528 34784
rect 44208 34848 44528 34849
rect 44208 34784 44216 34848
rect 44280 34784 44296 34848
rect 44360 34784 44376 34848
rect 44440 34784 44456 34848
rect 44520 34784 44528 34848
rect 44208 34783 44528 34784
rect 54208 34848 54528 34849
rect 54208 34784 54216 34848
rect 54280 34784 54296 34848
rect 54360 34784 54376 34848
rect 54440 34784 54456 34848
rect 54520 34784 54528 34848
rect 54208 34783 54528 34784
rect 64208 34848 64528 34849
rect 64208 34784 64216 34848
rect 64280 34784 64296 34848
rect 64360 34784 64376 34848
rect 64440 34784 64456 34848
rect 64520 34784 64528 34848
rect 69200 34824 70000 34854
rect 64208 34783 64528 34784
rect 32765 34642 32831 34645
rect 33869 34642 33935 34645
rect 32765 34640 33935 34642
rect 32765 34584 32770 34640
rect 32826 34584 33874 34640
rect 33930 34584 33935 34640
rect 32765 34582 33935 34584
rect 32765 34579 32831 34582
rect 33869 34579 33935 34582
rect 9208 34304 9528 34305
rect 0 34234 800 34264
rect 9208 34240 9216 34304
rect 9280 34240 9296 34304
rect 9360 34240 9376 34304
rect 9440 34240 9456 34304
rect 9520 34240 9528 34304
rect 9208 34239 9528 34240
rect 19208 34304 19528 34305
rect 19208 34240 19216 34304
rect 19280 34240 19296 34304
rect 19360 34240 19376 34304
rect 19440 34240 19456 34304
rect 19520 34240 19528 34304
rect 19208 34239 19528 34240
rect 29208 34304 29528 34305
rect 29208 34240 29216 34304
rect 29280 34240 29296 34304
rect 29360 34240 29376 34304
rect 29440 34240 29456 34304
rect 29520 34240 29528 34304
rect 29208 34239 29528 34240
rect 39208 34304 39528 34305
rect 39208 34240 39216 34304
rect 39280 34240 39296 34304
rect 39360 34240 39376 34304
rect 39440 34240 39456 34304
rect 39520 34240 39528 34304
rect 39208 34239 39528 34240
rect 49208 34304 49528 34305
rect 49208 34240 49216 34304
rect 49280 34240 49296 34304
rect 49360 34240 49376 34304
rect 49440 34240 49456 34304
rect 49520 34240 49528 34304
rect 49208 34239 49528 34240
rect 59208 34304 59528 34305
rect 59208 34240 59216 34304
rect 59280 34240 59296 34304
rect 59360 34240 59376 34304
rect 59440 34240 59456 34304
rect 59520 34240 59528 34304
rect 59208 34239 59528 34240
rect 1853 34234 1919 34237
rect 0 34232 1919 34234
rect 0 34176 1858 34232
rect 1914 34176 1919 34232
rect 0 34174 1919 34176
rect 0 34144 800 34174
rect 1853 34171 1919 34174
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 14208 33760 14528 33761
rect 14208 33696 14216 33760
rect 14280 33696 14296 33760
rect 14360 33696 14376 33760
rect 14440 33696 14456 33760
rect 14520 33696 14528 33760
rect 14208 33695 14528 33696
rect 24208 33760 24528 33761
rect 24208 33696 24216 33760
rect 24280 33696 24296 33760
rect 24360 33696 24376 33760
rect 24440 33696 24456 33760
rect 24520 33696 24528 33760
rect 24208 33695 24528 33696
rect 34208 33760 34528 33761
rect 34208 33696 34216 33760
rect 34280 33696 34296 33760
rect 34360 33696 34376 33760
rect 34440 33696 34456 33760
rect 34520 33696 34528 33760
rect 34208 33695 34528 33696
rect 44208 33760 44528 33761
rect 44208 33696 44216 33760
rect 44280 33696 44296 33760
rect 44360 33696 44376 33760
rect 44440 33696 44456 33760
rect 44520 33696 44528 33760
rect 44208 33695 44528 33696
rect 54208 33760 54528 33761
rect 54208 33696 54216 33760
rect 54280 33696 54296 33760
rect 54360 33696 54376 33760
rect 54440 33696 54456 33760
rect 54520 33696 54528 33760
rect 54208 33695 54528 33696
rect 64208 33760 64528 33761
rect 64208 33696 64216 33760
rect 64280 33696 64296 33760
rect 64360 33696 64376 33760
rect 64440 33696 64456 33760
rect 64520 33696 64528 33760
rect 64208 33695 64528 33696
rect 65149 33554 65215 33557
rect 69200 33554 70000 33584
rect 65149 33552 70000 33554
rect 65149 33496 65154 33552
rect 65210 33496 70000 33552
rect 65149 33494 70000 33496
rect 65149 33491 65215 33494
rect 69200 33464 70000 33494
rect 9208 33216 9528 33217
rect 9208 33152 9216 33216
rect 9280 33152 9296 33216
rect 9360 33152 9376 33216
rect 9440 33152 9456 33216
rect 9520 33152 9528 33216
rect 9208 33151 9528 33152
rect 19208 33216 19528 33217
rect 19208 33152 19216 33216
rect 19280 33152 19296 33216
rect 19360 33152 19376 33216
rect 19440 33152 19456 33216
rect 19520 33152 19528 33216
rect 19208 33151 19528 33152
rect 29208 33216 29528 33217
rect 29208 33152 29216 33216
rect 29280 33152 29296 33216
rect 29360 33152 29376 33216
rect 29440 33152 29456 33216
rect 29520 33152 29528 33216
rect 29208 33151 29528 33152
rect 39208 33216 39528 33217
rect 39208 33152 39216 33216
rect 39280 33152 39296 33216
rect 39360 33152 39376 33216
rect 39440 33152 39456 33216
rect 39520 33152 39528 33216
rect 39208 33151 39528 33152
rect 49208 33216 49528 33217
rect 49208 33152 49216 33216
rect 49280 33152 49296 33216
rect 49360 33152 49376 33216
rect 49440 33152 49456 33216
rect 49520 33152 49528 33216
rect 49208 33151 49528 33152
rect 59208 33216 59528 33217
rect 59208 33152 59216 33216
rect 59280 33152 59296 33216
rect 59360 33152 59376 33216
rect 59440 33152 59456 33216
rect 59520 33152 59528 33216
rect 59208 33151 59528 33152
rect 0 32920 800 33040
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 14208 32672 14528 32673
rect 14208 32608 14216 32672
rect 14280 32608 14296 32672
rect 14360 32608 14376 32672
rect 14440 32608 14456 32672
rect 14520 32608 14528 32672
rect 14208 32607 14528 32608
rect 24208 32672 24528 32673
rect 24208 32608 24216 32672
rect 24280 32608 24296 32672
rect 24360 32608 24376 32672
rect 24440 32608 24456 32672
rect 24520 32608 24528 32672
rect 24208 32607 24528 32608
rect 34208 32672 34528 32673
rect 34208 32608 34216 32672
rect 34280 32608 34296 32672
rect 34360 32608 34376 32672
rect 34440 32608 34456 32672
rect 34520 32608 34528 32672
rect 34208 32607 34528 32608
rect 44208 32672 44528 32673
rect 44208 32608 44216 32672
rect 44280 32608 44296 32672
rect 44360 32608 44376 32672
rect 44440 32608 44456 32672
rect 44520 32608 44528 32672
rect 44208 32607 44528 32608
rect 54208 32672 54528 32673
rect 54208 32608 54216 32672
rect 54280 32608 54296 32672
rect 54360 32608 54376 32672
rect 54440 32608 54456 32672
rect 54520 32608 54528 32672
rect 54208 32607 54528 32608
rect 64208 32672 64528 32673
rect 64208 32608 64216 32672
rect 64280 32608 64296 32672
rect 64360 32608 64376 32672
rect 64440 32608 64456 32672
rect 64520 32608 64528 32672
rect 64208 32607 64528 32608
rect 7189 32466 7255 32469
rect 38694 32466 38700 32468
rect 7189 32464 38700 32466
rect 7189 32408 7194 32464
rect 7250 32408 38700 32464
rect 7189 32406 38700 32408
rect 7189 32403 7255 32406
rect 38694 32404 38700 32406
rect 38764 32404 38770 32468
rect 68093 32330 68159 32333
rect 69200 32330 70000 32360
rect 68093 32328 70000 32330
rect 68093 32272 68098 32328
rect 68154 32272 70000 32328
rect 68093 32270 70000 32272
rect 68093 32267 68159 32270
rect 69200 32240 70000 32270
rect 9208 32128 9528 32129
rect 9208 32064 9216 32128
rect 9280 32064 9296 32128
rect 9360 32064 9376 32128
rect 9440 32064 9456 32128
rect 9520 32064 9528 32128
rect 9208 32063 9528 32064
rect 19208 32128 19528 32129
rect 19208 32064 19216 32128
rect 19280 32064 19296 32128
rect 19360 32064 19376 32128
rect 19440 32064 19456 32128
rect 19520 32064 19528 32128
rect 19208 32063 19528 32064
rect 29208 32128 29528 32129
rect 29208 32064 29216 32128
rect 29280 32064 29296 32128
rect 29360 32064 29376 32128
rect 29440 32064 29456 32128
rect 29520 32064 29528 32128
rect 29208 32063 29528 32064
rect 39208 32128 39528 32129
rect 39208 32064 39216 32128
rect 39280 32064 39296 32128
rect 39360 32064 39376 32128
rect 39440 32064 39456 32128
rect 39520 32064 39528 32128
rect 39208 32063 39528 32064
rect 49208 32128 49528 32129
rect 49208 32064 49216 32128
rect 49280 32064 49296 32128
rect 49360 32064 49376 32128
rect 49440 32064 49456 32128
rect 49520 32064 49528 32128
rect 49208 32063 49528 32064
rect 59208 32128 59528 32129
rect 59208 32064 59216 32128
rect 59280 32064 59296 32128
rect 59360 32064 59376 32128
rect 59440 32064 59456 32128
rect 59520 32064 59528 32128
rect 59208 32063 59528 32064
rect 0 31650 800 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 800 31590
rect 1577 31587 1643 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 14208 31584 14528 31585
rect 14208 31520 14216 31584
rect 14280 31520 14296 31584
rect 14360 31520 14376 31584
rect 14440 31520 14456 31584
rect 14520 31520 14528 31584
rect 14208 31519 14528 31520
rect 24208 31584 24528 31585
rect 24208 31520 24216 31584
rect 24280 31520 24296 31584
rect 24360 31520 24376 31584
rect 24440 31520 24456 31584
rect 24520 31520 24528 31584
rect 24208 31519 24528 31520
rect 34208 31584 34528 31585
rect 34208 31520 34216 31584
rect 34280 31520 34296 31584
rect 34360 31520 34376 31584
rect 34440 31520 34456 31584
rect 34520 31520 34528 31584
rect 34208 31519 34528 31520
rect 44208 31584 44528 31585
rect 44208 31520 44216 31584
rect 44280 31520 44296 31584
rect 44360 31520 44376 31584
rect 44440 31520 44456 31584
rect 44520 31520 44528 31584
rect 44208 31519 44528 31520
rect 54208 31584 54528 31585
rect 54208 31520 54216 31584
rect 54280 31520 54296 31584
rect 54360 31520 54376 31584
rect 54440 31520 54456 31584
rect 54520 31520 54528 31584
rect 54208 31519 54528 31520
rect 64208 31584 64528 31585
rect 64208 31520 64216 31584
rect 64280 31520 64296 31584
rect 64360 31520 64376 31584
rect 64440 31520 64456 31584
rect 64520 31520 64528 31584
rect 64208 31519 64528 31520
rect 9208 31040 9528 31041
rect 9208 30976 9216 31040
rect 9280 30976 9296 31040
rect 9360 30976 9376 31040
rect 9440 30976 9456 31040
rect 9520 30976 9528 31040
rect 9208 30975 9528 30976
rect 19208 31040 19528 31041
rect 19208 30976 19216 31040
rect 19280 30976 19296 31040
rect 19360 30976 19376 31040
rect 19440 30976 19456 31040
rect 19520 30976 19528 31040
rect 19208 30975 19528 30976
rect 29208 31040 29528 31041
rect 29208 30976 29216 31040
rect 29280 30976 29296 31040
rect 29360 30976 29376 31040
rect 29440 30976 29456 31040
rect 29520 30976 29528 31040
rect 29208 30975 29528 30976
rect 39208 31040 39528 31041
rect 39208 30976 39216 31040
rect 39280 30976 39296 31040
rect 39360 30976 39376 31040
rect 39440 30976 39456 31040
rect 39520 30976 39528 31040
rect 39208 30975 39528 30976
rect 49208 31040 49528 31041
rect 49208 30976 49216 31040
rect 49280 30976 49296 31040
rect 49360 30976 49376 31040
rect 49440 30976 49456 31040
rect 49520 30976 49528 31040
rect 49208 30975 49528 30976
rect 59208 31040 59528 31041
rect 59208 30976 59216 31040
rect 59280 30976 59296 31040
rect 59360 30976 59376 31040
rect 59440 30976 59456 31040
rect 59520 30976 59528 31040
rect 59208 30975 59528 30976
rect 68093 30970 68159 30973
rect 69200 30970 70000 31000
rect 68093 30968 70000 30970
rect 68093 30912 68098 30968
rect 68154 30912 70000 30968
rect 68093 30910 70000 30912
rect 68093 30907 68159 30910
rect 69200 30880 70000 30910
rect 4208 30496 4528 30497
rect 0 30426 800 30456
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 14208 30496 14528 30497
rect 14208 30432 14216 30496
rect 14280 30432 14296 30496
rect 14360 30432 14376 30496
rect 14440 30432 14456 30496
rect 14520 30432 14528 30496
rect 14208 30431 14528 30432
rect 24208 30496 24528 30497
rect 24208 30432 24216 30496
rect 24280 30432 24296 30496
rect 24360 30432 24376 30496
rect 24440 30432 24456 30496
rect 24520 30432 24528 30496
rect 24208 30431 24528 30432
rect 34208 30496 34528 30497
rect 34208 30432 34216 30496
rect 34280 30432 34296 30496
rect 34360 30432 34376 30496
rect 34440 30432 34456 30496
rect 34520 30432 34528 30496
rect 34208 30431 34528 30432
rect 44208 30496 44528 30497
rect 44208 30432 44216 30496
rect 44280 30432 44296 30496
rect 44360 30432 44376 30496
rect 44440 30432 44456 30496
rect 44520 30432 44528 30496
rect 44208 30431 44528 30432
rect 54208 30496 54528 30497
rect 54208 30432 54216 30496
rect 54280 30432 54296 30496
rect 54360 30432 54376 30496
rect 54440 30432 54456 30496
rect 54520 30432 54528 30496
rect 54208 30431 54528 30432
rect 64208 30496 64528 30497
rect 64208 30432 64216 30496
rect 64280 30432 64296 30496
rect 64360 30432 64376 30496
rect 64440 30432 64456 30496
rect 64520 30432 64528 30496
rect 64208 30431 64528 30432
rect 1761 30426 1827 30429
rect 0 30424 1827 30426
rect 0 30368 1766 30424
rect 1822 30368 1827 30424
rect 0 30366 1827 30368
rect 0 30336 800 30366
rect 1761 30363 1827 30366
rect 9208 29952 9528 29953
rect 9208 29888 9216 29952
rect 9280 29888 9296 29952
rect 9360 29888 9376 29952
rect 9440 29888 9456 29952
rect 9520 29888 9528 29952
rect 9208 29887 9528 29888
rect 19208 29952 19528 29953
rect 19208 29888 19216 29952
rect 19280 29888 19296 29952
rect 19360 29888 19376 29952
rect 19440 29888 19456 29952
rect 19520 29888 19528 29952
rect 19208 29887 19528 29888
rect 29208 29952 29528 29953
rect 29208 29888 29216 29952
rect 29280 29888 29296 29952
rect 29360 29888 29376 29952
rect 29440 29888 29456 29952
rect 29520 29888 29528 29952
rect 29208 29887 29528 29888
rect 39208 29952 39528 29953
rect 39208 29888 39216 29952
rect 39280 29888 39296 29952
rect 39360 29888 39376 29952
rect 39440 29888 39456 29952
rect 39520 29888 39528 29952
rect 39208 29887 39528 29888
rect 49208 29952 49528 29953
rect 49208 29888 49216 29952
rect 49280 29888 49296 29952
rect 49360 29888 49376 29952
rect 49440 29888 49456 29952
rect 49520 29888 49528 29952
rect 49208 29887 49528 29888
rect 59208 29952 59528 29953
rect 59208 29888 59216 29952
rect 59280 29888 59296 29952
rect 59360 29888 59376 29952
rect 59440 29888 59456 29952
rect 59520 29888 59528 29952
rect 59208 29887 59528 29888
rect 68093 29610 68159 29613
rect 69200 29610 70000 29640
rect 68093 29608 70000 29610
rect 68093 29552 68098 29608
rect 68154 29552 70000 29608
rect 68093 29550 70000 29552
rect 68093 29547 68159 29550
rect 69200 29520 70000 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 14208 29408 14528 29409
rect 14208 29344 14216 29408
rect 14280 29344 14296 29408
rect 14360 29344 14376 29408
rect 14440 29344 14456 29408
rect 14520 29344 14528 29408
rect 14208 29343 14528 29344
rect 24208 29408 24528 29409
rect 24208 29344 24216 29408
rect 24280 29344 24296 29408
rect 24360 29344 24376 29408
rect 24440 29344 24456 29408
rect 24520 29344 24528 29408
rect 24208 29343 24528 29344
rect 34208 29408 34528 29409
rect 34208 29344 34216 29408
rect 34280 29344 34296 29408
rect 34360 29344 34376 29408
rect 34440 29344 34456 29408
rect 34520 29344 34528 29408
rect 34208 29343 34528 29344
rect 44208 29408 44528 29409
rect 44208 29344 44216 29408
rect 44280 29344 44296 29408
rect 44360 29344 44376 29408
rect 44440 29344 44456 29408
rect 44520 29344 44528 29408
rect 44208 29343 44528 29344
rect 54208 29408 54528 29409
rect 54208 29344 54216 29408
rect 54280 29344 54296 29408
rect 54360 29344 54376 29408
rect 54440 29344 54456 29408
rect 54520 29344 54528 29408
rect 54208 29343 54528 29344
rect 64208 29408 64528 29409
rect 64208 29344 64216 29408
rect 64280 29344 64296 29408
rect 64360 29344 64376 29408
rect 64440 29344 64456 29408
rect 64520 29344 64528 29408
rect 64208 29343 64528 29344
rect 0 29066 800 29096
rect 1761 29066 1827 29069
rect 0 29064 1827 29066
rect 0 29008 1766 29064
rect 1822 29008 1827 29064
rect 0 29006 1827 29008
rect 0 28976 800 29006
rect 1761 29003 1827 29006
rect 9208 28864 9528 28865
rect 9208 28800 9216 28864
rect 9280 28800 9296 28864
rect 9360 28800 9376 28864
rect 9440 28800 9456 28864
rect 9520 28800 9528 28864
rect 9208 28799 9528 28800
rect 19208 28864 19528 28865
rect 19208 28800 19216 28864
rect 19280 28800 19296 28864
rect 19360 28800 19376 28864
rect 19440 28800 19456 28864
rect 19520 28800 19528 28864
rect 19208 28799 19528 28800
rect 29208 28864 29528 28865
rect 29208 28800 29216 28864
rect 29280 28800 29296 28864
rect 29360 28800 29376 28864
rect 29440 28800 29456 28864
rect 29520 28800 29528 28864
rect 29208 28799 29528 28800
rect 39208 28864 39528 28865
rect 39208 28800 39216 28864
rect 39280 28800 39296 28864
rect 39360 28800 39376 28864
rect 39440 28800 39456 28864
rect 39520 28800 39528 28864
rect 39208 28799 39528 28800
rect 49208 28864 49528 28865
rect 49208 28800 49216 28864
rect 49280 28800 49296 28864
rect 49360 28800 49376 28864
rect 49440 28800 49456 28864
rect 49520 28800 49528 28864
rect 49208 28799 49528 28800
rect 59208 28864 59528 28865
rect 59208 28800 59216 28864
rect 59280 28800 59296 28864
rect 59360 28800 59376 28864
rect 59440 28800 59456 28864
rect 59520 28800 59528 28864
rect 59208 28799 59528 28800
rect 66161 28386 66227 28389
rect 69200 28386 70000 28416
rect 66161 28384 70000 28386
rect 66161 28328 66166 28384
rect 66222 28328 70000 28384
rect 66161 28326 70000 28328
rect 66161 28323 66227 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 14208 28320 14528 28321
rect 14208 28256 14216 28320
rect 14280 28256 14296 28320
rect 14360 28256 14376 28320
rect 14440 28256 14456 28320
rect 14520 28256 14528 28320
rect 14208 28255 14528 28256
rect 24208 28320 24528 28321
rect 24208 28256 24216 28320
rect 24280 28256 24296 28320
rect 24360 28256 24376 28320
rect 24440 28256 24456 28320
rect 24520 28256 24528 28320
rect 24208 28255 24528 28256
rect 34208 28320 34528 28321
rect 34208 28256 34216 28320
rect 34280 28256 34296 28320
rect 34360 28256 34376 28320
rect 34440 28256 34456 28320
rect 34520 28256 34528 28320
rect 34208 28255 34528 28256
rect 44208 28320 44528 28321
rect 44208 28256 44216 28320
rect 44280 28256 44296 28320
rect 44360 28256 44376 28320
rect 44440 28256 44456 28320
rect 44520 28256 44528 28320
rect 44208 28255 44528 28256
rect 54208 28320 54528 28321
rect 54208 28256 54216 28320
rect 54280 28256 54296 28320
rect 54360 28256 54376 28320
rect 54440 28256 54456 28320
rect 54520 28256 54528 28320
rect 54208 28255 54528 28256
rect 64208 28320 64528 28321
rect 64208 28256 64216 28320
rect 64280 28256 64296 28320
rect 64360 28256 64376 28320
rect 64440 28256 64456 28320
rect 64520 28256 64528 28320
rect 69200 28296 70000 28326
rect 64208 28255 64528 28256
rect 0 27752 800 27872
rect 9208 27776 9528 27777
rect 9208 27712 9216 27776
rect 9280 27712 9296 27776
rect 9360 27712 9376 27776
rect 9440 27712 9456 27776
rect 9520 27712 9528 27776
rect 9208 27711 9528 27712
rect 19208 27776 19528 27777
rect 19208 27712 19216 27776
rect 19280 27712 19296 27776
rect 19360 27712 19376 27776
rect 19440 27712 19456 27776
rect 19520 27712 19528 27776
rect 19208 27711 19528 27712
rect 29208 27776 29528 27777
rect 29208 27712 29216 27776
rect 29280 27712 29296 27776
rect 29360 27712 29376 27776
rect 29440 27712 29456 27776
rect 29520 27712 29528 27776
rect 29208 27711 29528 27712
rect 39208 27776 39528 27777
rect 39208 27712 39216 27776
rect 39280 27712 39296 27776
rect 39360 27712 39376 27776
rect 39440 27712 39456 27776
rect 39520 27712 39528 27776
rect 39208 27711 39528 27712
rect 49208 27776 49528 27777
rect 49208 27712 49216 27776
rect 49280 27712 49296 27776
rect 49360 27712 49376 27776
rect 49440 27712 49456 27776
rect 49520 27712 49528 27776
rect 49208 27711 49528 27712
rect 59208 27776 59528 27777
rect 59208 27712 59216 27776
rect 59280 27712 59296 27776
rect 59360 27712 59376 27776
rect 59440 27712 59456 27776
rect 59520 27712 59528 27776
rect 59208 27711 59528 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 14208 27232 14528 27233
rect 14208 27168 14216 27232
rect 14280 27168 14296 27232
rect 14360 27168 14376 27232
rect 14440 27168 14456 27232
rect 14520 27168 14528 27232
rect 14208 27167 14528 27168
rect 24208 27232 24528 27233
rect 24208 27168 24216 27232
rect 24280 27168 24296 27232
rect 24360 27168 24376 27232
rect 24440 27168 24456 27232
rect 24520 27168 24528 27232
rect 24208 27167 24528 27168
rect 34208 27232 34528 27233
rect 34208 27168 34216 27232
rect 34280 27168 34296 27232
rect 34360 27168 34376 27232
rect 34440 27168 34456 27232
rect 34520 27168 34528 27232
rect 34208 27167 34528 27168
rect 44208 27232 44528 27233
rect 44208 27168 44216 27232
rect 44280 27168 44296 27232
rect 44360 27168 44376 27232
rect 44440 27168 44456 27232
rect 44520 27168 44528 27232
rect 44208 27167 44528 27168
rect 54208 27232 54528 27233
rect 54208 27168 54216 27232
rect 54280 27168 54296 27232
rect 54360 27168 54376 27232
rect 54440 27168 54456 27232
rect 54520 27168 54528 27232
rect 54208 27167 54528 27168
rect 64208 27232 64528 27233
rect 64208 27168 64216 27232
rect 64280 27168 64296 27232
rect 64360 27168 64376 27232
rect 64440 27168 64456 27232
rect 64520 27168 64528 27232
rect 64208 27167 64528 27168
rect 68093 27026 68159 27029
rect 69200 27026 70000 27056
rect 68093 27024 70000 27026
rect 68093 26968 68098 27024
rect 68154 26968 70000 27024
rect 68093 26966 70000 26968
rect 68093 26963 68159 26966
rect 69200 26936 70000 26966
rect 9208 26688 9528 26689
rect 9208 26624 9216 26688
rect 9280 26624 9296 26688
rect 9360 26624 9376 26688
rect 9440 26624 9456 26688
rect 9520 26624 9528 26688
rect 9208 26623 9528 26624
rect 19208 26688 19528 26689
rect 19208 26624 19216 26688
rect 19280 26624 19296 26688
rect 19360 26624 19376 26688
rect 19440 26624 19456 26688
rect 19520 26624 19528 26688
rect 19208 26623 19528 26624
rect 29208 26688 29528 26689
rect 29208 26624 29216 26688
rect 29280 26624 29296 26688
rect 29360 26624 29376 26688
rect 29440 26624 29456 26688
rect 29520 26624 29528 26688
rect 29208 26623 29528 26624
rect 39208 26688 39528 26689
rect 39208 26624 39216 26688
rect 39280 26624 39296 26688
rect 39360 26624 39376 26688
rect 39440 26624 39456 26688
rect 39520 26624 39528 26688
rect 39208 26623 39528 26624
rect 49208 26688 49528 26689
rect 49208 26624 49216 26688
rect 49280 26624 49296 26688
rect 49360 26624 49376 26688
rect 49440 26624 49456 26688
rect 49520 26624 49528 26688
rect 49208 26623 49528 26624
rect 59208 26688 59528 26689
rect 59208 26624 59216 26688
rect 59280 26624 59296 26688
rect 59360 26624 59376 26688
rect 59440 26624 59456 26688
rect 59520 26624 59528 26688
rect 59208 26623 59528 26624
rect 0 26482 800 26512
rect 1577 26482 1643 26485
rect 0 26480 1643 26482
rect 0 26424 1582 26480
rect 1638 26424 1643 26480
rect 0 26422 1643 26424
rect 0 26392 800 26422
rect 1577 26419 1643 26422
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 14208 26144 14528 26145
rect 14208 26080 14216 26144
rect 14280 26080 14296 26144
rect 14360 26080 14376 26144
rect 14440 26080 14456 26144
rect 14520 26080 14528 26144
rect 14208 26079 14528 26080
rect 24208 26144 24528 26145
rect 24208 26080 24216 26144
rect 24280 26080 24296 26144
rect 24360 26080 24376 26144
rect 24440 26080 24456 26144
rect 24520 26080 24528 26144
rect 24208 26079 24528 26080
rect 34208 26144 34528 26145
rect 34208 26080 34216 26144
rect 34280 26080 34296 26144
rect 34360 26080 34376 26144
rect 34440 26080 34456 26144
rect 34520 26080 34528 26144
rect 34208 26079 34528 26080
rect 44208 26144 44528 26145
rect 44208 26080 44216 26144
rect 44280 26080 44296 26144
rect 44360 26080 44376 26144
rect 44440 26080 44456 26144
rect 44520 26080 44528 26144
rect 44208 26079 44528 26080
rect 54208 26144 54528 26145
rect 54208 26080 54216 26144
rect 54280 26080 54296 26144
rect 54360 26080 54376 26144
rect 54440 26080 54456 26144
rect 54520 26080 54528 26144
rect 54208 26079 54528 26080
rect 64208 26144 64528 26145
rect 64208 26080 64216 26144
rect 64280 26080 64296 26144
rect 64360 26080 64376 26144
rect 64440 26080 64456 26144
rect 64520 26080 64528 26144
rect 64208 26079 64528 26080
rect 68093 25666 68159 25669
rect 69200 25666 70000 25696
rect 68093 25664 70000 25666
rect 68093 25608 68098 25664
rect 68154 25608 70000 25664
rect 68093 25606 70000 25608
rect 68093 25603 68159 25606
rect 9208 25600 9528 25601
rect 9208 25536 9216 25600
rect 9280 25536 9296 25600
rect 9360 25536 9376 25600
rect 9440 25536 9456 25600
rect 9520 25536 9528 25600
rect 9208 25535 9528 25536
rect 19208 25600 19528 25601
rect 19208 25536 19216 25600
rect 19280 25536 19296 25600
rect 19360 25536 19376 25600
rect 19440 25536 19456 25600
rect 19520 25536 19528 25600
rect 19208 25535 19528 25536
rect 29208 25600 29528 25601
rect 29208 25536 29216 25600
rect 29280 25536 29296 25600
rect 29360 25536 29376 25600
rect 29440 25536 29456 25600
rect 29520 25536 29528 25600
rect 29208 25535 29528 25536
rect 39208 25600 39528 25601
rect 39208 25536 39216 25600
rect 39280 25536 39296 25600
rect 39360 25536 39376 25600
rect 39440 25536 39456 25600
rect 39520 25536 39528 25600
rect 39208 25535 39528 25536
rect 49208 25600 49528 25601
rect 49208 25536 49216 25600
rect 49280 25536 49296 25600
rect 49360 25536 49376 25600
rect 49440 25536 49456 25600
rect 49520 25536 49528 25600
rect 49208 25535 49528 25536
rect 59208 25600 59528 25601
rect 59208 25536 59216 25600
rect 59280 25536 59296 25600
rect 59360 25536 59376 25600
rect 59440 25536 59456 25600
rect 59520 25536 59528 25600
rect 69200 25576 70000 25606
rect 59208 25535 59528 25536
rect 0 25258 800 25288
rect 1761 25258 1827 25261
rect 0 25256 1827 25258
rect 0 25200 1766 25256
rect 1822 25200 1827 25256
rect 0 25198 1827 25200
rect 0 25168 800 25198
rect 1761 25195 1827 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 14208 25056 14528 25057
rect 14208 24992 14216 25056
rect 14280 24992 14296 25056
rect 14360 24992 14376 25056
rect 14440 24992 14456 25056
rect 14520 24992 14528 25056
rect 14208 24991 14528 24992
rect 24208 25056 24528 25057
rect 24208 24992 24216 25056
rect 24280 24992 24296 25056
rect 24360 24992 24376 25056
rect 24440 24992 24456 25056
rect 24520 24992 24528 25056
rect 24208 24991 24528 24992
rect 34208 25056 34528 25057
rect 34208 24992 34216 25056
rect 34280 24992 34296 25056
rect 34360 24992 34376 25056
rect 34440 24992 34456 25056
rect 34520 24992 34528 25056
rect 34208 24991 34528 24992
rect 44208 25056 44528 25057
rect 44208 24992 44216 25056
rect 44280 24992 44296 25056
rect 44360 24992 44376 25056
rect 44440 24992 44456 25056
rect 44520 24992 44528 25056
rect 44208 24991 44528 24992
rect 54208 25056 54528 25057
rect 54208 24992 54216 25056
rect 54280 24992 54296 25056
rect 54360 24992 54376 25056
rect 54440 24992 54456 25056
rect 54520 24992 54528 25056
rect 54208 24991 54528 24992
rect 64208 25056 64528 25057
rect 64208 24992 64216 25056
rect 64280 24992 64296 25056
rect 64360 24992 64376 25056
rect 64440 24992 64456 25056
rect 64520 24992 64528 25056
rect 64208 24991 64528 24992
rect 9208 24512 9528 24513
rect 9208 24448 9216 24512
rect 9280 24448 9296 24512
rect 9360 24448 9376 24512
rect 9440 24448 9456 24512
rect 9520 24448 9528 24512
rect 9208 24447 9528 24448
rect 19208 24512 19528 24513
rect 19208 24448 19216 24512
rect 19280 24448 19296 24512
rect 19360 24448 19376 24512
rect 19440 24448 19456 24512
rect 19520 24448 19528 24512
rect 19208 24447 19528 24448
rect 29208 24512 29528 24513
rect 29208 24448 29216 24512
rect 29280 24448 29296 24512
rect 29360 24448 29376 24512
rect 29440 24448 29456 24512
rect 29520 24448 29528 24512
rect 29208 24447 29528 24448
rect 39208 24512 39528 24513
rect 39208 24448 39216 24512
rect 39280 24448 39296 24512
rect 39360 24448 39376 24512
rect 39440 24448 39456 24512
rect 39520 24448 39528 24512
rect 39208 24447 39528 24448
rect 49208 24512 49528 24513
rect 49208 24448 49216 24512
rect 49280 24448 49296 24512
rect 49360 24448 49376 24512
rect 49440 24448 49456 24512
rect 49520 24448 49528 24512
rect 49208 24447 49528 24448
rect 59208 24512 59528 24513
rect 59208 24448 59216 24512
rect 59280 24448 59296 24512
rect 59360 24448 59376 24512
rect 59440 24448 59456 24512
rect 59520 24448 59528 24512
rect 59208 24447 59528 24448
rect 68093 24306 68159 24309
rect 69200 24306 70000 24336
rect 68093 24304 70000 24306
rect 68093 24248 68098 24304
rect 68154 24248 70000 24304
rect 68093 24246 70000 24248
rect 68093 24243 68159 24246
rect 69200 24216 70000 24246
rect 4208 23968 4528 23969
rect 0 23898 800 23928
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 14208 23968 14528 23969
rect 14208 23904 14216 23968
rect 14280 23904 14296 23968
rect 14360 23904 14376 23968
rect 14440 23904 14456 23968
rect 14520 23904 14528 23968
rect 14208 23903 14528 23904
rect 24208 23968 24528 23969
rect 24208 23904 24216 23968
rect 24280 23904 24296 23968
rect 24360 23904 24376 23968
rect 24440 23904 24456 23968
rect 24520 23904 24528 23968
rect 24208 23903 24528 23904
rect 34208 23968 34528 23969
rect 34208 23904 34216 23968
rect 34280 23904 34296 23968
rect 34360 23904 34376 23968
rect 34440 23904 34456 23968
rect 34520 23904 34528 23968
rect 34208 23903 34528 23904
rect 44208 23968 44528 23969
rect 44208 23904 44216 23968
rect 44280 23904 44296 23968
rect 44360 23904 44376 23968
rect 44440 23904 44456 23968
rect 44520 23904 44528 23968
rect 44208 23903 44528 23904
rect 54208 23968 54528 23969
rect 54208 23904 54216 23968
rect 54280 23904 54296 23968
rect 54360 23904 54376 23968
rect 54440 23904 54456 23968
rect 54520 23904 54528 23968
rect 54208 23903 54528 23904
rect 64208 23968 64528 23969
rect 64208 23904 64216 23968
rect 64280 23904 64296 23968
rect 64360 23904 64376 23968
rect 64440 23904 64456 23968
rect 64520 23904 64528 23968
rect 64208 23903 64528 23904
rect 1853 23898 1919 23901
rect 0 23896 1919 23898
rect 0 23840 1858 23896
rect 1914 23840 1919 23896
rect 0 23838 1919 23840
rect 0 23808 800 23838
rect 1853 23835 1919 23838
rect 9208 23424 9528 23425
rect 9208 23360 9216 23424
rect 9280 23360 9296 23424
rect 9360 23360 9376 23424
rect 9440 23360 9456 23424
rect 9520 23360 9528 23424
rect 9208 23359 9528 23360
rect 19208 23424 19528 23425
rect 19208 23360 19216 23424
rect 19280 23360 19296 23424
rect 19360 23360 19376 23424
rect 19440 23360 19456 23424
rect 19520 23360 19528 23424
rect 19208 23359 19528 23360
rect 29208 23424 29528 23425
rect 29208 23360 29216 23424
rect 29280 23360 29296 23424
rect 29360 23360 29376 23424
rect 29440 23360 29456 23424
rect 29520 23360 29528 23424
rect 29208 23359 29528 23360
rect 39208 23424 39528 23425
rect 39208 23360 39216 23424
rect 39280 23360 39296 23424
rect 39360 23360 39376 23424
rect 39440 23360 39456 23424
rect 39520 23360 39528 23424
rect 39208 23359 39528 23360
rect 49208 23424 49528 23425
rect 49208 23360 49216 23424
rect 49280 23360 49296 23424
rect 49360 23360 49376 23424
rect 49440 23360 49456 23424
rect 49520 23360 49528 23424
rect 49208 23359 49528 23360
rect 59208 23424 59528 23425
rect 59208 23360 59216 23424
rect 59280 23360 59296 23424
rect 59360 23360 59376 23424
rect 59440 23360 59456 23424
rect 59520 23360 59528 23424
rect 59208 23359 59528 23360
rect 68093 23082 68159 23085
rect 69200 23082 70000 23112
rect 68093 23080 70000 23082
rect 68093 23024 68098 23080
rect 68154 23024 70000 23080
rect 68093 23022 70000 23024
rect 68093 23019 68159 23022
rect 69200 22992 70000 23022
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 14208 22880 14528 22881
rect 14208 22816 14216 22880
rect 14280 22816 14296 22880
rect 14360 22816 14376 22880
rect 14440 22816 14456 22880
rect 14520 22816 14528 22880
rect 14208 22815 14528 22816
rect 24208 22880 24528 22881
rect 24208 22816 24216 22880
rect 24280 22816 24296 22880
rect 24360 22816 24376 22880
rect 24440 22816 24456 22880
rect 24520 22816 24528 22880
rect 24208 22815 24528 22816
rect 34208 22880 34528 22881
rect 34208 22816 34216 22880
rect 34280 22816 34296 22880
rect 34360 22816 34376 22880
rect 34440 22816 34456 22880
rect 34520 22816 34528 22880
rect 34208 22815 34528 22816
rect 44208 22880 44528 22881
rect 44208 22816 44216 22880
rect 44280 22816 44296 22880
rect 44360 22816 44376 22880
rect 44440 22816 44456 22880
rect 44520 22816 44528 22880
rect 44208 22815 44528 22816
rect 54208 22880 54528 22881
rect 54208 22816 54216 22880
rect 54280 22816 54296 22880
rect 54360 22816 54376 22880
rect 54440 22816 54456 22880
rect 54520 22816 54528 22880
rect 54208 22815 54528 22816
rect 64208 22880 64528 22881
rect 64208 22816 64216 22880
rect 64280 22816 64296 22880
rect 64360 22816 64376 22880
rect 64440 22816 64456 22880
rect 64520 22816 64528 22880
rect 64208 22815 64528 22816
rect 0 22584 800 22704
rect 9208 22336 9528 22337
rect 9208 22272 9216 22336
rect 9280 22272 9296 22336
rect 9360 22272 9376 22336
rect 9440 22272 9456 22336
rect 9520 22272 9528 22336
rect 9208 22271 9528 22272
rect 19208 22336 19528 22337
rect 19208 22272 19216 22336
rect 19280 22272 19296 22336
rect 19360 22272 19376 22336
rect 19440 22272 19456 22336
rect 19520 22272 19528 22336
rect 19208 22271 19528 22272
rect 29208 22336 29528 22337
rect 29208 22272 29216 22336
rect 29280 22272 29296 22336
rect 29360 22272 29376 22336
rect 29440 22272 29456 22336
rect 29520 22272 29528 22336
rect 29208 22271 29528 22272
rect 39208 22336 39528 22337
rect 39208 22272 39216 22336
rect 39280 22272 39296 22336
rect 39360 22272 39376 22336
rect 39440 22272 39456 22336
rect 39520 22272 39528 22336
rect 39208 22271 39528 22272
rect 49208 22336 49528 22337
rect 49208 22272 49216 22336
rect 49280 22272 49296 22336
rect 49360 22272 49376 22336
rect 49440 22272 49456 22336
rect 49520 22272 49528 22336
rect 49208 22271 49528 22272
rect 59208 22336 59528 22337
rect 59208 22272 59216 22336
rect 59280 22272 59296 22336
rect 59360 22272 59376 22336
rect 59440 22272 59456 22336
rect 59520 22272 59528 22336
rect 59208 22271 59528 22272
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 14208 21792 14528 21793
rect 14208 21728 14216 21792
rect 14280 21728 14296 21792
rect 14360 21728 14376 21792
rect 14440 21728 14456 21792
rect 14520 21728 14528 21792
rect 14208 21727 14528 21728
rect 24208 21792 24528 21793
rect 24208 21728 24216 21792
rect 24280 21728 24296 21792
rect 24360 21728 24376 21792
rect 24440 21728 24456 21792
rect 24520 21728 24528 21792
rect 24208 21727 24528 21728
rect 34208 21792 34528 21793
rect 34208 21728 34216 21792
rect 34280 21728 34296 21792
rect 34360 21728 34376 21792
rect 34440 21728 34456 21792
rect 34520 21728 34528 21792
rect 34208 21727 34528 21728
rect 44208 21792 44528 21793
rect 44208 21728 44216 21792
rect 44280 21728 44296 21792
rect 44360 21728 44376 21792
rect 44440 21728 44456 21792
rect 44520 21728 44528 21792
rect 44208 21727 44528 21728
rect 54208 21792 54528 21793
rect 54208 21728 54216 21792
rect 54280 21728 54296 21792
rect 54360 21728 54376 21792
rect 54440 21728 54456 21792
rect 54520 21728 54528 21792
rect 54208 21727 54528 21728
rect 64208 21792 64528 21793
rect 64208 21728 64216 21792
rect 64280 21728 64296 21792
rect 64360 21728 64376 21792
rect 64440 21728 64456 21792
rect 64520 21728 64528 21792
rect 64208 21727 64528 21728
rect 68093 21722 68159 21725
rect 69200 21722 70000 21752
rect 68093 21720 70000 21722
rect 68093 21664 68098 21720
rect 68154 21664 70000 21720
rect 68093 21662 70000 21664
rect 68093 21659 68159 21662
rect 69200 21632 70000 21662
rect 7373 21450 7439 21453
rect 39062 21450 39068 21452
rect 7373 21448 39068 21450
rect 7373 21392 7378 21448
rect 7434 21392 39068 21448
rect 7373 21390 39068 21392
rect 7373 21387 7439 21390
rect 39062 21388 39068 21390
rect 39132 21388 39138 21452
rect 0 21314 800 21344
rect 1393 21314 1459 21317
rect 0 21312 1459 21314
rect 0 21256 1398 21312
rect 1454 21256 1459 21312
rect 0 21254 1459 21256
rect 0 21224 800 21254
rect 1393 21251 1459 21254
rect 9208 21248 9528 21249
rect 9208 21184 9216 21248
rect 9280 21184 9296 21248
rect 9360 21184 9376 21248
rect 9440 21184 9456 21248
rect 9520 21184 9528 21248
rect 9208 21183 9528 21184
rect 19208 21248 19528 21249
rect 19208 21184 19216 21248
rect 19280 21184 19296 21248
rect 19360 21184 19376 21248
rect 19440 21184 19456 21248
rect 19520 21184 19528 21248
rect 19208 21183 19528 21184
rect 29208 21248 29528 21249
rect 29208 21184 29216 21248
rect 29280 21184 29296 21248
rect 29360 21184 29376 21248
rect 29440 21184 29456 21248
rect 29520 21184 29528 21248
rect 29208 21183 29528 21184
rect 39208 21248 39528 21249
rect 39208 21184 39216 21248
rect 39280 21184 39296 21248
rect 39360 21184 39376 21248
rect 39440 21184 39456 21248
rect 39520 21184 39528 21248
rect 39208 21183 39528 21184
rect 49208 21248 49528 21249
rect 49208 21184 49216 21248
rect 49280 21184 49296 21248
rect 49360 21184 49376 21248
rect 49440 21184 49456 21248
rect 49520 21184 49528 21248
rect 49208 21183 49528 21184
rect 59208 21248 59528 21249
rect 59208 21184 59216 21248
rect 59280 21184 59296 21248
rect 59360 21184 59376 21248
rect 59440 21184 59456 21248
rect 59520 21184 59528 21248
rect 59208 21183 59528 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 14208 20704 14528 20705
rect 14208 20640 14216 20704
rect 14280 20640 14296 20704
rect 14360 20640 14376 20704
rect 14440 20640 14456 20704
rect 14520 20640 14528 20704
rect 14208 20639 14528 20640
rect 24208 20704 24528 20705
rect 24208 20640 24216 20704
rect 24280 20640 24296 20704
rect 24360 20640 24376 20704
rect 24440 20640 24456 20704
rect 24520 20640 24528 20704
rect 24208 20639 24528 20640
rect 34208 20704 34528 20705
rect 34208 20640 34216 20704
rect 34280 20640 34296 20704
rect 34360 20640 34376 20704
rect 34440 20640 34456 20704
rect 34520 20640 34528 20704
rect 34208 20639 34528 20640
rect 44208 20704 44528 20705
rect 44208 20640 44216 20704
rect 44280 20640 44296 20704
rect 44360 20640 44376 20704
rect 44440 20640 44456 20704
rect 44520 20640 44528 20704
rect 44208 20639 44528 20640
rect 54208 20704 54528 20705
rect 54208 20640 54216 20704
rect 54280 20640 54296 20704
rect 54360 20640 54376 20704
rect 54440 20640 54456 20704
rect 54520 20640 54528 20704
rect 54208 20639 54528 20640
rect 64208 20704 64528 20705
rect 64208 20640 64216 20704
rect 64280 20640 64296 20704
rect 64360 20640 64376 20704
rect 64440 20640 64456 20704
rect 64520 20640 64528 20704
rect 64208 20639 64528 20640
rect 68093 20362 68159 20365
rect 69200 20362 70000 20392
rect 68093 20360 70000 20362
rect 68093 20304 68098 20360
rect 68154 20304 70000 20360
rect 68093 20302 70000 20304
rect 68093 20299 68159 20302
rect 69200 20272 70000 20302
rect 9208 20160 9528 20161
rect 0 20090 800 20120
rect 9208 20096 9216 20160
rect 9280 20096 9296 20160
rect 9360 20096 9376 20160
rect 9440 20096 9456 20160
rect 9520 20096 9528 20160
rect 9208 20095 9528 20096
rect 19208 20160 19528 20161
rect 19208 20096 19216 20160
rect 19280 20096 19296 20160
rect 19360 20096 19376 20160
rect 19440 20096 19456 20160
rect 19520 20096 19528 20160
rect 19208 20095 19528 20096
rect 29208 20160 29528 20161
rect 29208 20096 29216 20160
rect 29280 20096 29296 20160
rect 29360 20096 29376 20160
rect 29440 20096 29456 20160
rect 29520 20096 29528 20160
rect 29208 20095 29528 20096
rect 39208 20160 39528 20161
rect 39208 20096 39216 20160
rect 39280 20096 39296 20160
rect 39360 20096 39376 20160
rect 39440 20096 39456 20160
rect 39520 20096 39528 20160
rect 39208 20095 39528 20096
rect 49208 20160 49528 20161
rect 49208 20096 49216 20160
rect 49280 20096 49296 20160
rect 49360 20096 49376 20160
rect 49440 20096 49456 20160
rect 49520 20096 49528 20160
rect 49208 20095 49528 20096
rect 59208 20160 59528 20161
rect 59208 20096 59216 20160
rect 59280 20096 59296 20160
rect 59360 20096 59376 20160
rect 59440 20096 59456 20160
rect 59520 20096 59528 20160
rect 59208 20095 59528 20096
rect 1853 20090 1919 20093
rect 0 20088 1919 20090
rect 0 20032 1858 20088
rect 1914 20032 1919 20088
rect 0 20030 1919 20032
rect 0 20000 800 20030
rect 1853 20027 1919 20030
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 14208 19616 14528 19617
rect 14208 19552 14216 19616
rect 14280 19552 14296 19616
rect 14360 19552 14376 19616
rect 14440 19552 14456 19616
rect 14520 19552 14528 19616
rect 14208 19551 14528 19552
rect 24208 19616 24528 19617
rect 24208 19552 24216 19616
rect 24280 19552 24296 19616
rect 24360 19552 24376 19616
rect 24440 19552 24456 19616
rect 24520 19552 24528 19616
rect 24208 19551 24528 19552
rect 34208 19616 34528 19617
rect 34208 19552 34216 19616
rect 34280 19552 34296 19616
rect 34360 19552 34376 19616
rect 34440 19552 34456 19616
rect 34520 19552 34528 19616
rect 34208 19551 34528 19552
rect 44208 19616 44528 19617
rect 44208 19552 44216 19616
rect 44280 19552 44296 19616
rect 44360 19552 44376 19616
rect 44440 19552 44456 19616
rect 44520 19552 44528 19616
rect 44208 19551 44528 19552
rect 54208 19616 54528 19617
rect 54208 19552 54216 19616
rect 54280 19552 54296 19616
rect 54360 19552 54376 19616
rect 54440 19552 54456 19616
rect 54520 19552 54528 19616
rect 54208 19551 54528 19552
rect 64208 19616 64528 19617
rect 64208 19552 64216 19616
rect 64280 19552 64296 19616
rect 64360 19552 64376 19616
rect 64440 19552 64456 19616
rect 64520 19552 64528 19616
rect 64208 19551 64528 19552
rect 68093 19138 68159 19141
rect 69200 19138 70000 19168
rect 68093 19136 70000 19138
rect 68093 19080 68098 19136
rect 68154 19080 70000 19136
rect 68093 19078 70000 19080
rect 68093 19075 68159 19078
rect 9208 19072 9528 19073
rect 9208 19008 9216 19072
rect 9280 19008 9296 19072
rect 9360 19008 9376 19072
rect 9440 19008 9456 19072
rect 9520 19008 9528 19072
rect 9208 19007 9528 19008
rect 39208 19072 39528 19073
rect 39208 19008 39216 19072
rect 39280 19008 39296 19072
rect 39360 19008 39376 19072
rect 39440 19008 39456 19072
rect 39520 19008 39528 19072
rect 39208 19007 39528 19008
rect 49208 19072 49528 19073
rect 49208 19008 49216 19072
rect 49280 19008 49296 19072
rect 49360 19008 49376 19072
rect 49440 19008 49456 19072
rect 49520 19008 49528 19072
rect 49208 19007 49528 19008
rect 59208 19072 59528 19073
rect 59208 19008 59216 19072
rect 59280 19008 59296 19072
rect 59360 19008 59376 19072
rect 59440 19008 59456 19072
rect 59520 19008 59528 19072
rect 69200 19048 70000 19078
rect 59208 19007 59528 19008
rect 0 18730 800 18760
rect 1761 18730 1827 18733
rect 0 18728 1827 18730
rect 0 18672 1766 18728
rect 1822 18672 1827 18728
rect 0 18670 1827 18672
rect 0 18640 800 18670
rect 1761 18667 1827 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 14208 18528 14528 18529
rect 14208 18464 14216 18528
rect 14280 18464 14296 18528
rect 14360 18464 14376 18528
rect 14440 18464 14456 18528
rect 14520 18464 14528 18528
rect 14208 18463 14528 18464
rect 44208 18528 44528 18529
rect 44208 18464 44216 18528
rect 44280 18464 44296 18528
rect 44360 18464 44376 18528
rect 44440 18464 44456 18528
rect 44520 18464 44528 18528
rect 44208 18463 44528 18464
rect 54208 18528 54528 18529
rect 54208 18464 54216 18528
rect 54280 18464 54296 18528
rect 54360 18464 54376 18528
rect 54440 18464 54456 18528
rect 54520 18464 54528 18528
rect 54208 18463 54528 18464
rect 64208 18528 64528 18529
rect 64208 18464 64216 18528
rect 64280 18464 64296 18528
rect 64360 18464 64376 18528
rect 64440 18464 64456 18528
rect 64520 18464 64528 18528
rect 64208 18463 64528 18464
rect 9208 17984 9528 17985
rect 9208 17920 9216 17984
rect 9280 17920 9296 17984
rect 9360 17920 9376 17984
rect 9440 17920 9456 17984
rect 9520 17920 9528 17984
rect 9208 17919 9528 17920
rect 39208 17984 39528 17985
rect 39208 17920 39216 17984
rect 39280 17920 39296 17984
rect 39360 17920 39376 17984
rect 39440 17920 39456 17984
rect 39520 17920 39528 17984
rect 39208 17919 39528 17920
rect 49208 17984 49528 17985
rect 49208 17920 49216 17984
rect 49280 17920 49296 17984
rect 49360 17920 49376 17984
rect 49440 17920 49456 17984
rect 49520 17920 49528 17984
rect 49208 17919 49528 17920
rect 59208 17984 59528 17985
rect 59208 17920 59216 17984
rect 59280 17920 59296 17984
rect 59360 17920 59376 17984
rect 59440 17920 59456 17984
rect 59520 17920 59528 17984
rect 59208 17919 59528 17920
rect 68093 17778 68159 17781
rect 69200 17778 70000 17808
rect 68093 17776 70000 17778
rect 68093 17720 68098 17776
rect 68154 17720 70000 17776
rect 68093 17718 70000 17720
rect 68093 17715 68159 17718
rect 69200 17688 70000 17718
rect 4208 17440 4528 17441
rect 0 17280 800 17400
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 14208 17440 14528 17441
rect 14208 17376 14216 17440
rect 14280 17376 14296 17440
rect 14360 17376 14376 17440
rect 14440 17376 14456 17440
rect 14520 17376 14528 17440
rect 14208 17375 14528 17376
rect 44208 17440 44528 17441
rect 44208 17376 44216 17440
rect 44280 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44528 17440
rect 44208 17375 44528 17376
rect 54208 17440 54528 17441
rect 54208 17376 54216 17440
rect 54280 17376 54296 17440
rect 54360 17376 54376 17440
rect 54440 17376 54456 17440
rect 54520 17376 54528 17440
rect 54208 17375 54528 17376
rect 64208 17440 64528 17441
rect 64208 17376 64216 17440
rect 64280 17376 64296 17440
rect 64360 17376 64376 17440
rect 64440 17376 64456 17440
rect 64520 17376 64528 17440
rect 64208 17375 64528 17376
rect 22093 17234 22159 17237
rect 39798 17234 39804 17236
rect 22093 17232 39804 17234
rect 22093 17176 22098 17232
rect 22154 17176 39804 17232
rect 22093 17174 39804 17176
rect 22093 17171 22159 17174
rect 39798 17172 39804 17174
rect 39868 17172 39874 17236
rect 9208 16896 9528 16897
rect 9208 16832 9216 16896
rect 9280 16832 9296 16896
rect 9360 16832 9376 16896
rect 9440 16832 9456 16896
rect 9520 16832 9528 16896
rect 9208 16831 9528 16832
rect 39208 16896 39528 16897
rect 39208 16832 39216 16896
rect 39280 16832 39296 16896
rect 39360 16832 39376 16896
rect 39440 16832 39456 16896
rect 39520 16832 39528 16896
rect 39208 16831 39528 16832
rect 49208 16896 49528 16897
rect 49208 16832 49216 16896
rect 49280 16832 49296 16896
rect 49360 16832 49376 16896
rect 49440 16832 49456 16896
rect 49520 16832 49528 16896
rect 49208 16831 49528 16832
rect 59208 16896 59528 16897
rect 59208 16832 59216 16896
rect 59280 16832 59296 16896
rect 59360 16832 59376 16896
rect 59440 16832 59456 16896
rect 59520 16832 59528 16896
rect 59208 16831 59528 16832
rect 29208 16438 29528 16476
rect 29208 16374 29216 16438
rect 29280 16374 29296 16438
rect 29360 16374 29376 16438
rect 29440 16374 29456 16438
rect 29520 16374 29528 16438
rect 29208 16358 29528 16374
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 14208 16352 14528 16353
rect 14208 16288 14216 16352
rect 14280 16288 14296 16352
rect 14360 16288 14376 16352
rect 14440 16288 14456 16352
rect 14520 16288 14528 16352
rect 14208 16287 14528 16288
rect 29208 16294 29216 16358
rect 29280 16294 29296 16358
rect 29360 16294 29376 16358
rect 29440 16294 29456 16358
rect 29520 16294 29528 16358
rect 68093 16418 68159 16421
rect 69200 16418 70000 16448
rect 68093 16416 70000 16418
rect 68093 16360 68098 16416
rect 68154 16360 70000 16416
rect 68093 16358 70000 16360
rect 68093 16355 68159 16358
rect 29208 16278 29528 16294
rect 44208 16352 44528 16353
rect 44208 16288 44216 16352
rect 44280 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44528 16352
rect 44208 16287 44528 16288
rect 54208 16352 54528 16353
rect 54208 16288 54216 16352
rect 54280 16288 54296 16352
rect 54360 16288 54376 16352
rect 54440 16288 54456 16352
rect 54520 16288 54528 16352
rect 54208 16287 54528 16288
rect 64208 16352 64528 16353
rect 64208 16288 64216 16352
rect 64280 16288 64296 16352
rect 64360 16288 64376 16352
rect 64440 16288 64456 16352
rect 64520 16288 64528 16352
rect 69200 16328 70000 16358
rect 64208 16287 64528 16288
rect 29208 16214 29216 16278
rect 29280 16214 29296 16278
rect 29360 16214 29376 16278
rect 29440 16214 29456 16278
rect 29520 16214 29528 16278
rect 29208 16198 29528 16214
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 29208 16134 29216 16198
rect 29280 16134 29296 16198
rect 29360 16134 29376 16198
rect 29440 16134 29456 16198
rect 29520 16134 29528 16198
rect 29208 16118 29528 16134
rect 29208 16054 29216 16118
rect 29280 16054 29296 16118
rect 29360 16054 29376 16118
rect 29440 16054 29456 16118
rect 29520 16054 29528 16118
rect 29208 16016 29528 16054
rect 9208 15808 9528 15809
rect 9208 15744 9216 15808
rect 9280 15744 9296 15808
rect 9360 15744 9376 15808
rect 9440 15744 9456 15808
rect 9520 15744 9528 15808
rect 9208 15743 9528 15744
rect 39208 15808 39528 15809
rect 39208 15744 39216 15808
rect 39280 15744 39296 15808
rect 39360 15744 39376 15808
rect 39440 15744 39456 15808
rect 39520 15744 39528 15808
rect 39208 15743 39528 15744
rect 49208 15808 49528 15809
rect 49208 15744 49216 15808
rect 49280 15744 49296 15808
rect 49360 15744 49376 15808
rect 49440 15744 49456 15808
rect 49520 15744 49528 15808
rect 49208 15743 49528 15744
rect 59208 15808 59528 15809
rect 59208 15744 59216 15808
rect 59280 15744 59296 15808
rect 59360 15744 59376 15808
rect 59440 15744 59456 15808
rect 59520 15744 59528 15808
rect 59208 15743 59528 15744
rect 24208 15638 24528 15676
rect 24208 15574 24216 15638
rect 24280 15574 24296 15638
rect 24360 15574 24376 15638
rect 24440 15574 24456 15638
rect 24520 15574 24528 15638
rect 24208 15558 24528 15574
rect 24208 15494 24216 15558
rect 24280 15494 24296 15558
rect 24360 15494 24376 15558
rect 24440 15494 24456 15558
rect 24520 15494 24528 15558
rect 24208 15478 24528 15494
rect 24208 15414 24216 15478
rect 24280 15414 24296 15478
rect 24360 15414 24376 15478
rect 24440 15414 24456 15478
rect 24520 15414 24528 15478
rect 24208 15398 24528 15414
rect 24208 15334 24216 15398
rect 24280 15334 24296 15398
rect 24360 15334 24376 15398
rect 24440 15334 24456 15398
rect 24520 15334 24528 15398
rect 24208 15318 24528 15334
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 14208 15264 14528 15265
rect 14208 15200 14216 15264
rect 14280 15200 14296 15264
rect 14360 15200 14376 15264
rect 14440 15200 14456 15264
rect 14520 15200 14528 15264
rect 24208 15254 24216 15318
rect 24280 15254 24296 15318
rect 24360 15254 24376 15318
rect 24440 15254 24456 15318
rect 24520 15254 24528 15318
rect 24208 15216 24528 15254
rect 44208 15264 44528 15265
rect 14208 15199 14528 15200
rect 44208 15200 44216 15264
rect 44280 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44528 15264
rect 44208 15199 44528 15200
rect 54208 15264 54528 15265
rect 54208 15200 54216 15264
rect 54280 15200 54296 15264
rect 54360 15200 54376 15264
rect 54440 15200 54456 15264
rect 54520 15200 54528 15264
rect 54208 15199 54528 15200
rect 64208 15264 64528 15265
rect 64208 15200 64216 15264
rect 64280 15200 64296 15264
rect 64360 15200 64376 15264
rect 64440 15200 64456 15264
rect 64520 15200 64528 15264
rect 64208 15199 64528 15200
rect 68093 15058 68159 15061
rect 69200 15058 70000 15088
rect 68093 15056 70000 15058
rect 68093 15000 68098 15056
rect 68154 15000 70000 15056
rect 68093 14998 70000 15000
rect 68093 14995 68159 14998
rect 69200 14968 70000 14998
rect 0 14786 800 14816
rect 1853 14786 1919 14789
rect 0 14784 1919 14786
rect 0 14728 1858 14784
rect 1914 14728 1919 14784
rect 0 14726 1919 14728
rect 0 14696 800 14726
rect 1853 14723 1919 14726
rect 9208 14720 9528 14721
rect 9208 14656 9216 14720
rect 9280 14656 9296 14720
rect 9360 14656 9376 14720
rect 9440 14656 9456 14720
rect 9520 14656 9528 14720
rect 9208 14655 9528 14656
rect 39208 14720 39528 14721
rect 39208 14656 39216 14720
rect 39280 14656 39296 14720
rect 39360 14656 39376 14720
rect 39440 14656 39456 14720
rect 39520 14656 39528 14720
rect 39208 14655 39528 14656
rect 49208 14720 49528 14721
rect 49208 14656 49216 14720
rect 49280 14656 49296 14720
rect 49360 14656 49376 14720
rect 49440 14656 49456 14720
rect 49520 14656 49528 14720
rect 49208 14655 49528 14656
rect 59208 14720 59528 14721
rect 59208 14656 59216 14720
rect 59280 14656 59296 14720
rect 59360 14656 59376 14720
rect 59440 14656 59456 14720
rect 59520 14656 59528 14720
rect 59208 14655 59528 14656
rect 40166 14452 40172 14516
rect 40236 14514 40242 14516
rect 41505 14514 41571 14517
rect 40236 14512 41571 14514
rect 40236 14456 41510 14512
rect 41566 14456 41571 14512
rect 40236 14454 41571 14456
rect 40236 14452 40242 14454
rect 41505 14451 41571 14454
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 14208 14176 14528 14177
rect 14208 14112 14216 14176
rect 14280 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14528 14176
rect 14208 14111 14528 14112
rect 44208 14176 44528 14177
rect 44208 14112 44216 14176
rect 44280 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44528 14176
rect 44208 14111 44528 14112
rect 54208 14176 54528 14177
rect 54208 14112 54216 14176
rect 54280 14112 54296 14176
rect 54360 14112 54376 14176
rect 54440 14112 54456 14176
rect 54520 14112 54528 14176
rect 54208 14111 54528 14112
rect 64208 14176 64528 14177
rect 64208 14112 64216 14176
rect 64280 14112 64296 14176
rect 64360 14112 64376 14176
rect 64440 14112 64456 14176
rect 64520 14112 64528 14176
rect 64208 14111 64528 14112
rect 15694 13772 15700 13836
rect 15764 13834 15770 13836
rect 15837 13834 15903 13837
rect 16297 13836 16363 13837
rect 15764 13832 15903 13834
rect 15764 13776 15842 13832
rect 15898 13776 15903 13832
rect 15764 13774 15903 13776
rect 15764 13772 15770 13774
rect 15837 13771 15903 13774
rect 16246 13772 16252 13836
rect 16316 13834 16363 13836
rect 68093 13834 68159 13837
rect 69200 13834 70000 13864
rect 16316 13832 16408 13834
rect 16358 13776 16408 13832
rect 16316 13774 16408 13776
rect 68093 13832 70000 13834
rect 68093 13776 68098 13832
rect 68154 13776 70000 13832
rect 68093 13774 70000 13776
rect 16316 13772 16363 13774
rect 16297 13771 16363 13772
rect 68093 13771 68159 13774
rect 69200 13744 70000 13774
rect 9208 13632 9528 13633
rect 0 13562 800 13592
rect 9208 13568 9216 13632
rect 9280 13568 9296 13632
rect 9360 13568 9376 13632
rect 9440 13568 9456 13632
rect 9520 13568 9528 13632
rect 9208 13567 9528 13568
rect 39208 13632 39528 13633
rect 39208 13568 39216 13632
rect 39280 13568 39296 13632
rect 39360 13568 39376 13632
rect 39440 13568 39456 13632
rect 39520 13568 39528 13632
rect 39208 13567 39528 13568
rect 49208 13632 49528 13633
rect 49208 13568 49216 13632
rect 49280 13568 49296 13632
rect 49360 13568 49376 13632
rect 49440 13568 49456 13632
rect 49520 13568 49528 13632
rect 49208 13567 49528 13568
rect 59208 13632 59528 13633
rect 59208 13568 59216 13632
rect 59280 13568 59296 13632
rect 59360 13568 59376 13632
rect 59440 13568 59456 13632
rect 59520 13568 59528 13632
rect 59208 13567 59528 13568
rect 1853 13562 1919 13565
rect 0 13560 1919 13562
rect 0 13504 1858 13560
rect 1914 13504 1919 13560
rect 0 13502 1919 13504
rect 0 13472 800 13502
rect 1853 13499 1919 13502
rect 13537 13156 13603 13157
rect 13486 13092 13492 13156
rect 13556 13154 13603 13156
rect 13556 13152 13648 13154
rect 13598 13096 13648 13152
rect 13556 13094 13648 13096
rect 13556 13092 13603 13094
rect 39062 13092 39068 13156
rect 39132 13154 39138 13156
rect 39205 13154 39271 13157
rect 39132 13152 39271 13154
rect 39132 13096 39210 13152
rect 39266 13096 39271 13152
rect 39132 13094 39271 13096
rect 39132 13092 39138 13094
rect 13537 13091 13603 13092
rect 39205 13091 39271 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 14208 13088 14528 13089
rect 14208 13024 14216 13088
rect 14280 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14528 13088
rect 14208 13023 14528 13024
rect 44208 13088 44528 13089
rect 44208 13024 44216 13088
rect 44280 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44528 13088
rect 44208 13023 44528 13024
rect 54208 13088 54528 13089
rect 54208 13024 54216 13088
rect 54280 13024 54296 13088
rect 54360 13024 54376 13088
rect 54440 13024 54456 13088
rect 54520 13024 54528 13088
rect 54208 13023 54528 13024
rect 64208 13088 64528 13089
rect 64208 13024 64216 13088
rect 64280 13024 64296 13088
rect 64360 13024 64376 13088
rect 64440 13024 64456 13088
rect 64520 13024 64528 13088
rect 64208 13023 64528 13024
rect 39798 12956 39804 13020
rect 39868 13018 39874 13020
rect 39941 13018 40007 13021
rect 39868 13016 40007 13018
rect 39868 12960 39946 13016
rect 40002 12960 40007 13016
rect 39868 12958 40007 12960
rect 39868 12956 39874 12958
rect 39941 12955 40007 12958
rect 13118 12548 13124 12612
rect 13188 12610 13194 12612
rect 13353 12610 13419 12613
rect 13188 12608 13419 12610
rect 13188 12552 13358 12608
rect 13414 12552 13419 12608
rect 13188 12550 13419 12552
rect 13188 12548 13194 12550
rect 13353 12547 13419 12550
rect 40718 12548 40724 12612
rect 40788 12610 40794 12612
rect 40861 12610 40927 12613
rect 40788 12608 40927 12610
rect 40788 12552 40866 12608
rect 40922 12552 40927 12608
rect 40788 12550 40927 12552
rect 40788 12548 40794 12550
rect 40861 12547 40927 12550
rect 9208 12544 9528 12545
rect 9208 12480 9216 12544
rect 9280 12480 9296 12544
rect 9360 12480 9376 12544
rect 9440 12480 9456 12544
rect 9520 12480 9528 12544
rect 9208 12479 9528 12480
rect 39208 12544 39528 12545
rect 39208 12480 39216 12544
rect 39280 12480 39296 12544
rect 39360 12480 39376 12544
rect 39440 12480 39456 12544
rect 39520 12480 39528 12544
rect 39208 12479 39528 12480
rect 49208 12544 49528 12545
rect 49208 12480 49216 12544
rect 49280 12480 49296 12544
rect 49360 12480 49376 12544
rect 49440 12480 49456 12544
rect 49520 12480 49528 12544
rect 49208 12479 49528 12480
rect 59208 12544 59528 12545
rect 59208 12480 59216 12544
rect 59280 12480 59296 12544
rect 59360 12480 59376 12544
rect 59440 12480 59456 12544
rect 59520 12480 59528 12544
rect 59208 12479 59528 12480
rect 39614 12412 39620 12476
rect 39684 12474 39690 12476
rect 39757 12474 39823 12477
rect 39684 12472 39823 12474
rect 39684 12416 39762 12472
rect 39818 12416 39823 12472
rect 39684 12414 39823 12416
rect 39684 12412 39690 12414
rect 39757 12411 39823 12414
rect 68093 12474 68159 12477
rect 69200 12474 70000 12504
rect 68093 12472 70000 12474
rect 68093 12416 68098 12472
rect 68154 12416 70000 12472
rect 68093 12414 70000 12416
rect 68093 12411 68159 12414
rect 69200 12384 70000 12414
rect 17493 12338 17559 12341
rect 46933 12338 46999 12341
rect 17493 12336 46999 12338
rect 17493 12280 17498 12336
rect 17554 12280 46938 12336
rect 46994 12280 46999 12336
rect 17493 12278 46999 12280
rect 17493 12275 17559 12278
rect 46933 12275 46999 12278
rect 0 12112 800 12232
rect 13905 12202 13971 12205
rect 37917 12202 37983 12205
rect 39757 12204 39823 12205
rect 13905 12200 37983 12202
rect 13905 12144 13910 12200
rect 13966 12144 37922 12200
rect 37978 12144 37983 12200
rect 13905 12142 37983 12144
rect 13905 12139 13971 12142
rect 37917 12139 37983 12142
rect 38694 12140 38700 12204
rect 38764 12202 38770 12204
rect 39757 12202 39804 12204
rect 38764 12200 39804 12202
rect 38764 12144 39762 12200
rect 38764 12142 39804 12144
rect 38764 12140 38770 12142
rect 39757 12140 39804 12142
rect 39868 12140 39874 12204
rect 39757 12139 39823 12140
rect 16113 12066 16179 12069
rect 38285 12066 38351 12069
rect 16113 12064 38351 12066
rect 16113 12008 16118 12064
rect 16174 12008 38290 12064
rect 38346 12008 38351 12064
rect 16113 12006 38351 12008
rect 16113 12003 16179 12006
rect 38285 12003 38351 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 14208 12000 14528 12001
rect 14208 11936 14216 12000
rect 14280 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14528 12000
rect 14208 11935 14528 11936
rect 44208 12000 44528 12001
rect 44208 11936 44216 12000
rect 44280 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44528 12000
rect 44208 11935 44528 11936
rect 54208 12000 54528 12001
rect 54208 11936 54216 12000
rect 54280 11936 54296 12000
rect 54360 11936 54376 12000
rect 54440 11936 54456 12000
rect 54520 11936 54528 12000
rect 54208 11935 54528 11936
rect 64208 12000 64528 12001
rect 64208 11936 64216 12000
rect 64280 11936 64296 12000
rect 64360 11936 64376 12000
rect 64440 11936 64456 12000
rect 64520 11936 64528 12000
rect 64208 11935 64528 11936
rect 24208 11907 24528 11935
rect 24208 11843 24216 11907
rect 24280 11843 24296 11907
rect 24360 11843 24376 11907
rect 24440 11843 24456 11907
rect 24520 11843 24528 11907
rect 24208 11827 24528 11843
rect 24208 11763 24216 11827
rect 24280 11763 24296 11827
rect 24360 11763 24376 11827
rect 24440 11763 24456 11827
rect 24520 11763 24528 11827
rect 24208 11747 24528 11763
rect 24208 11683 24216 11747
rect 24280 11683 24296 11747
rect 24360 11683 24376 11747
rect 24440 11683 24456 11747
rect 24520 11683 24528 11747
rect 24208 11667 24528 11683
rect 14825 11660 14891 11661
rect 14774 11596 14780 11660
rect 14844 11658 14891 11660
rect 14844 11656 14936 11658
rect 14886 11600 14936 11656
rect 14844 11598 14936 11600
rect 24208 11603 24216 11667
rect 24280 11603 24296 11667
rect 24360 11603 24376 11667
rect 24440 11603 24456 11667
rect 24520 11603 24528 11667
rect 14844 11596 14891 11598
rect 14825 11595 14891 11596
rect 24208 11575 24528 11603
rect 34208 11907 34528 11935
rect 34208 11843 34216 11907
rect 34280 11843 34296 11907
rect 34360 11843 34376 11907
rect 34440 11843 34456 11907
rect 34520 11843 34528 11907
rect 34208 11827 34528 11843
rect 34208 11763 34216 11827
rect 34280 11763 34296 11827
rect 34360 11763 34376 11827
rect 34440 11763 34456 11827
rect 34520 11763 34528 11827
rect 34208 11747 34528 11763
rect 34208 11683 34216 11747
rect 34280 11683 34296 11747
rect 34360 11683 34376 11747
rect 34440 11683 34456 11747
rect 34520 11683 34528 11747
rect 34208 11667 34528 11683
rect 34208 11603 34216 11667
rect 34280 11603 34296 11667
rect 34360 11603 34376 11667
rect 34440 11603 34456 11667
rect 34520 11603 34528 11667
rect 34208 11575 34528 11603
rect 9208 11456 9528 11457
rect 9208 11392 9216 11456
rect 9280 11392 9296 11456
rect 9360 11392 9376 11456
rect 9440 11392 9456 11456
rect 9520 11392 9528 11456
rect 9208 11391 9528 11392
rect 39208 11456 39528 11457
rect 39208 11392 39216 11456
rect 39280 11392 39296 11456
rect 39360 11392 39376 11456
rect 39440 11392 39456 11456
rect 39520 11392 39528 11456
rect 39208 11391 39528 11392
rect 49208 11456 49528 11457
rect 49208 11392 49216 11456
rect 49280 11392 49296 11456
rect 49360 11392 49376 11456
rect 49440 11392 49456 11456
rect 49520 11392 49528 11456
rect 49208 11391 49528 11392
rect 59208 11456 59528 11457
rect 59208 11392 59216 11456
rect 59280 11392 59296 11456
rect 59360 11392 59376 11456
rect 59440 11392 59456 11456
rect 59520 11392 59528 11456
rect 59208 11391 59528 11392
rect 13813 11388 13879 11389
rect 13813 11386 13860 11388
rect 13768 11384 13860 11386
rect 13768 11328 13818 11384
rect 13768 11326 13860 11328
rect 13813 11324 13860 11326
rect 13924 11324 13930 11388
rect 39665 11386 39731 11389
rect 43805 11386 43871 11389
rect 39665 11384 43871 11386
rect 39665 11328 39670 11384
rect 39726 11328 43810 11384
rect 43866 11328 43871 11384
rect 39665 11326 43871 11328
rect 13813 11323 13879 11324
rect 39665 11323 39731 11326
rect 43805 11323 43871 11326
rect 9673 11252 9739 11253
rect 9622 11188 9628 11252
rect 9692 11250 9739 11252
rect 18321 11250 18387 11253
rect 45369 11250 45435 11253
rect 9692 11248 9784 11250
rect 9734 11192 9784 11248
rect 9692 11190 9784 11192
rect 18321 11248 45435 11250
rect 18321 11192 18326 11248
rect 18382 11192 45374 11248
rect 45430 11192 45435 11248
rect 18321 11190 45435 11192
rect 9692 11188 9739 11190
rect 9673 11187 9739 11188
rect 18321 11187 18387 11190
rect 45369 11187 45435 11190
rect 2681 11114 2747 11117
rect 39665 11114 39731 11117
rect 2681 11112 39731 11114
rect 2681 11056 2686 11112
rect 2742 11056 39670 11112
rect 39726 11056 39731 11112
rect 2681 11054 39731 11056
rect 2681 11051 2747 11054
rect 39665 11051 39731 11054
rect 42333 11114 42399 11117
rect 42558 11114 42564 11116
rect 42333 11112 42564 11114
rect 42333 11056 42338 11112
rect 42394 11056 42564 11112
rect 42333 11054 42564 11056
rect 42333 11051 42399 11054
rect 42558 11052 42564 11054
rect 42628 11114 42634 11116
rect 42701 11114 42767 11117
rect 42628 11112 42767 11114
rect 42628 11056 42706 11112
rect 42762 11056 42767 11112
rect 42628 11054 42767 11056
rect 42628 11052 42634 11054
rect 42701 11051 42767 11054
rect 68093 11114 68159 11117
rect 69200 11114 70000 11144
rect 68093 11112 70000 11114
rect 68093 11056 68098 11112
rect 68154 11056 70000 11112
rect 68093 11054 70000 11056
rect 68093 11051 68159 11054
rect 69200 11024 70000 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 44081 10978 44147 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 17174 10976 44147 10978
rect 17174 10920 44086 10976
rect 44142 10920 44147 10976
rect 17174 10918 44147 10920
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 14208 10912 14528 10913
rect 14208 10848 14216 10912
rect 14280 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14528 10912
rect 14208 10847 14528 10848
rect 9949 10706 10015 10709
rect 17174 10706 17234 10918
rect 44081 10915 44147 10918
rect 44208 10912 44528 10913
rect 44208 10848 44216 10912
rect 44280 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44528 10912
rect 44208 10847 44528 10848
rect 54208 10912 54528 10913
rect 54208 10848 54216 10912
rect 54280 10848 54296 10912
rect 54360 10848 54376 10912
rect 54440 10848 54456 10912
rect 54520 10848 54528 10912
rect 54208 10847 54528 10848
rect 64208 10912 64528 10913
rect 64208 10848 64216 10912
rect 64280 10848 64296 10912
rect 64360 10848 64376 10912
rect 64440 10848 64456 10912
rect 64520 10848 64528 10912
rect 64208 10847 64528 10848
rect 18229 10842 18295 10845
rect 41965 10842 42031 10845
rect 18229 10840 42031 10842
rect 18229 10784 18234 10840
rect 18290 10784 41970 10840
rect 42026 10784 42031 10840
rect 18229 10782 42031 10784
rect 18229 10779 18295 10782
rect 41965 10779 42031 10782
rect 9949 10704 17234 10706
rect 9949 10648 9954 10704
rect 10010 10648 17234 10704
rect 9949 10646 17234 10648
rect 9949 10643 10015 10646
rect 29208 10633 29528 10661
rect 14457 10570 14523 10573
rect 14774 10570 14780 10572
rect 14457 10568 14780 10570
rect 14457 10512 14462 10568
rect 14518 10512 14780 10568
rect 14457 10510 14780 10512
rect 14457 10507 14523 10510
rect 14774 10508 14780 10510
rect 14844 10508 14850 10572
rect 29208 10569 29216 10633
rect 29280 10569 29296 10633
rect 29360 10569 29376 10633
rect 29440 10569 29456 10633
rect 29520 10569 29528 10633
rect 29208 10553 29528 10569
rect 29208 10489 29216 10553
rect 29280 10489 29296 10553
rect 29360 10489 29376 10553
rect 29440 10489 29456 10553
rect 29520 10489 29528 10553
rect 40125 10570 40191 10573
rect 40350 10570 40356 10572
rect 40125 10568 40356 10570
rect 40125 10512 40130 10568
rect 40186 10512 40356 10568
rect 40125 10510 40356 10512
rect 40125 10507 40191 10510
rect 40350 10508 40356 10510
rect 40420 10508 40426 10572
rect 29208 10473 29528 10489
rect 29208 10409 29216 10473
rect 29280 10409 29296 10473
rect 29360 10409 29376 10473
rect 29440 10409 29456 10473
rect 29520 10409 29528 10473
rect 29208 10393 29528 10409
rect 9208 10368 9528 10369
rect 9208 10304 9216 10368
rect 9280 10304 9296 10368
rect 9360 10304 9376 10368
rect 9440 10304 9456 10368
rect 9520 10304 9528 10368
rect 9208 10303 9528 10304
rect 29208 10329 29216 10393
rect 29280 10329 29296 10393
rect 29360 10329 29376 10393
rect 29440 10329 29456 10393
rect 29520 10329 29528 10393
rect 29208 10301 29528 10329
rect 39208 10368 39528 10369
rect 39208 10304 39216 10368
rect 39280 10304 39296 10368
rect 39360 10304 39376 10368
rect 39440 10304 39456 10368
rect 39520 10304 39528 10368
rect 39208 10303 39528 10304
rect 49208 10368 49528 10369
rect 49208 10304 49216 10368
rect 49280 10304 49296 10368
rect 49360 10304 49376 10368
rect 49440 10304 49456 10368
rect 49520 10304 49528 10368
rect 49208 10303 49528 10304
rect 59208 10368 59528 10369
rect 59208 10304 59216 10368
rect 59280 10304 59296 10368
rect 59360 10304 59376 10368
rect 59440 10304 59456 10368
rect 59520 10304 59528 10368
rect 59208 10303 59528 10304
rect 14825 10298 14891 10301
rect 14825 10296 15210 10298
rect 14825 10240 14830 10296
rect 14886 10240 15210 10296
rect 14825 10238 15210 10240
rect 14825 10235 14891 10238
rect 14733 10162 14799 10165
rect 14733 10160 14842 10162
rect 14733 10104 14738 10160
rect 14794 10104 14842 10160
rect 14733 10099 14842 10104
rect 11605 10028 11671 10029
rect 11605 10026 11652 10028
rect 11560 10024 11652 10026
rect 11560 9968 11610 10024
rect 11560 9966 11652 9968
rect 11605 9964 11652 9966
rect 11716 9964 11722 10028
rect 14549 10026 14615 10029
rect 14549 10024 14658 10026
rect 14549 9968 14554 10024
rect 14610 9968 14658 10024
rect 11605 9963 11671 9964
rect 14549 9963 14658 9968
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 14208 9824 14528 9825
rect 14208 9760 14216 9824
rect 14280 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14528 9824
rect 14208 9759 14528 9760
rect 14365 9690 14431 9693
rect 14598 9690 14658 9963
rect 14782 9693 14842 10099
rect 15150 10029 15210 10238
rect 15150 10024 15259 10029
rect 40861 10026 40927 10029
rect 15150 9968 15198 10024
rect 15254 9968 15259 10024
rect 15150 9966 15259 9968
rect 15193 9963 15259 9966
rect 40542 10024 40927 10026
rect 40542 9968 40866 10024
rect 40922 9968 40927 10024
rect 40542 9966 40927 9968
rect 14365 9688 14658 9690
rect 0 9618 800 9648
rect 14365 9632 14370 9688
rect 14426 9632 14658 9688
rect 14365 9630 14658 9632
rect 14733 9688 14842 9693
rect 14733 9632 14738 9688
rect 14794 9632 14842 9688
rect 14733 9630 14842 9632
rect 14365 9627 14431 9630
rect 14733 9627 14799 9630
rect 1761 9618 1827 9621
rect 0 9616 1827 9618
rect 0 9560 1766 9616
rect 1822 9560 1827 9616
rect 0 9558 1827 9560
rect 0 9528 800 9558
rect 1761 9555 1827 9558
rect 16205 9482 16271 9485
rect 16205 9480 16314 9482
rect 16205 9424 16210 9480
rect 16266 9424 16314 9480
rect 16205 9419 16314 9424
rect 38878 9420 38884 9484
rect 38948 9482 38954 9484
rect 39481 9482 39547 9485
rect 38948 9480 39547 9482
rect 38948 9424 39486 9480
rect 39542 9424 39547 9480
rect 38948 9422 39547 9424
rect 38948 9420 38954 9422
rect 39481 9419 39547 9422
rect 14774 9284 14780 9348
rect 14844 9346 14850 9348
rect 14917 9346 14983 9349
rect 14844 9344 14983 9346
rect 14844 9288 14922 9344
rect 14978 9288 14983 9344
rect 14844 9286 14983 9288
rect 14844 9284 14850 9286
rect 14917 9283 14983 9286
rect 9208 9280 9528 9281
rect 9208 9216 9216 9280
rect 9280 9216 9296 9280
rect 9360 9216 9376 9280
rect 9440 9216 9456 9280
rect 9520 9216 9528 9280
rect 9208 9215 9528 9216
rect 14089 9076 14155 9077
rect 14038 9012 14044 9076
rect 14108 9074 14155 9076
rect 14108 9072 14200 9074
rect 14150 9016 14200 9072
rect 14108 9014 14200 9016
rect 14108 9012 14155 9014
rect 14089 9011 14155 9012
rect 14365 8938 14431 8941
rect 14590 8938 14596 8940
rect 14365 8936 14596 8938
rect 14365 8880 14370 8936
rect 14426 8880 14596 8936
rect 14365 8878 14596 8880
rect 14365 8875 14431 8878
rect 14590 8876 14596 8878
rect 14660 8876 14666 8940
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 14208 8736 14528 8737
rect 14208 8672 14216 8736
rect 14280 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14528 8736
rect 14208 8671 14528 8672
rect 12249 8532 12315 8533
rect 12198 8468 12204 8532
rect 12268 8530 12315 8532
rect 12268 8528 12360 8530
rect 12310 8472 12360 8528
rect 12268 8470 12360 8472
rect 12268 8468 12315 8470
rect 12249 8467 12315 8468
rect 0 8394 800 8424
rect 16254 8397 16314 9419
rect 24208 9358 24528 9386
rect 24208 9294 24216 9358
rect 24280 9294 24296 9358
rect 24360 9294 24376 9358
rect 24440 9294 24456 9358
rect 24520 9294 24528 9358
rect 24208 9278 24528 9294
rect 24208 9214 24216 9278
rect 24280 9214 24296 9278
rect 24360 9214 24376 9278
rect 24440 9214 24456 9278
rect 24520 9214 24528 9278
rect 24208 9198 24528 9214
rect 24208 9134 24216 9198
rect 24280 9134 24296 9198
rect 24360 9134 24376 9198
rect 24440 9134 24456 9198
rect 24520 9134 24528 9198
rect 24208 9118 24528 9134
rect 17217 9074 17283 9077
rect 17217 9072 17418 9074
rect 17217 9016 17222 9072
rect 17278 9016 17418 9072
rect 24208 9054 24216 9118
rect 24280 9054 24296 9118
rect 24360 9054 24376 9118
rect 24440 9054 24456 9118
rect 24520 9054 24528 9118
rect 24208 9026 24528 9054
rect 34208 9358 34528 9386
rect 34208 9294 34216 9358
rect 34280 9294 34296 9358
rect 34360 9294 34376 9358
rect 34440 9294 34456 9358
rect 34520 9294 34528 9358
rect 34208 9278 34528 9294
rect 34208 9214 34216 9278
rect 34280 9214 34296 9278
rect 34360 9214 34376 9278
rect 34440 9214 34456 9278
rect 34520 9214 34528 9278
rect 39208 9280 39528 9281
rect 39208 9216 39216 9280
rect 39280 9216 39296 9280
rect 39360 9216 39376 9280
rect 39440 9216 39456 9280
rect 39520 9216 39528 9280
rect 39208 9215 39528 9216
rect 34208 9198 34528 9214
rect 40542 9213 40602 9966
rect 40861 9963 40927 9966
rect 68093 9890 68159 9893
rect 69200 9890 70000 9920
rect 68093 9888 70000 9890
rect 68093 9832 68098 9888
rect 68154 9832 70000 9888
rect 68093 9830 70000 9832
rect 68093 9827 68159 9830
rect 44208 9824 44528 9825
rect 44208 9760 44216 9824
rect 44280 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44528 9824
rect 44208 9759 44528 9760
rect 54208 9824 54528 9825
rect 54208 9760 54216 9824
rect 54280 9760 54296 9824
rect 54360 9760 54376 9824
rect 54440 9760 54456 9824
rect 54520 9760 54528 9824
rect 54208 9759 54528 9760
rect 64208 9824 64528 9825
rect 64208 9760 64216 9824
rect 64280 9760 64296 9824
rect 64360 9760 64376 9824
rect 64440 9760 64456 9824
rect 64520 9760 64528 9824
rect 69200 9800 70000 9830
rect 64208 9759 64528 9760
rect 43846 9420 43852 9484
rect 43916 9482 43922 9484
rect 43989 9482 44055 9485
rect 43916 9480 44055 9482
rect 43916 9424 43994 9480
rect 44050 9424 44055 9480
rect 43916 9422 44055 9424
rect 43916 9420 43922 9422
rect 43989 9419 44055 9422
rect 49208 9280 49528 9281
rect 49208 9216 49216 9280
rect 49280 9216 49296 9280
rect 49360 9216 49376 9280
rect 49440 9216 49456 9280
rect 49520 9216 49528 9280
rect 49208 9215 49528 9216
rect 59208 9280 59528 9281
rect 59208 9216 59216 9280
rect 59280 9216 59296 9280
rect 59360 9216 59376 9280
rect 59440 9216 59456 9280
rect 59520 9216 59528 9280
rect 59208 9215 59528 9216
rect 34208 9134 34216 9198
rect 34280 9134 34296 9198
rect 34360 9134 34376 9198
rect 34440 9134 34456 9198
rect 34520 9134 34528 9198
rect 40493 9208 40602 9213
rect 40493 9152 40498 9208
rect 40554 9152 40602 9208
rect 40493 9150 40602 9152
rect 40493 9147 40559 9150
rect 40902 9148 40908 9212
rect 40972 9210 40978 9212
rect 43621 9210 43687 9213
rect 40972 9208 43687 9210
rect 40972 9152 43626 9208
rect 43682 9152 43687 9208
rect 40972 9150 43687 9152
rect 40972 9148 40978 9150
rect 43621 9147 43687 9150
rect 34208 9118 34528 9134
rect 34208 9054 34216 9118
rect 34280 9054 34296 9118
rect 34360 9054 34376 9118
rect 34440 9054 34456 9118
rect 34520 9054 34528 9118
rect 34208 9026 34528 9054
rect 39021 9074 39087 9077
rect 40166 9074 40172 9076
rect 39021 9072 40172 9074
rect 17217 9014 17418 9016
rect 17217 9011 17283 9014
rect 17358 8802 17418 9014
rect 39021 9016 39026 9072
rect 39082 9016 40172 9072
rect 39021 9014 40172 9016
rect 39021 9011 39087 9014
rect 40166 9012 40172 9014
rect 40236 9012 40242 9076
rect 41454 9012 41460 9076
rect 41524 9074 41530 9076
rect 42885 9074 42951 9077
rect 41524 9072 42951 9074
rect 41524 9016 42890 9072
rect 42946 9016 42951 9072
rect 41524 9014 42951 9016
rect 41524 9012 41530 9014
rect 42885 9011 42951 9014
rect 39849 8938 39915 8941
rect 42333 8940 42399 8941
rect 39982 8938 39988 8940
rect 39849 8936 39988 8938
rect 39849 8880 39854 8936
rect 39910 8880 39988 8936
rect 39849 8878 39988 8880
rect 39849 8875 39915 8878
rect 39982 8876 39988 8878
rect 40052 8876 40058 8940
rect 42333 8936 42380 8940
rect 42444 8938 42450 8940
rect 42333 8880 42338 8936
rect 42333 8876 42380 8880
rect 42444 8878 42490 8938
rect 42444 8876 42450 8878
rect 44030 8876 44036 8940
rect 44100 8938 44106 8940
rect 44265 8938 44331 8941
rect 44100 8936 44331 8938
rect 44100 8880 44270 8936
rect 44326 8880 44331 8936
rect 44100 8878 44331 8880
rect 44100 8876 44106 8878
rect 42333 8875 42399 8876
rect 44265 8875 44331 8878
rect 17493 8802 17559 8805
rect 17358 8800 17559 8802
rect 17358 8744 17498 8800
rect 17554 8744 17559 8800
rect 17358 8742 17559 8744
rect 17493 8739 17559 8742
rect 44208 8736 44528 8737
rect 44208 8672 44216 8736
rect 44280 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44528 8736
rect 44208 8671 44528 8672
rect 54208 8736 54528 8737
rect 54208 8672 54216 8736
rect 54280 8672 54296 8736
rect 54360 8672 54376 8736
rect 54440 8672 54456 8736
rect 54520 8672 54528 8736
rect 54208 8671 54528 8672
rect 64208 8736 64528 8737
rect 64208 8672 64216 8736
rect 64280 8672 64296 8736
rect 64360 8672 64376 8736
rect 64440 8672 64456 8736
rect 64520 8672 64528 8736
rect 64208 8671 64528 8672
rect 39389 8530 39455 8533
rect 40350 8530 40356 8532
rect 39389 8528 40356 8530
rect 39389 8472 39394 8528
rect 39450 8472 40356 8528
rect 39389 8470 40356 8472
rect 39389 8467 39455 8470
rect 40350 8468 40356 8470
rect 40420 8468 40426 8532
rect 44950 8468 44956 8532
rect 45020 8530 45026 8532
rect 45093 8530 45159 8533
rect 45020 8528 45159 8530
rect 45020 8472 45098 8528
rect 45154 8472 45159 8528
rect 45020 8470 45159 8472
rect 45020 8468 45026 8470
rect 45093 8467 45159 8470
rect 68093 8530 68159 8533
rect 69200 8530 70000 8560
rect 68093 8528 70000 8530
rect 68093 8472 68098 8528
rect 68154 8472 70000 8528
rect 68093 8470 70000 8472
rect 68093 8467 68159 8470
rect 69200 8440 70000 8470
rect 1761 8394 1827 8397
rect 0 8392 1827 8394
rect 0 8336 1766 8392
rect 1822 8336 1827 8392
rect 0 8334 1827 8336
rect 16254 8392 16363 8397
rect 16254 8336 16302 8392
rect 16358 8336 16363 8392
rect 16254 8334 16363 8336
rect 0 8304 800 8334
rect 1761 8331 1827 8334
rect 16297 8331 16363 8334
rect 41321 8260 41387 8261
rect 41270 8196 41276 8260
rect 41340 8258 41387 8260
rect 41340 8256 41432 8258
rect 41382 8200 41432 8256
rect 41340 8198 41432 8200
rect 41340 8196 41387 8198
rect 41321 8195 41387 8196
rect 9208 8192 9528 8193
rect 9208 8128 9216 8192
rect 9280 8128 9296 8192
rect 9360 8128 9376 8192
rect 9440 8128 9456 8192
rect 9520 8128 9528 8192
rect 9208 8127 9528 8128
rect 39208 8192 39528 8193
rect 39208 8128 39216 8192
rect 39280 8128 39296 8192
rect 39360 8128 39376 8192
rect 39440 8128 39456 8192
rect 39520 8128 39528 8192
rect 39208 8127 39528 8128
rect 49208 8192 49528 8193
rect 49208 8128 49216 8192
rect 49280 8128 49296 8192
rect 49360 8128 49376 8192
rect 49440 8128 49456 8192
rect 49520 8128 49528 8192
rect 49208 8127 49528 8128
rect 59208 8192 59528 8193
rect 59208 8128 59216 8192
rect 59280 8128 59296 8192
rect 59360 8128 59376 8192
rect 59440 8128 59456 8192
rect 59520 8128 59528 8192
rect 59208 8127 59528 8128
rect 29208 8083 29528 8111
rect 29208 8019 29216 8083
rect 29280 8019 29296 8083
rect 29360 8019 29376 8083
rect 29440 8019 29456 8083
rect 29520 8019 29528 8083
rect 29208 8003 29528 8019
rect 29208 7939 29216 8003
rect 29280 7939 29296 8003
rect 29360 7939 29376 8003
rect 29440 7939 29456 8003
rect 29520 7939 29528 8003
rect 29208 7923 29528 7939
rect 29208 7859 29216 7923
rect 29280 7859 29296 7923
rect 29360 7859 29376 7923
rect 29440 7859 29456 7923
rect 29520 7859 29528 7923
rect 29208 7843 29528 7859
rect 46841 7852 46907 7853
rect 29208 7779 29216 7843
rect 29280 7779 29296 7843
rect 29360 7779 29376 7843
rect 29440 7779 29456 7843
rect 29520 7779 29528 7843
rect 46790 7788 46796 7852
rect 46860 7850 46907 7852
rect 46860 7848 46952 7850
rect 46902 7792 46952 7848
rect 46860 7790 46952 7792
rect 46860 7788 46907 7790
rect 46841 7787 46907 7788
rect 29208 7751 29528 7779
rect 13629 7716 13695 7717
rect 13629 7714 13676 7716
rect 13584 7712 13676 7714
rect 13584 7656 13634 7712
rect 13584 7654 13676 7656
rect 13629 7652 13676 7654
rect 13740 7652 13746 7716
rect 13629 7651 13695 7652
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 14208 7648 14528 7649
rect 14208 7584 14216 7648
rect 14280 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14528 7648
rect 14208 7583 14528 7584
rect 44208 7648 44528 7649
rect 44208 7584 44216 7648
rect 44280 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44528 7648
rect 44208 7583 44528 7584
rect 54208 7648 54528 7649
rect 54208 7584 54216 7648
rect 54280 7584 54296 7648
rect 54360 7584 54376 7648
rect 54440 7584 54456 7648
rect 54520 7584 54528 7648
rect 54208 7583 54528 7584
rect 64208 7648 64528 7649
rect 64208 7584 64216 7648
rect 64280 7584 64296 7648
rect 64360 7584 64376 7648
rect 64440 7584 64456 7648
rect 64520 7584 64528 7648
rect 64208 7583 64528 7584
rect 11421 7442 11487 7445
rect 38745 7442 38811 7445
rect 38878 7442 38884 7444
rect 11421 7440 11530 7442
rect 11421 7384 11426 7440
rect 11482 7384 11530 7440
rect 11421 7379 11530 7384
rect 38745 7440 38884 7442
rect 38745 7384 38750 7440
rect 38806 7384 38884 7440
rect 38745 7382 38884 7384
rect 38745 7379 38811 7382
rect 38878 7380 38884 7382
rect 38948 7380 38954 7444
rect 5390 7108 5396 7172
rect 5460 7170 5466 7172
rect 5717 7170 5783 7173
rect 5460 7168 5783 7170
rect 5460 7112 5722 7168
rect 5778 7112 5783 7168
rect 5460 7110 5783 7112
rect 5460 7108 5466 7110
rect 5717 7107 5783 7110
rect 9208 7104 9528 7105
rect 0 7034 800 7064
rect 9208 7040 9216 7104
rect 9280 7040 9296 7104
rect 9360 7040 9376 7104
rect 9440 7040 9456 7104
rect 9520 7040 9528 7104
rect 9208 7039 9528 7040
rect 1577 7034 1643 7037
rect 0 7032 1643 7034
rect 0 6976 1582 7032
rect 1638 6976 1643 7032
rect 0 6974 1643 6976
rect 0 6944 800 6974
rect 1577 6971 1643 6974
rect 11470 6898 11530 7379
rect 68093 7170 68159 7173
rect 69200 7170 70000 7200
rect 68093 7168 70000 7170
rect 68093 7112 68098 7168
rect 68154 7112 70000 7168
rect 68093 7110 70000 7112
rect 68093 7107 68159 7110
rect 39208 7104 39528 7105
rect 39208 7040 39216 7104
rect 39280 7040 39296 7104
rect 39360 7040 39376 7104
rect 39440 7040 39456 7104
rect 39520 7040 39528 7104
rect 39208 7039 39528 7040
rect 49208 7104 49528 7105
rect 49208 7040 49216 7104
rect 49280 7040 49296 7104
rect 49360 7040 49376 7104
rect 49440 7040 49456 7104
rect 49520 7040 49528 7104
rect 49208 7039 49528 7040
rect 59208 7104 59528 7105
rect 59208 7040 59216 7104
rect 59280 7040 59296 7104
rect 59360 7040 59376 7104
rect 59440 7040 59456 7104
rect 59520 7040 59528 7104
rect 69200 7080 70000 7110
rect 59208 7039 59528 7040
rect 15837 7034 15903 7037
rect 39665 7036 39731 7037
rect 15837 7032 16130 7034
rect 15837 6976 15842 7032
rect 15898 6976 16130 7032
rect 15837 6974 16130 6976
rect 15837 6971 15903 6974
rect 12157 6898 12223 6901
rect 11470 6896 12223 6898
rect 11470 6840 12162 6896
rect 12218 6840 12223 6896
rect 11470 6838 12223 6840
rect 12157 6835 12223 6838
rect 16070 6765 16130 6974
rect 39614 6972 39620 7036
rect 39684 7034 39731 7036
rect 39684 7032 39776 7034
rect 39726 6976 39776 7032
rect 39684 6974 39776 6976
rect 39684 6972 39731 6974
rect 39665 6971 39731 6972
rect 35157 6898 35223 6901
rect 42885 6898 42951 6901
rect 35157 6896 42951 6898
rect 35157 6840 35162 6896
rect 35218 6840 42890 6896
rect 42946 6840 42951 6896
rect 35157 6838 42951 6840
rect 24208 6809 24528 6837
rect 16070 6760 16179 6765
rect 16070 6704 16118 6760
rect 16174 6704 16179 6760
rect 16070 6702 16179 6704
rect 16113 6699 16179 6702
rect 24208 6745 24216 6809
rect 24280 6745 24296 6809
rect 24360 6745 24376 6809
rect 24440 6745 24456 6809
rect 24520 6745 24528 6809
rect 24208 6729 24528 6745
rect 24208 6665 24216 6729
rect 24280 6665 24296 6729
rect 24360 6665 24376 6729
rect 24440 6665 24456 6729
rect 24520 6665 24528 6729
rect 24208 6649 24528 6665
rect 24208 6585 24216 6649
rect 24280 6585 24296 6649
rect 24360 6585 24376 6649
rect 24440 6585 24456 6649
rect 24520 6585 24528 6649
rect 24208 6569 24528 6585
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 14208 6560 14528 6561
rect 14208 6496 14216 6560
rect 14280 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14528 6560
rect 14208 6495 14528 6496
rect 24208 6505 24216 6569
rect 24280 6505 24296 6569
rect 24360 6505 24376 6569
rect 24440 6505 24456 6569
rect 24520 6505 24528 6569
rect 24208 6477 24528 6505
rect 34208 6809 34528 6837
rect 35157 6835 35223 6838
rect 42885 6835 42951 6838
rect 65241 6898 65307 6901
rect 65793 6898 65859 6901
rect 65241 6896 65859 6898
rect 65241 6840 65246 6896
rect 65302 6840 65798 6896
rect 65854 6840 65859 6896
rect 65241 6838 65859 6840
rect 65241 6835 65307 6838
rect 65793 6835 65859 6838
rect 34208 6745 34216 6809
rect 34280 6745 34296 6809
rect 34360 6745 34376 6809
rect 34440 6745 34456 6809
rect 34520 6745 34528 6809
rect 34208 6729 34528 6745
rect 34208 6665 34216 6729
rect 34280 6665 34296 6729
rect 34360 6665 34376 6729
rect 34440 6665 34456 6729
rect 34520 6665 34528 6729
rect 34208 6649 34528 6665
rect 34208 6585 34216 6649
rect 34280 6585 34296 6649
rect 34360 6585 34376 6649
rect 34440 6585 34456 6649
rect 34520 6585 34528 6649
rect 34208 6569 34528 6585
rect 34208 6505 34216 6569
rect 34280 6505 34296 6569
rect 34360 6505 34376 6569
rect 34440 6505 34456 6569
rect 34520 6505 34528 6569
rect 39849 6626 39915 6629
rect 40401 6626 40467 6629
rect 39849 6624 40467 6626
rect 39849 6568 39854 6624
rect 39910 6568 40406 6624
rect 40462 6568 40467 6624
rect 39849 6566 40467 6568
rect 39849 6563 39915 6566
rect 40401 6563 40467 6566
rect 34208 6477 34528 6505
rect 44208 6560 44528 6561
rect 44208 6496 44216 6560
rect 44280 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44528 6560
rect 44208 6495 44528 6496
rect 54208 6560 54528 6561
rect 54208 6496 54216 6560
rect 54280 6496 54296 6560
rect 54360 6496 54376 6560
rect 54440 6496 54456 6560
rect 54520 6496 54528 6560
rect 54208 6495 54528 6496
rect 64208 6560 64528 6561
rect 64208 6496 64216 6560
rect 64280 6496 64296 6560
rect 64360 6496 64376 6560
rect 64440 6496 64456 6560
rect 64520 6496 64528 6560
rect 64208 6495 64528 6496
rect 36721 6490 36787 6493
rect 41689 6490 41755 6493
rect 36721 6488 41755 6490
rect 36721 6432 36726 6488
rect 36782 6432 41694 6488
rect 41750 6432 41755 6488
rect 36721 6430 41755 6432
rect 36721 6427 36787 6430
rect 41689 6427 41755 6430
rect 14457 6354 14523 6357
rect 14590 6354 14596 6356
rect 14457 6352 14596 6354
rect 14457 6296 14462 6352
rect 14518 6296 14596 6352
rect 14457 6294 14596 6296
rect 14457 6291 14523 6294
rect 14590 6292 14596 6294
rect 14660 6292 14666 6356
rect 18781 6354 18847 6357
rect 37917 6354 37983 6357
rect 18781 6352 37983 6354
rect 18781 6296 18786 6352
rect 18842 6296 37922 6352
rect 37978 6296 37983 6352
rect 18781 6294 37983 6296
rect 18781 6291 18847 6294
rect 37917 6291 37983 6294
rect 23933 6218 23999 6221
rect 65241 6218 65307 6221
rect 23933 6216 65307 6218
rect 23933 6160 23938 6216
rect 23994 6160 65246 6216
rect 65302 6160 65307 6216
rect 23933 6158 65307 6160
rect 23933 6155 23999 6158
rect 65241 6155 65307 6158
rect 15285 6082 15351 6085
rect 15469 6082 15535 6085
rect 23933 6082 23999 6085
rect 15285 6080 23999 6082
rect 15285 6024 15290 6080
rect 15346 6024 15474 6080
rect 15530 6024 23938 6080
rect 23994 6024 23999 6080
rect 15285 6022 23999 6024
rect 15285 6019 15351 6022
rect 15469 6019 15535 6022
rect 23933 6019 23999 6022
rect 30414 6020 30420 6084
rect 30484 6082 30490 6084
rect 38653 6082 38719 6085
rect 30484 6080 38719 6082
rect 30484 6024 38658 6080
rect 38714 6024 38719 6080
rect 30484 6022 38719 6024
rect 30484 6020 30490 6022
rect 38653 6019 38719 6022
rect 40493 6082 40559 6085
rect 41137 6082 41203 6085
rect 40493 6080 41203 6082
rect 40493 6024 40498 6080
rect 40554 6024 41142 6080
rect 41198 6024 41203 6080
rect 40493 6022 41203 6024
rect 40493 6019 40559 6022
rect 41137 6019 41203 6022
rect 42006 6020 42012 6084
rect 42076 6082 42082 6084
rect 43069 6082 43135 6085
rect 42076 6080 43135 6082
rect 42076 6024 43074 6080
rect 43130 6024 43135 6080
rect 42076 6022 43135 6024
rect 42076 6020 42082 6022
rect 43069 6019 43135 6022
rect 9208 6016 9528 6017
rect 9208 5952 9216 6016
rect 9280 5952 9296 6016
rect 9360 5952 9376 6016
rect 9440 5952 9456 6016
rect 9520 5952 9528 6016
rect 9208 5951 9528 5952
rect 39208 6016 39528 6017
rect 39208 5952 39216 6016
rect 39280 5952 39296 6016
rect 39360 5952 39376 6016
rect 39440 5952 39456 6016
rect 39520 5952 39528 6016
rect 39208 5951 39528 5952
rect 49208 6016 49528 6017
rect 49208 5952 49216 6016
rect 49280 5952 49296 6016
rect 49360 5952 49376 6016
rect 49440 5952 49456 6016
rect 49520 5952 49528 6016
rect 49208 5951 49528 5952
rect 59208 6016 59528 6017
rect 59208 5952 59216 6016
rect 59280 5952 59296 6016
rect 59360 5952 59376 6016
rect 59440 5952 59456 6016
rect 59520 5952 59528 6016
rect 59208 5951 59528 5952
rect 13169 5946 13235 5949
rect 23473 5946 23539 5949
rect 13169 5944 23539 5946
rect 13169 5888 13174 5944
rect 13230 5888 23478 5944
rect 23534 5888 23539 5944
rect 13169 5886 23539 5888
rect 13169 5883 13235 5886
rect 23473 5883 23539 5886
rect 27654 5884 27660 5948
rect 27724 5946 27730 5948
rect 38561 5946 38627 5949
rect 42333 5946 42399 5949
rect 27724 5944 38627 5946
rect 27724 5888 38566 5944
rect 38622 5888 38627 5944
rect 27724 5886 38627 5888
rect 27724 5884 27730 5886
rect 38561 5883 38627 5886
rect 39622 5944 42399 5946
rect 39622 5888 42338 5944
rect 42394 5888 42399 5944
rect 39622 5886 42399 5888
rect 0 5810 800 5840
rect 1761 5810 1827 5813
rect 0 5808 1827 5810
rect 0 5752 1766 5808
rect 1822 5752 1827 5808
rect 0 5750 1827 5752
rect 0 5720 800 5750
rect 1761 5747 1827 5750
rect 13629 5810 13695 5813
rect 18873 5810 18939 5813
rect 13629 5808 18939 5810
rect 13629 5752 13634 5808
rect 13690 5752 18878 5808
rect 18934 5752 18939 5808
rect 13629 5750 18939 5752
rect 13629 5747 13695 5750
rect 18873 5747 18939 5750
rect 33133 5810 33199 5813
rect 39622 5810 39682 5886
rect 42333 5883 42399 5886
rect 46657 5812 46723 5813
rect 33133 5808 39682 5810
rect 33133 5752 33138 5808
rect 33194 5752 39682 5808
rect 33133 5750 39682 5752
rect 33133 5747 33199 5750
rect 46606 5748 46612 5812
rect 46676 5810 46723 5812
rect 68093 5810 68159 5813
rect 69200 5810 70000 5840
rect 46676 5808 46768 5810
rect 46718 5752 46768 5808
rect 46676 5750 46768 5752
rect 68093 5808 70000 5810
rect 68093 5752 68098 5808
rect 68154 5752 70000 5808
rect 68093 5750 70000 5752
rect 46676 5748 46723 5750
rect 46657 5747 46723 5748
rect 68093 5747 68159 5750
rect 69200 5720 70000 5750
rect 16573 5674 16639 5677
rect 21173 5674 21239 5677
rect 16573 5672 21239 5674
rect 16573 5616 16578 5672
rect 16634 5616 21178 5672
rect 21234 5616 21239 5672
rect 16573 5614 21239 5616
rect 16573 5611 16639 5614
rect 21173 5611 21239 5614
rect 39205 5674 39271 5677
rect 59537 5674 59603 5677
rect 60641 5674 60707 5677
rect 39205 5672 60707 5674
rect 39205 5616 39210 5672
rect 39266 5616 59542 5672
rect 59598 5616 60646 5672
rect 60702 5616 60707 5672
rect 39205 5614 60707 5616
rect 39205 5611 39271 5614
rect 59537 5611 59603 5614
rect 60641 5611 60707 5614
rect 30598 5476 30604 5540
rect 30668 5538 30674 5540
rect 40033 5538 40099 5541
rect 30668 5536 40099 5538
rect 30668 5480 40038 5536
rect 40094 5480 40099 5536
rect 30668 5478 40099 5480
rect 30668 5476 30674 5478
rect 40033 5475 40099 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 14208 5472 14528 5473
rect 14208 5408 14216 5472
rect 14280 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14528 5472
rect 14208 5407 14528 5408
rect 44208 5472 44528 5473
rect 44208 5408 44216 5472
rect 44280 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44528 5472
rect 44208 5407 44528 5408
rect 54208 5472 54528 5473
rect 54208 5408 54216 5472
rect 54280 5408 54296 5472
rect 54360 5408 54376 5472
rect 54440 5408 54456 5472
rect 54520 5408 54528 5472
rect 54208 5407 54528 5408
rect 64208 5472 64528 5473
rect 64208 5408 64216 5472
rect 64280 5408 64296 5472
rect 64360 5408 64376 5472
rect 64440 5408 64456 5472
rect 64520 5408 64528 5472
rect 64208 5407 64528 5408
rect 31886 5340 31892 5404
rect 31956 5402 31962 5404
rect 43345 5402 43411 5405
rect 31956 5400 43411 5402
rect 31956 5344 43350 5400
rect 43406 5344 43411 5400
rect 31956 5342 43411 5344
rect 31956 5340 31962 5342
rect 43345 5339 43411 5342
rect 3969 5266 4035 5269
rect 17217 5266 17283 5269
rect 3969 5264 17283 5266
rect 3969 5208 3974 5264
rect 4030 5208 17222 5264
rect 17278 5208 17283 5264
rect 3969 5206 17283 5208
rect 3969 5203 4035 5206
rect 17217 5203 17283 5206
rect 30046 5204 30052 5268
rect 30116 5266 30122 5268
rect 41781 5266 41847 5269
rect 55949 5268 56015 5269
rect 55949 5266 55996 5268
rect 30116 5264 41847 5266
rect 30116 5208 41786 5264
rect 41842 5208 41847 5264
rect 30116 5206 41847 5208
rect 55904 5264 55996 5266
rect 55904 5208 55954 5264
rect 55904 5206 55996 5208
rect 30116 5204 30122 5206
rect 41781 5203 41847 5206
rect 55949 5204 55996 5206
rect 56060 5204 56066 5268
rect 55949 5203 56015 5204
rect 5441 5132 5507 5133
rect 5390 5068 5396 5132
rect 5460 5130 5507 5132
rect 33041 5130 33107 5133
rect 68277 5130 68343 5133
rect 5460 5128 5552 5130
rect 5502 5072 5552 5128
rect 5460 5070 5552 5072
rect 33041 5128 68343 5130
rect 33041 5072 33046 5128
rect 33102 5072 68282 5128
rect 68338 5072 68343 5128
rect 33041 5070 68343 5072
rect 5460 5068 5507 5070
rect 5441 5067 5507 5068
rect 33041 5067 33107 5070
rect 68277 5067 68343 5070
rect 53598 4932 53604 4996
rect 53668 4994 53674 4996
rect 53741 4994 53807 4997
rect 54937 4996 55003 4997
rect 53668 4992 53807 4994
rect 53668 4936 53746 4992
rect 53802 4936 53807 4992
rect 53668 4934 53807 4936
rect 53668 4932 53674 4934
rect 53741 4931 53807 4934
rect 54886 4932 54892 4996
rect 54956 4994 55003 4996
rect 54956 4992 55048 4994
rect 54998 4936 55048 4992
rect 54956 4934 55048 4936
rect 54956 4932 55003 4934
rect 54937 4931 55003 4932
rect 9208 4928 9528 4929
rect 9208 4864 9216 4928
rect 9280 4864 9296 4928
rect 9360 4864 9376 4928
rect 9440 4864 9456 4928
rect 9520 4864 9528 4928
rect 9208 4863 9528 4864
rect 39208 4928 39528 4929
rect 39208 4864 39216 4928
rect 39280 4864 39296 4928
rect 39360 4864 39376 4928
rect 39440 4864 39456 4928
rect 39520 4864 39528 4928
rect 39208 4863 39528 4864
rect 49208 4928 49528 4929
rect 49208 4864 49216 4928
rect 49280 4864 49296 4928
rect 49360 4864 49376 4928
rect 49440 4864 49456 4928
rect 49520 4864 49528 4928
rect 49208 4863 49528 4864
rect 59208 4928 59528 4929
rect 59208 4864 59216 4928
rect 59280 4864 59296 4928
rect 59360 4864 59376 4928
rect 59440 4864 59456 4928
rect 59520 4864 59528 4928
rect 59208 4863 59528 4864
rect 16205 4858 16271 4861
rect 24117 4858 24183 4861
rect 16205 4856 24183 4858
rect 16205 4800 16210 4856
rect 16266 4800 24122 4856
rect 24178 4800 24183 4856
rect 16205 4798 24183 4800
rect 16205 4795 16271 4798
rect 24117 4795 24183 4798
rect 31150 4660 31156 4724
rect 31220 4722 31226 4724
rect 39021 4722 39087 4725
rect 31220 4720 39087 4722
rect 31220 4664 39026 4720
rect 39082 4664 39087 4720
rect 31220 4662 39087 4664
rect 31220 4660 31226 4662
rect 39021 4659 39087 4662
rect 39849 4722 39915 4725
rect 40902 4722 40908 4724
rect 39849 4720 40908 4722
rect 39849 4664 39854 4720
rect 39910 4664 40908 4720
rect 39849 4662 40908 4664
rect 39849 4659 39915 4662
rect 40902 4660 40908 4662
rect 40972 4660 40978 4724
rect 42609 4722 42675 4725
rect 43621 4722 43687 4725
rect 42609 4720 43687 4722
rect 42609 4664 42614 4720
rect 42670 4664 43626 4720
rect 43682 4664 43687 4720
rect 42609 4662 43687 4664
rect 42609 4659 42675 4662
rect 43621 4659 43687 4662
rect 39665 4586 39731 4589
rect 39982 4586 39988 4588
rect 39665 4584 39988 4586
rect 39665 4528 39670 4584
rect 39726 4528 39988 4584
rect 39665 4526 39988 4528
rect 39665 4523 39731 4526
rect 39982 4524 39988 4526
rect 40052 4524 40058 4588
rect 41137 4586 41203 4589
rect 44173 4586 44239 4589
rect 64689 4588 64755 4589
rect 41137 4584 44239 4586
rect 41137 4528 41142 4584
rect 41198 4528 44178 4584
rect 44234 4528 44239 4584
rect 41137 4526 44239 4528
rect 41137 4523 41203 4526
rect 44173 4523 44239 4526
rect 64638 4524 64644 4588
rect 64708 4586 64755 4588
rect 67541 4586 67607 4589
rect 69200 4586 70000 4616
rect 64708 4584 64800 4586
rect 64750 4528 64800 4584
rect 64708 4526 64800 4528
rect 67541 4584 70000 4586
rect 67541 4528 67546 4584
rect 67602 4528 70000 4584
rect 67541 4526 70000 4528
rect 64708 4524 64755 4526
rect 64689 4523 64755 4524
rect 67541 4523 67607 4526
rect 69200 4496 70000 4526
rect 0 4450 800 4480
rect 1853 4450 1919 4453
rect 0 4448 1919 4450
rect 0 4392 1858 4448
rect 1914 4392 1919 4448
rect 0 4390 1919 4392
rect 0 4360 800 4390
rect 1853 4387 1919 4390
rect 38878 4388 38884 4452
rect 38948 4450 38954 4452
rect 43345 4450 43411 4453
rect 38948 4448 43411 4450
rect 38948 4392 43350 4448
rect 43406 4392 43411 4448
rect 38948 4390 43411 4392
rect 38948 4388 38954 4390
rect 43345 4387 43411 4390
rect 46197 4450 46263 4453
rect 48497 4450 48563 4453
rect 46197 4448 48563 4450
rect 46197 4392 46202 4448
rect 46258 4392 48502 4448
rect 48558 4392 48563 4448
rect 46197 4390 48563 4392
rect 46197 4387 46263 4390
rect 48497 4387 48563 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 14208 4384 14528 4385
rect 14208 4320 14216 4384
rect 14280 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14528 4384
rect 14208 4319 14528 4320
rect 44208 4384 44528 4385
rect 44208 4320 44216 4384
rect 44280 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44528 4384
rect 44208 4319 44528 4320
rect 54208 4384 54528 4385
rect 54208 4320 54216 4384
rect 54280 4320 54296 4384
rect 54360 4320 54376 4384
rect 54440 4320 54456 4384
rect 54520 4320 54528 4384
rect 54208 4319 54528 4320
rect 64208 4384 64528 4385
rect 64208 4320 64216 4384
rect 64280 4320 64296 4384
rect 64360 4320 64376 4384
rect 64440 4320 64456 4384
rect 64520 4320 64528 4384
rect 64208 4319 64528 4320
rect 6821 4178 6887 4181
rect 16481 4178 16547 4181
rect 6821 4176 16547 4178
rect 6821 4120 6826 4176
rect 6882 4120 16486 4176
rect 16542 4120 16547 4176
rect 6821 4118 16547 4120
rect 6821 4115 6887 4118
rect 16481 4115 16547 4118
rect 38653 4178 38719 4181
rect 39389 4178 39455 4181
rect 38653 4176 39455 4178
rect 38653 4120 38658 4176
rect 38714 4120 39394 4176
rect 39450 4120 39455 4176
rect 38653 4118 39455 4120
rect 38653 4115 38719 4118
rect 39389 4115 39455 4118
rect 9213 4042 9279 4045
rect 9078 4040 9279 4042
rect 9078 3984 9218 4040
rect 9274 3984 9279 4040
rect 9078 3982 9279 3984
rect 8937 3906 9003 3909
rect 9078 3906 9138 3982
rect 9213 3979 9279 3982
rect 11646 3980 11652 4044
rect 11716 4042 11722 4044
rect 12249 4042 12315 4045
rect 11716 4040 12315 4042
rect 11716 3984 12254 4040
rect 12310 3984 12315 4040
rect 11716 3982 12315 3984
rect 11716 3980 11722 3982
rect 12249 3979 12315 3982
rect 13670 3980 13676 4044
rect 13740 4042 13746 4044
rect 14457 4042 14523 4045
rect 13740 4040 14523 4042
rect 13740 3984 14462 4040
rect 14518 3984 14523 4040
rect 13740 3982 14523 3984
rect 13740 3980 13746 3982
rect 14457 3979 14523 3982
rect 16205 4044 16271 4045
rect 16205 4040 16252 4044
rect 16316 4042 16322 4044
rect 43253 4042 43319 4045
rect 16205 3984 16210 4040
rect 16205 3980 16252 3984
rect 16316 3982 16362 4042
rect 31710 4040 43319 4042
rect 31710 3984 43258 4040
rect 43314 3984 43319 4040
rect 31710 3982 43319 3984
rect 16316 3980 16322 3982
rect 16205 3979 16271 3980
rect 8937 3904 9138 3906
rect 8937 3848 8942 3904
rect 8998 3848 9138 3904
rect 8937 3846 9138 3848
rect 11053 3906 11119 3909
rect 13537 3906 13603 3909
rect 11053 3904 13603 3906
rect 11053 3848 11058 3904
rect 11114 3848 13542 3904
rect 13598 3848 13603 3904
rect 11053 3846 13603 3848
rect 8937 3843 9003 3846
rect 11053 3843 11119 3846
rect 13537 3843 13603 3846
rect 13997 3908 14063 3909
rect 13997 3904 14044 3908
rect 14108 3906 14114 3908
rect 14365 3906 14431 3909
rect 21633 3906 21699 3909
rect 31710 3906 31770 3982
rect 43253 3979 43319 3982
rect 49734 3980 49740 4044
rect 49804 4042 49810 4044
rect 49877 4042 49943 4045
rect 49804 4040 49943 4042
rect 49804 3984 49882 4040
rect 49938 3984 49943 4040
rect 49804 3982 49943 3984
rect 49804 3980 49810 3982
rect 49877 3979 49943 3982
rect 13997 3848 14002 3904
rect 13997 3844 14044 3848
rect 14108 3846 14154 3906
rect 14365 3904 21699 3906
rect 14365 3848 14370 3904
rect 14426 3848 21638 3904
rect 21694 3848 21699 3904
rect 14365 3846 21699 3848
rect 14108 3844 14114 3846
rect 13997 3843 14063 3844
rect 14365 3843 14431 3846
rect 21633 3843 21699 3846
rect 26926 3846 31770 3906
rect 32397 3906 32463 3909
rect 38878 3906 38884 3908
rect 32397 3904 38884 3906
rect 32397 3848 32402 3904
rect 32458 3848 38884 3904
rect 32397 3846 38884 3848
rect 9208 3840 9528 3841
rect 9208 3776 9216 3840
rect 9280 3776 9296 3840
rect 9360 3776 9376 3840
rect 9440 3776 9456 3840
rect 9520 3776 9528 3840
rect 9208 3775 9528 3776
rect 9622 3708 9628 3772
rect 9692 3770 9698 3772
rect 9765 3770 9831 3773
rect 9692 3768 9831 3770
rect 9692 3712 9770 3768
rect 9826 3712 9831 3768
rect 9692 3710 9831 3712
rect 9692 3708 9698 3710
rect 9765 3707 9831 3710
rect 11513 3770 11579 3773
rect 12065 3770 12131 3773
rect 11513 3768 11852 3770
rect 11513 3712 11518 3768
rect 11574 3712 11852 3768
rect 11513 3710 11852 3712
rect 11513 3707 11579 3710
rect 10041 3634 10107 3637
rect 10501 3634 10567 3637
rect 10041 3632 10567 3634
rect 10041 3576 10046 3632
rect 10102 3576 10506 3632
rect 10562 3576 10567 3632
rect 10041 3574 10567 3576
rect 10041 3571 10107 3574
rect 10501 3571 10567 3574
rect 9857 3498 9923 3501
rect 9814 3496 9923 3498
rect 9814 3440 9862 3496
rect 9918 3440 9923 3496
rect 9814 3435 9923 3440
rect 11792 3498 11852 3710
rect 12022 3768 12131 3770
rect 12022 3712 12070 3768
rect 12126 3712 12131 3768
rect 12022 3707 12131 3712
rect 12198 3708 12204 3772
rect 12268 3770 12274 3772
rect 12433 3770 12499 3773
rect 12268 3768 12499 3770
rect 12268 3712 12438 3768
rect 12494 3712 12499 3768
rect 12268 3710 12499 3712
rect 12268 3708 12274 3710
rect 12433 3707 12499 3710
rect 13353 3770 13419 3773
rect 13486 3770 13492 3772
rect 13353 3768 13492 3770
rect 13353 3712 13358 3768
rect 13414 3712 13492 3768
rect 13353 3710 13492 3712
rect 13353 3707 13419 3710
rect 13486 3708 13492 3710
rect 13556 3708 13562 3772
rect 15469 3770 15535 3773
rect 22645 3770 22711 3773
rect 15469 3768 22711 3770
rect 15469 3712 15474 3768
rect 15530 3712 22650 3768
rect 22706 3712 22711 3768
rect 15469 3710 22711 3712
rect 15469 3707 15535 3710
rect 22645 3707 22711 3710
rect 12022 3634 12082 3707
rect 16573 3634 16639 3637
rect 12022 3632 16639 3634
rect 12022 3576 16578 3632
rect 16634 3576 16639 3632
rect 12022 3574 16639 3576
rect 16573 3571 16639 3574
rect 17493 3498 17559 3501
rect 26926 3498 26986 3846
rect 32397 3843 32463 3846
rect 38878 3844 38884 3846
rect 38948 3844 38954 3908
rect 46565 3906 46631 3909
rect 47853 3906 47919 3909
rect 46565 3904 47919 3906
rect 46565 3848 46570 3904
rect 46626 3848 47858 3904
rect 47914 3848 47919 3904
rect 46565 3846 47919 3848
rect 46565 3843 46631 3846
rect 47853 3843 47919 3846
rect 49877 3906 49943 3909
rect 50705 3906 50771 3909
rect 49877 3904 50771 3906
rect 49877 3848 49882 3904
rect 49938 3848 50710 3904
rect 50766 3848 50771 3904
rect 49877 3846 50771 3848
rect 49877 3843 49943 3846
rect 50705 3843 50771 3846
rect 65149 3906 65215 3909
rect 65149 3904 65258 3906
rect 65149 3848 65154 3904
rect 65210 3848 65258 3904
rect 65149 3843 65258 3848
rect 39208 3840 39528 3841
rect 39208 3776 39216 3840
rect 39280 3776 39296 3840
rect 39360 3776 39376 3840
rect 39440 3776 39456 3840
rect 39520 3776 39528 3840
rect 39208 3775 39528 3776
rect 49208 3840 49528 3841
rect 49208 3776 49216 3840
rect 49280 3776 49296 3840
rect 49360 3776 49376 3840
rect 49440 3776 49456 3840
rect 49520 3776 49528 3840
rect 49208 3775 49528 3776
rect 59208 3840 59528 3841
rect 59208 3776 59216 3840
rect 59280 3776 59296 3840
rect 59360 3776 59376 3840
rect 59440 3776 59456 3840
rect 59520 3776 59528 3840
rect 59208 3775 59528 3776
rect 28206 3708 28212 3772
rect 28276 3770 28282 3772
rect 33726 3770 33732 3772
rect 28276 3710 33732 3770
rect 28276 3708 28282 3710
rect 33726 3708 33732 3710
rect 33796 3708 33802 3772
rect 33961 3770 34027 3773
rect 35985 3770 36051 3773
rect 39021 3770 39087 3773
rect 33961 3768 36051 3770
rect 33961 3712 33966 3768
rect 34022 3712 35990 3768
rect 36046 3712 36051 3768
rect 33961 3710 36051 3712
rect 33961 3707 34027 3710
rect 35985 3707 36051 3710
rect 38518 3768 39087 3770
rect 38518 3712 39026 3768
rect 39082 3712 39087 3768
rect 38518 3710 39087 3712
rect 28022 3572 28028 3636
rect 28092 3634 28098 3636
rect 32765 3634 32831 3637
rect 28092 3632 32831 3634
rect 28092 3576 32770 3632
rect 32826 3576 32831 3632
rect 28092 3574 32831 3576
rect 28092 3572 28098 3574
rect 32765 3571 32831 3574
rect 33041 3634 33107 3637
rect 38518 3634 38578 3710
rect 39021 3707 39087 3710
rect 43713 3770 43779 3773
rect 55949 3772 56015 3773
rect 44030 3770 44036 3772
rect 43713 3768 44036 3770
rect 43713 3712 43718 3768
rect 43774 3712 44036 3768
rect 43713 3710 44036 3712
rect 43713 3707 43779 3710
rect 44030 3708 44036 3710
rect 44100 3708 44106 3772
rect 55949 3768 55996 3772
rect 56060 3770 56066 3772
rect 55949 3712 55954 3768
rect 55949 3708 55996 3712
rect 56060 3710 56106 3770
rect 56060 3708 56066 3710
rect 55949 3707 56015 3708
rect 33041 3632 38578 3634
rect 33041 3576 33046 3632
rect 33102 3576 38578 3632
rect 33041 3574 38578 3576
rect 38653 3634 38719 3637
rect 44541 3634 44607 3637
rect 45645 3634 45711 3637
rect 38653 3632 45711 3634
rect 38653 3576 38658 3632
rect 38714 3576 44546 3632
rect 44602 3576 45650 3632
rect 45706 3576 45711 3632
rect 38653 3574 45711 3576
rect 33041 3571 33107 3574
rect 38653 3571 38719 3574
rect 44541 3571 44607 3574
rect 45645 3571 45711 3574
rect 11792 3438 14658 3498
rect 4208 3296 4528 3297
rect 0 3226 800 3256
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 1577 3226 1643 3229
rect 0 3224 1643 3226
rect 0 3168 1582 3224
rect 1638 3168 1643 3224
rect 0 3166 1643 3168
rect 0 3136 800 3166
rect 1577 3163 1643 3166
rect 9814 2821 9874 3435
rect 14598 3362 14658 3438
rect 17493 3496 26986 3498
rect 17493 3440 17498 3496
rect 17554 3440 26986 3496
rect 17493 3438 26986 3440
rect 31845 3498 31911 3501
rect 39757 3498 39823 3501
rect 31845 3496 39823 3498
rect 31845 3440 31850 3496
rect 31906 3440 39762 3496
rect 39818 3440 39823 3496
rect 31845 3438 39823 3440
rect 17493 3435 17559 3438
rect 31845 3435 31911 3438
rect 39757 3435 39823 3438
rect 45093 3498 45159 3501
rect 48405 3498 48471 3501
rect 45093 3496 48471 3498
rect 45093 3440 45098 3496
rect 45154 3440 48410 3496
rect 48466 3440 48471 3496
rect 45093 3438 48471 3440
rect 65198 3498 65258 3843
rect 67449 3634 67515 3637
rect 67406 3632 67515 3634
rect 67406 3576 67454 3632
rect 67510 3576 67515 3632
rect 67406 3571 67515 3576
rect 65517 3498 65583 3501
rect 65198 3496 65583 3498
rect 65198 3440 65522 3496
rect 65578 3440 65583 3496
rect 65198 3438 65583 3440
rect 45093 3435 45159 3438
rect 48405 3435 48471 3438
rect 65517 3435 65583 3438
rect 19057 3362 19123 3365
rect 14598 3360 19123 3362
rect 14598 3304 19062 3360
rect 19118 3304 19123 3360
rect 14598 3302 19123 3304
rect 19057 3299 19123 3302
rect 33869 3362 33935 3365
rect 38653 3362 38719 3365
rect 33869 3360 38719 3362
rect 33869 3304 33874 3360
rect 33930 3304 38658 3360
rect 38714 3304 38719 3360
rect 33869 3302 38719 3304
rect 33869 3299 33935 3302
rect 38653 3299 38719 3302
rect 39062 3300 39068 3364
rect 39132 3362 39138 3364
rect 39205 3362 39271 3365
rect 39132 3360 39271 3362
rect 39132 3304 39210 3360
rect 39266 3304 39271 3360
rect 39132 3302 39271 3304
rect 39132 3300 39138 3302
rect 39205 3299 39271 3302
rect 39481 3362 39547 3365
rect 39798 3362 39804 3364
rect 39481 3360 39804 3362
rect 39481 3304 39486 3360
rect 39542 3304 39804 3360
rect 39481 3302 39804 3304
rect 39481 3299 39547 3302
rect 39798 3300 39804 3302
rect 39868 3300 39874 3364
rect 41689 3362 41755 3365
rect 42057 3362 42123 3365
rect 41689 3360 42123 3362
rect 41689 3304 41694 3360
rect 41750 3304 42062 3360
rect 42118 3304 42123 3360
rect 41689 3302 42123 3304
rect 41689 3299 41755 3302
rect 42057 3299 42123 3302
rect 45461 3362 45527 3365
rect 46790 3362 46796 3364
rect 45461 3360 46796 3362
rect 45461 3304 45466 3360
rect 45522 3304 46796 3360
rect 45461 3302 46796 3304
rect 45461 3299 45527 3302
rect 46790 3300 46796 3302
rect 46860 3300 46866 3364
rect 14208 3296 14528 3297
rect 14208 3232 14216 3296
rect 14280 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14528 3296
rect 44208 3296 44528 3297
rect 14208 3231 14528 3232
rect 24208 3222 24528 3260
rect 44208 3232 44216 3296
rect 44280 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44528 3296
rect 44208 3231 44528 3232
rect 54208 3296 54528 3297
rect 54208 3232 54216 3296
rect 54280 3232 54296 3296
rect 54360 3232 54376 3296
rect 54440 3232 54456 3296
rect 54520 3232 54528 3296
rect 54208 3231 54528 3232
rect 64208 3296 64528 3297
rect 64208 3232 64216 3296
rect 64280 3232 64296 3296
rect 64360 3232 64376 3296
rect 64440 3232 64456 3296
rect 64520 3232 64528 3296
rect 64208 3231 64528 3232
rect 67406 3229 67466 3571
rect 24208 3158 24216 3222
rect 24280 3158 24296 3222
rect 24360 3158 24376 3222
rect 24440 3158 24456 3222
rect 24520 3158 24528 3222
rect 34697 3226 34763 3229
rect 42885 3226 42951 3229
rect 34697 3224 42951 3226
rect 34697 3168 34702 3224
rect 34758 3168 42890 3224
rect 42946 3168 42951 3224
rect 34697 3166 42951 3168
rect 34697 3163 34763 3166
rect 42885 3163 42951 3166
rect 47577 3226 47643 3229
rect 50889 3226 50955 3229
rect 51073 3226 51139 3229
rect 47577 3224 47778 3226
rect 47577 3168 47582 3224
rect 47638 3168 47778 3224
rect 47577 3166 47778 3168
rect 47577 3163 47643 3166
rect 24208 3142 24528 3158
rect 15694 3028 15700 3092
rect 15764 3090 15770 3092
rect 15929 3090 15995 3093
rect 15764 3088 15995 3090
rect 15764 3032 15934 3088
rect 15990 3032 15995 3088
rect 15764 3030 15995 3032
rect 15764 3028 15770 3030
rect 15929 3027 15995 3030
rect 24208 3078 24216 3142
rect 24280 3078 24296 3142
rect 24360 3078 24376 3142
rect 24440 3078 24456 3142
rect 24520 3078 24528 3142
rect 24208 3062 24528 3078
rect 24208 2998 24216 3062
rect 24280 2998 24296 3062
rect 24360 2998 24376 3062
rect 24440 2998 24456 3062
rect 24520 2998 24528 3062
rect 35985 3090 36051 3093
rect 40493 3090 40559 3093
rect 40677 3092 40743 3093
rect 41413 3092 41479 3093
rect 40677 3090 40724 3092
rect 35985 3088 40559 3090
rect 35985 3032 35990 3088
rect 36046 3032 40498 3088
rect 40554 3032 40559 3088
rect 35985 3030 40559 3032
rect 40632 3088 40724 3090
rect 40632 3032 40682 3088
rect 40632 3030 40724 3032
rect 35985 3027 36051 3030
rect 40493 3027 40559 3030
rect 40677 3028 40724 3030
rect 40788 3028 40794 3092
rect 41413 3090 41460 3092
rect 41368 3088 41460 3090
rect 41368 3032 41418 3088
rect 41368 3030 41460 3032
rect 41413 3028 41460 3030
rect 41524 3028 41530 3092
rect 42374 3028 42380 3092
rect 42444 3090 42450 3092
rect 42701 3090 42767 3093
rect 42444 3088 42767 3090
rect 42444 3032 42706 3088
rect 42762 3032 42767 3088
rect 42444 3030 42767 3032
rect 42444 3028 42450 3030
rect 40677 3027 40743 3028
rect 41413 3027 41479 3028
rect 42701 3027 42767 3030
rect 43713 3090 43779 3093
rect 43846 3090 43852 3092
rect 43713 3088 43852 3090
rect 43713 3032 43718 3088
rect 43774 3032 43852 3088
rect 43713 3030 43852 3032
rect 43713 3027 43779 3030
rect 43846 3028 43852 3030
rect 43916 3028 43922 3092
rect 24208 2982 24528 2998
rect 13721 2954 13787 2957
rect 18873 2954 18939 2957
rect 19149 2954 19215 2957
rect 13721 2952 14106 2954
rect 13721 2896 13726 2952
rect 13782 2896 14106 2952
rect 13721 2894 14106 2896
rect 13721 2891 13787 2894
rect 5257 2818 5323 2821
rect 5993 2818 6059 2821
rect 5257 2816 6059 2818
rect 5257 2760 5262 2816
rect 5318 2760 5998 2816
rect 6054 2760 6059 2816
rect 5257 2758 6059 2760
rect 5257 2755 5323 2758
rect 5993 2755 6059 2758
rect 9765 2816 9874 2821
rect 9765 2760 9770 2816
rect 9826 2760 9874 2816
rect 9765 2758 9874 2760
rect 9765 2755 9831 2758
rect 9208 2752 9528 2753
rect 9208 2688 9216 2752
rect 9280 2688 9296 2752
rect 9360 2688 9376 2752
rect 9440 2688 9456 2752
rect 9520 2688 9528 2752
rect 9208 2687 9528 2688
rect 13077 2684 13143 2685
rect 13813 2684 13879 2685
rect 13077 2680 13124 2684
rect 13188 2682 13194 2684
rect 13077 2624 13082 2680
rect 13077 2620 13124 2624
rect 13188 2622 13234 2682
rect 13813 2680 13860 2684
rect 13924 2682 13930 2684
rect 14046 2682 14106 2894
rect 18873 2952 19215 2954
rect 18873 2896 18878 2952
rect 18934 2896 19154 2952
rect 19210 2896 19215 2952
rect 18873 2894 19215 2896
rect 18873 2891 18939 2894
rect 19149 2891 19215 2894
rect 24208 2918 24216 2982
rect 24280 2918 24296 2982
rect 24360 2918 24376 2982
rect 24440 2918 24456 2982
rect 24520 2918 24528 2982
rect 47718 2957 47778 3166
rect 50889 3224 51139 3226
rect 50889 3168 50894 3224
rect 50950 3168 51078 3224
rect 51134 3168 51139 3224
rect 50889 3166 51139 3168
rect 67406 3224 67515 3229
rect 67406 3168 67454 3224
rect 67510 3168 67515 3224
rect 67406 3166 67515 3168
rect 50889 3163 50955 3166
rect 51073 3163 51139 3166
rect 67449 3163 67515 3166
rect 68093 3226 68159 3229
rect 69200 3226 70000 3256
rect 68093 3224 70000 3226
rect 68093 3168 68098 3224
rect 68154 3168 70000 3224
rect 68093 3166 70000 3168
rect 68093 3163 68159 3166
rect 69200 3136 70000 3166
rect 48681 3090 48747 3093
rect 48681 3088 49802 3090
rect 48681 3032 48686 3088
rect 48742 3032 49802 3088
rect 48681 3030 49802 3032
rect 48681 3027 48747 3030
rect 24208 2902 24528 2918
rect 24208 2838 24216 2902
rect 24280 2838 24296 2902
rect 24360 2838 24376 2902
rect 24440 2838 24456 2902
rect 24520 2838 24528 2902
rect 33910 2892 33916 2956
rect 33980 2954 33986 2956
rect 41045 2954 41111 2957
rect 33980 2952 41111 2954
rect 33980 2896 41050 2952
rect 41106 2896 41111 2952
rect 33980 2894 41111 2896
rect 47718 2952 47827 2957
rect 47718 2896 47766 2952
rect 47822 2896 47827 2952
rect 47718 2894 47827 2896
rect 33980 2892 33986 2894
rect 41045 2891 41111 2894
rect 47761 2891 47827 2894
rect 14917 2818 14983 2821
rect 16205 2818 16271 2821
rect 14917 2816 16271 2818
rect 14917 2760 14922 2816
rect 14978 2760 16210 2816
rect 16266 2760 16271 2816
rect 14917 2758 16271 2760
rect 14917 2755 14983 2758
rect 16205 2755 16271 2758
rect 18321 2818 18387 2821
rect 18873 2818 18939 2821
rect 18321 2816 18939 2818
rect 18321 2760 18326 2816
rect 18382 2760 18878 2816
rect 18934 2760 18939 2816
rect 24208 2800 24528 2838
rect 34697 2818 34763 2821
rect 35065 2818 35131 2821
rect 34697 2816 35131 2818
rect 18321 2758 18939 2760
rect 18321 2755 18387 2758
rect 18873 2755 18939 2758
rect 34697 2760 34702 2816
rect 34758 2760 35070 2816
rect 35126 2760 35131 2816
rect 34697 2758 35131 2760
rect 34697 2755 34763 2758
rect 35065 2755 35131 2758
rect 40125 2818 40191 2821
rect 41965 2818 42031 2821
rect 40125 2816 42031 2818
rect 40125 2760 40130 2816
rect 40186 2760 41970 2816
rect 42026 2760 42031 2816
rect 40125 2758 42031 2760
rect 40125 2755 40191 2758
rect 41965 2755 42031 2758
rect 43161 2818 43227 2821
rect 43529 2818 43595 2821
rect 43161 2816 43595 2818
rect 43161 2760 43166 2816
rect 43222 2760 43534 2816
rect 43590 2760 43595 2816
rect 43161 2758 43595 2760
rect 43161 2755 43227 2758
rect 43529 2755 43595 2758
rect 44541 2818 44607 2821
rect 44950 2818 44956 2820
rect 44541 2816 44956 2818
rect 44541 2760 44546 2816
rect 44602 2760 44956 2816
rect 44541 2758 44956 2760
rect 44541 2755 44607 2758
rect 44950 2756 44956 2758
rect 45020 2756 45026 2820
rect 49049 2818 49115 2821
rect 48638 2816 49115 2818
rect 48638 2760 49054 2816
rect 49110 2760 49115 2816
rect 48638 2758 49115 2760
rect 39208 2752 39528 2753
rect 39208 2688 39216 2752
rect 39280 2688 39296 2752
rect 39360 2688 39376 2752
rect 39440 2688 39456 2752
rect 39520 2688 39528 2752
rect 39208 2687 39528 2688
rect 15193 2682 15259 2685
rect 13813 2624 13818 2680
rect 13188 2620 13194 2622
rect 13813 2620 13860 2624
rect 13924 2622 13970 2682
rect 14046 2680 15259 2682
rect 14046 2624 15198 2680
rect 15254 2624 15259 2680
rect 14046 2622 15259 2624
rect 13924 2620 13930 2622
rect 13077 2619 13143 2620
rect 13813 2619 13879 2620
rect 15193 2619 15259 2622
rect 18321 2682 18387 2685
rect 18873 2682 18939 2685
rect 18321 2680 18939 2682
rect 18321 2624 18326 2680
rect 18382 2624 18878 2680
rect 18934 2624 18939 2680
rect 18321 2622 18939 2624
rect 18321 2619 18387 2622
rect 18873 2619 18939 2622
rect 42425 2682 42491 2685
rect 42558 2682 42564 2684
rect 42425 2680 42564 2682
rect 42425 2624 42430 2680
rect 42486 2624 42564 2680
rect 42425 2622 42564 2624
rect 42425 2619 42491 2622
rect 42558 2620 42564 2622
rect 42628 2620 42634 2684
rect 38745 2546 38811 2549
rect 41597 2546 41663 2549
rect 38745 2544 41663 2546
rect 38745 2488 38750 2544
rect 38806 2488 41602 2544
rect 41658 2488 41663 2544
rect 38745 2486 41663 2488
rect 38745 2483 38811 2486
rect 41597 2483 41663 2486
rect 48497 2546 48563 2549
rect 48638 2546 48698 2758
rect 49049 2755 49115 2758
rect 49208 2752 49528 2753
rect 49208 2688 49216 2752
rect 49280 2688 49296 2752
rect 49360 2688 49376 2752
rect 49440 2688 49456 2752
rect 49520 2688 49528 2752
rect 49208 2687 49528 2688
rect 48497 2544 48698 2546
rect 48497 2488 48502 2544
rect 48558 2488 48698 2544
rect 48497 2486 48698 2488
rect 49742 2549 49802 3030
rect 49969 2954 50035 2957
rect 49926 2952 50035 2954
rect 49926 2896 49974 2952
rect 50030 2896 50035 2952
rect 49926 2891 50035 2896
rect 49742 2544 49851 2549
rect 49742 2488 49790 2544
rect 49846 2488 49851 2544
rect 49742 2486 49851 2488
rect 48497 2483 48563 2486
rect 49785 2483 49851 2486
rect 29208 2430 29528 2460
rect 29208 2366 29216 2430
rect 29280 2366 29296 2430
rect 29360 2366 29376 2430
rect 29440 2366 29456 2430
rect 29520 2366 29528 2430
rect 29208 2350 29528 2366
rect 29208 2286 29216 2350
rect 29280 2286 29296 2350
rect 29360 2286 29376 2350
rect 29440 2286 29456 2350
rect 29520 2286 29528 2350
rect 36629 2410 36695 2413
rect 42333 2410 42399 2413
rect 36629 2408 42399 2410
rect 36629 2352 36634 2408
rect 36690 2352 42338 2408
rect 42394 2352 42399 2408
rect 36629 2350 42399 2352
rect 36629 2347 36695 2350
rect 42333 2347 42399 2350
rect 48865 2410 48931 2413
rect 49926 2410 49986 2891
rect 59208 2752 59528 2753
rect 59208 2688 59216 2752
rect 59280 2688 59296 2752
rect 59360 2688 59376 2752
rect 59440 2688 59456 2752
rect 59520 2688 59528 2752
rect 59208 2687 59528 2688
rect 52269 2546 52335 2549
rect 53598 2546 53604 2548
rect 52269 2544 53604 2546
rect 52269 2488 52274 2544
rect 52330 2488 53604 2544
rect 52269 2486 53604 2488
rect 52269 2483 52335 2486
rect 53598 2484 53604 2486
rect 53668 2484 53674 2548
rect 48865 2408 49986 2410
rect 48865 2352 48870 2408
rect 48926 2352 49986 2408
rect 48865 2350 49986 2352
rect 48865 2347 48931 2350
rect 29208 2270 29528 2286
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 14208 2208 14528 2209
rect 14208 2144 14216 2208
rect 14280 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14528 2208
rect 29208 2206 29216 2270
rect 29280 2206 29296 2270
rect 29360 2206 29376 2270
rect 29440 2206 29456 2270
rect 29520 2206 29528 2270
rect 39205 2274 39271 2277
rect 42006 2274 42012 2276
rect 39205 2272 42012 2274
rect 39205 2216 39210 2272
rect 39266 2216 42012 2272
rect 39205 2214 42012 2216
rect 39205 2211 39271 2214
rect 42006 2212 42012 2214
rect 42076 2212 42082 2276
rect 49417 2274 49483 2277
rect 49734 2274 49740 2276
rect 49417 2272 49740 2274
rect 49417 2216 49422 2272
rect 49478 2216 49740 2272
rect 49417 2214 49740 2216
rect 49417 2211 49483 2214
rect 49734 2212 49740 2214
rect 49804 2212 49810 2276
rect 29208 2176 29528 2206
rect 44208 2208 44528 2209
rect 14208 2143 14528 2144
rect 44208 2144 44216 2208
rect 44280 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44528 2208
rect 44208 2143 44528 2144
rect 54208 2208 54528 2209
rect 54208 2144 54216 2208
rect 54280 2144 54296 2208
rect 54360 2144 54376 2208
rect 54440 2144 54456 2208
rect 54520 2144 54528 2208
rect 54208 2143 54528 2144
rect 64208 2208 64528 2209
rect 64208 2144 64216 2208
rect 64280 2144 64296 2208
rect 64360 2144 64376 2208
rect 64440 2144 64456 2208
rect 64520 2144 64528 2208
rect 64208 2143 64528 2144
rect 4521 2002 4587 2005
rect 5390 2002 5396 2004
rect 4521 2000 5396 2002
rect 4521 1944 4526 2000
rect 4582 1944 5396 2000
rect 4521 1942 5396 1944
rect 4521 1939 4587 1942
rect 5390 1940 5396 1942
rect 5460 1940 5466 2004
rect 38653 2002 38719 2005
rect 46606 2002 46612 2004
rect 38653 2000 46612 2002
rect 38653 1944 38658 2000
rect 38714 1944 46612 2000
rect 38653 1942 46612 1944
rect 38653 1939 38719 1942
rect 46606 1940 46612 1942
rect 46676 1940 46682 2004
rect 54385 2002 54451 2005
rect 54886 2002 54892 2004
rect 54385 2000 54892 2002
rect 54385 1944 54390 2000
rect 54446 1944 54892 2000
rect 54385 1942 54892 1944
rect 54385 1939 54451 1942
rect 54886 1940 54892 1942
rect 54956 1940 54962 2004
rect 64321 2002 64387 2005
rect 64638 2002 64644 2004
rect 64321 2000 64644 2002
rect 64321 1944 64326 2000
rect 64382 1944 64644 2000
rect 64321 1942 64644 1944
rect 64321 1939 64387 1942
rect 64638 1940 64644 1942
rect 64708 1940 64714 2004
rect 0 1866 800 1896
rect 1853 1866 1919 1869
rect 27705 1868 27771 1869
rect 28073 1868 28139 1869
rect 0 1864 1919 1866
rect 0 1808 1858 1864
rect 1914 1808 1919 1864
rect 0 1806 1919 1808
rect 0 1776 800 1806
rect 1853 1803 1919 1806
rect 27654 1804 27660 1868
rect 27724 1866 27771 1868
rect 27724 1864 27816 1866
rect 27766 1808 27816 1864
rect 27724 1806 27816 1808
rect 27724 1804 27771 1806
rect 28022 1804 28028 1868
rect 28092 1866 28139 1868
rect 29913 1866 29979 1869
rect 30046 1866 30052 1868
rect 28092 1864 28184 1866
rect 28134 1808 28184 1864
rect 28092 1806 28184 1808
rect 29913 1864 30052 1866
rect 29913 1808 29918 1864
rect 29974 1808 30052 1864
rect 29913 1806 30052 1808
rect 28092 1804 28139 1806
rect 27705 1803 27771 1804
rect 28073 1803 28139 1804
rect 29913 1803 29979 1806
rect 30046 1804 30052 1806
rect 30116 1804 30122 1868
rect 30189 1866 30255 1869
rect 30414 1866 30420 1868
rect 30189 1864 30420 1866
rect 30189 1808 30194 1864
rect 30250 1808 30420 1864
rect 30189 1806 30420 1808
rect 30189 1803 30255 1806
rect 30414 1804 30420 1806
rect 30484 1804 30490 1868
rect 31017 1866 31083 1869
rect 31150 1866 31156 1868
rect 31017 1864 31156 1866
rect 31017 1808 31022 1864
rect 31078 1808 31156 1864
rect 31017 1806 31156 1808
rect 31017 1803 31083 1806
rect 31150 1804 31156 1806
rect 31220 1804 31226 1868
rect 68185 1866 68251 1869
rect 69200 1866 70000 1896
rect 68185 1864 70000 1866
rect 68185 1808 68190 1864
rect 68246 1808 70000 1864
rect 68185 1806 70000 1808
rect 68185 1803 68251 1806
rect 69200 1776 70000 1806
rect 28165 1732 28231 1733
rect 28165 1730 28212 1732
rect 28120 1728 28212 1730
rect 28120 1672 28170 1728
rect 28120 1670 28212 1672
rect 28165 1668 28212 1670
rect 28276 1668 28282 1732
rect 28901 1730 28967 1733
rect 30598 1730 30604 1732
rect 28901 1728 30604 1730
rect 28901 1672 28906 1728
rect 28962 1672 30604 1728
rect 28901 1670 30604 1672
rect 28165 1667 28231 1668
rect 28901 1667 28967 1670
rect 30598 1668 30604 1670
rect 30668 1668 30674 1732
rect 39481 1322 39547 1325
rect 41270 1322 41276 1324
rect 39481 1320 41276 1322
rect 39481 1264 39486 1320
rect 39542 1264 41276 1320
rect 39481 1262 41276 1264
rect 39481 1259 39547 1262
rect 41270 1260 41276 1262
rect 41340 1260 41346 1324
rect 31845 1188 31911 1189
rect 31845 1186 31892 1188
rect 31800 1184 31892 1186
rect 31800 1128 31850 1184
rect 31800 1126 31892 1128
rect 31845 1124 31892 1126
rect 31956 1124 31962 1188
rect 31845 1123 31911 1124
rect 0 642 800 672
rect 2865 642 2931 645
rect 0 640 2931 642
rect 0 584 2870 640
rect 2926 584 2931 640
rect 0 582 2931 584
rect 0 552 800 582
rect 2865 579 2931 582
rect 66069 642 66135 645
rect 69200 642 70000 672
rect 66069 640 70000 642
rect 66069 584 66074 640
rect 66130 584 70000 640
rect 66069 582 70000 584
rect 66069 579 66135 582
rect 69200 552 70000 582
<< via3 >>
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 14216 67484 14280 67488
rect 14216 67428 14220 67484
rect 14220 67428 14276 67484
rect 14276 67428 14280 67484
rect 14216 67424 14280 67428
rect 14296 67484 14360 67488
rect 14296 67428 14300 67484
rect 14300 67428 14356 67484
rect 14356 67428 14360 67484
rect 14296 67424 14360 67428
rect 14376 67484 14440 67488
rect 14376 67428 14380 67484
rect 14380 67428 14436 67484
rect 14436 67428 14440 67484
rect 14376 67424 14440 67428
rect 14456 67484 14520 67488
rect 14456 67428 14460 67484
rect 14460 67428 14516 67484
rect 14516 67428 14520 67484
rect 14456 67424 14520 67428
rect 24216 67484 24280 67488
rect 24216 67428 24220 67484
rect 24220 67428 24276 67484
rect 24276 67428 24280 67484
rect 24216 67424 24280 67428
rect 24296 67484 24360 67488
rect 24296 67428 24300 67484
rect 24300 67428 24356 67484
rect 24356 67428 24360 67484
rect 24296 67424 24360 67428
rect 24376 67484 24440 67488
rect 24376 67428 24380 67484
rect 24380 67428 24436 67484
rect 24436 67428 24440 67484
rect 24376 67424 24440 67428
rect 24456 67484 24520 67488
rect 24456 67428 24460 67484
rect 24460 67428 24516 67484
rect 24516 67428 24520 67484
rect 24456 67424 24520 67428
rect 34216 67484 34280 67488
rect 34216 67428 34220 67484
rect 34220 67428 34276 67484
rect 34276 67428 34280 67484
rect 34216 67424 34280 67428
rect 34296 67484 34360 67488
rect 34296 67428 34300 67484
rect 34300 67428 34356 67484
rect 34356 67428 34360 67484
rect 34296 67424 34360 67428
rect 34376 67484 34440 67488
rect 34376 67428 34380 67484
rect 34380 67428 34436 67484
rect 34436 67428 34440 67484
rect 34376 67424 34440 67428
rect 34456 67484 34520 67488
rect 34456 67428 34460 67484
rect 34460 67428 34516 67484
rect 34516 67428 34520 67484
rect 34456 67424 34520 67428
rect 44216 67484 44280 67488
rect 44216 67428 44220 67484
rect 44220 67428 44276 67484
rect 44276 67428 44280 67484
rect 44216 67424 44280 67428
rect 44296 67484 44360 67488
rect 44296 67428 44300 67484
rect 44300 67428 44356 67484
rect 44356 67428 44360 67484
rect 44296 67424 44360 67428
rect 44376 67484 44440 67488
rect 44376 67428 44380 67484
rect 44380 67428 44436 67484
rect 44436 67428 44440 67484
rect 44376 67424 44440 67428
rect 44456 67484 44520 67488
rect 44456 67428 44460 67484
rect 44460 67428 44516 67484
rect 44516 67428 44520 67484
rect 44456 67424 44520 67428
rect 54216 67484 54280 67488
rect 54216 67428 54220 67484
rect 54220 67428 54276 67484
rect 54276 67428 54280 67484
rect 54216 67424 54280 67428
rect 54296 67484 54360 67488
rect 54296 67428 54300 67484
rect 54300 67428 54356 67484
rect 54356 67428 54360 67484
rect 54296 67424 54360 67428
rect 54376 67484 54440 67488
rect 54376 67428 54380 67484
rect 54380 67428 54436 67484
rect 54436 67428 54440 67484
rect 54376 67424 54440 67428
rect 54456 67484 54520 67488
rect 54456 67428 54460 67484
rect 54460 67428 54516 67484
rect 54516 67428 54520 67484
rect 54456 67424 54520 67428
rect 64216 67484 64280 67488
rect 64216 67428 64220 67484
rect 64220 67428 64276 67484
rect 64276 67428 64280 67484
rect 64216 67424 64280 67428
rect 64296 67484 64360 67488
rect 64296 67428 64300 67484
rect 64300 67428 64356 67484
rect 64356 67428 64360 67484
rect 64296 67424 64360 67428
rect 64376 67484 64440 67488
rect 64376 67428 64380 67484
rect 64380 67428 64436 67484
rect 64436 67428 64440 67484
rect 64376 67424 64440 67428
rect 64456 67484 64520 67488
rect 64456 67428 64460 67484
rect 64460 67428 64516 67484
rect 64516 67428 64520 67484
rect 64456 67424 64520 67428
rect 9216 66940 9280 66944
rect 9216 66884 9220 66940
rect 9220 66884 9276 66940
rect 9276 66884 9280 66940
rect 9216 66880 9280 66884
rect 9296 66940 9360 66944
rect 9296 66884 9300 66940
rect 9300 66884 9356 66940
rect 9356 66884 9360 66940
rect 9296 66880 9360 66884
rect 9376 66940 9440 66944
rect 9376 66884 9380 66940
rect 9380 66884 9436 66940
rect 9436 66884 9440 66940
rect 9376 66880 9440 66884
rect 9456 66940 9520 66944
rect 9456 66884 9460 66940
rect 9460 66884 9516 66940
rect 9516 66884 9520 66940
rect 9456 66880 9520 66884
rect 19216 66940 19280 66944
rect 19216 66884 19220 66940
rect 19220 66884 19276 66940
rect 19276 66884 19280 66940
rect 19216 66880 19280 66884
rect 19296 66940 19360 66944
rect 19296 66884 19300 66940
rect 19300 66884 19356 66940
rect 19356 66884 19360 66940
rect 19296 66880 19360 66884
rect 19376 66940 19440 66944
rect 19376 66884 19380 66940
rect 19380 66884 19436 66940
rect 19436 66884 19440 66940
rect 19376 66880 19440 66884
rect 19456 66940 19520 66944
rect 19456 66884 19460 66940
rect 19460 66884 19516 66940
rect 19516 66884 19520 66940
rect 19456 66880 19520 66884
rect 29216 66940 29280 66944
rect 29216 66884 29220 66940
rect 29220 66884 29276 66940
rect 29276 66884 29280 66940
rect 29216 66880 29280 66884
rect 29296 66940 29360 66944
rect 29296 66884 29300 66940
rect 29300 66884 29356 66940
rect 29356 66884 29360 66940
rect 29296 66880 29360 66884
rect 29376 66940 29440 66944
rect 29376 66884 29380 66940
rect 29380 66884 29436 66940
rect 29436 66884 29440 66940
rect 29376 66880 29440 66884
rect 29456 66940 29520 66944
rect 29456 66884 29460 66940
rect 29460 66884 29516 66940
rect 29516 66884 29520 66940
rect 29456 66880 29520 66884
rect 39216 66940 39280 66944
rect 39216 66884 39220 66940
rect 39220 66884 39276 66940
rect 39276 66884 39280 66940
rect 39216 66880 39280 66884
rect 39296 66940 39360 66944
rect 39296 66884 39300 66940
rect 39300 66884 39356 66940
rect 39356 66884 39360 66940
rect 39296 66880 39360 66884
rect 39376 66940 39440 66944
rect 39376 66884 39380 66940
rect 39380 66884 39436 66940
rect 39436 66884 39440 66940
rect 39376 66880 39440 66884
rect 39456 66940 39520 66944
rect 39456 66884 39460 66940
rect 39460 66884 39516 66940
rect 39516 66884 39520 66940
rect 39456 66880 39520 66884
rect 49216 66940 49280 66944
rect 49216 66884 49220 66940
rect 49220 66884 49276 66940
rect 49276 66884 49280 66940
rect 49216 66880 49280 66884
rect 49296 66940 49360 66944
rect 49296 66884 49300 66940
rect 49300 66884 49356 66940
rect 49356 66884 49360 66940
rect 49296 66880 49360 66884
rect 49376 66940 49440 66944
rect 49376 66884 49380 66940
rect 49380 66884 49436 66940
rect 49436 66884 49440 66940
rect 49376 66880 49440 66884
rect 49456 66940 49520 66944
rect 49456 66884 49460 66940
rect 49460 66884 49516 66940
rect 49516 66884 49520 66940
rect 49456 66880 49520 66884
rect 59216 66940 59280 66944
rect 59216 66884 59220 66940
rect 59220 66884 59276 66940
rect 59276 66884 59280 66940
rect 59216 66880 59280 66884
rect 59296 66940 59360 66944
rect 59296 66884 59300 66940
rect 59300 66884 59356 66940
rect 59356 66884 59360 66940
rect 59296 66880 59360 66884
rect 59376 66940 59440 66944
rect 59376 66884 59380 66940
rect 59380 66884 59436 66940
rect 59436 66884 59440 66940
rect 59376 66880 59440 66884
rect 59456 66940 59520 66944
rect 59456 66884 59460 66940
rect 59460 66884 59516 66940
rect 59516 66884 59520 66940
rect 59456 66880 59520 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 14216 66396 14280 66400
rect 14216 66340 14220 66396
rect 14220 66340 14276 66396
rect 14276 66340 14280 66396
rect 14216 66336 14280 66340
rect 14296 66396 14360 66400
rect 14296 66340 14300 66396
rect 14300 66340 14356 66396
rect 14356 66340 14360 66396
rect 14296 66336 14360 66340
rect 14376 66396 14440 66400
rect 14376 66340 14380 66396
rect 14380 66340 14436 66396
rect 14436 66340 14440 66396
rect 14376 66336 14440 66340
rect 14456 66396 14520 66400
rect 14456 66340 14460 66396
rect 14460 66340 14516 66396
rect 14516 66340 14520 66396
rect 14456 66336 14520 66340
rect 24216 66396 24280 66400
rect 24216 66340 24220 66396
rect 24220 66340 24276 66396
rect 24276 66340 24280 66396
rect 24216 66336 24280 66340
rect 24296 66396 24360 66400
rect 24296 66340 24300 66396
rect 24300 66340 24356 66396
rect 24356 66340 24360 66396
rect 24296 66336 24360 66340
rect 24376 66396 24440 66400
rect 24376 66340 24380 66396
rect 24380 66340 24436 66396
rect 24436 66340 24440 66396
rect 24376 66336 24440 66340
rect 24456 66396 24520 66400
rect 24456 66340 24460 66396
rect 24460 66340 24516 66396
rect 24516 66340 24520 66396
rect 24456 66336 24520 66340
rect 34216 66396 34280 66400
rect 34216 66340 34220 66396
rect 34220 66340 34276 66396
rect 34276 66340 34280 66396
rect 34216 66336 34280 66340
rect 34296 66396 34360 66400
rect 34296 66340 34300 66396
rect 34300 66340 34356 66396
rect 34356 66340 34360 66396
rect 34296 66336 34360 66340
rect 34376 66396 34440 66400
rect 34376 66340 34380 66396
rect 34380 66340 34436 66396
rect 34436 66340 34440 66396
rect 34376 66336 34440 66340
rect 34456 66396 34520 66400
rect 34456 66340 34460 66396
rect 34460 66340 34516 66396
rect 34516 66340 34520 66396
rect 34456 66336 34520 66340
rect 44216 66396 44280 66400
rect 44216 66340 44220 66396
rect 44220 66340 44276 66396
rect 44276 66340 44280 66396
rect 44216 66336 44280 66340
rect 44296 66396 44360 66400
rect 44296 66340 44300 66396
rect 44300 66340 44356 66396
rect 44356 66340 44360 66396
rect 44296 66336 44360 66340
rect 44376 66396 44440 66400
rect 44376 66340 44380 66396
rect 44380 66340 44436 66396
rect 44436 66340 44440 66396
rect 44376 66336 44440 66340
rect 44456 66396 44520 66400
rect 44456 66340 44460 66396
rect 44460 66340 44516 66396
rect 44516 66340 44520 66396
rect 44456 66336 44520 66340
rect 54216 66396 54280 66400
rect 54216 66340 54220 66396
rect 54220 66340 54276 66396
rect 54276 66340 54280 66396
rect 54216 66336 54280 66340
rect 54296 66396 54360 66400
rect 54296 66340 54300 66396
rect 54300 66340 54356 66396
rect 54356 66340 54360 66396
rect 54296 66336 54360 66340
rect 54376 66396 54440 66400
rect 54376 66340 54380 66396
rect 54380 66340 54436 66396
rect 54436 66340 54440 66396
rect 54376 66336 54440 66340
rect 54456 66396 54520 66400
rect 54456 66340 54460 66396
rect 54460 66340 54516 66396
rect 54516 66340 54520 66396
rect 54456 66336 54520 66340
rect 64216 66396 64280 66400
rect 64216 66340 64220 66396
rect 64220 66340 64276 66396
rect 64276 66340 64280 66396
rect 64216 66336 64280 66340
rect 64296 66396 64360 66400
rect 64296 66340 64300 66396
rect 64300 66340 64356 66396
rect 64356 66340 64360 66396
rect 64296 66336 64360 66340
rect 64376 66396 64440 66400
rect 64376 66340 64380 66396
rect 64380 66340 64436 66396
rect 64436 66340 64440 66396
rect 64376 66336 64440 66340
rect 64456 66396 64520 66400
rect 64456 66340 64460 66396
rect 64460 66340 64516 66396
rect 64516 66340 64520 66396
rect 64456 66336 64520 66340
rect 9216 65852 9280 65856
rect 9216 65796 9220 65852
rect 9220 65796 9276 65852
rect 9276 65796 9280 65852
rect 9216 65792 9280 65796
rect 9296 65852 9360 65856
rect 9296 65796 9300 65852
rect 9300 65796 9356 65852
rect 9356 65796 9360 65852
rect 9296 65792 9360 65796
rect 9376 65852 9440 65856
rect 9376 65796 9380 65852
rect 9380 65796 9436 65852
rect 9436 65796 9440 65852
rect 9376 65792 9440 65796
rect 9456 65852 9520 65856
rect 9456 65796 9460 65852
rect 9460 65796 9516 65852
rect 9516 65796 9520 65852
rect 9456 65792 9520 65796
rect 19216 65852 19280 65856
rect 19216 65796 19220 65852
rect 19220 65796 19276 65852
rect 19276 65796 19280 65852
rect 19216 65792 19280 65796
rect 19296 65852 19360 65856
rect 19296 65796 19300 65852
rect 19300 65796 19356 65852
rect 19356 65796 19360 65852
rect 19296 65792 19360 65796
rect 19376 65852 19440 65856
rect 19376 65796 19380 65852
rect 19380 65796 19436 65852
rect 19436 65796 19440 65852
rect 19376 65792 19440 65796
rect 19456 65852 19520 65856
rect 19456 65796 19460 65852
rect 19460 65796 19516 65852
rect 19516 65796 19520 65852
rect 19456 65792 19520 65796
rect 29216 65852 29280 65856
rect 29216 65796 29220 65852
rect 29220 65796 29276 65852
rect 29276 65796 29280 65852
rect 29216 65792 29280 65796
rect 29296 65852 29360 65856
rect 29296 65796 29300 65852
rect 29300 65796 29356 65852
rect 29356 65796 29360 65852
rect 29296 65792 29360 65796
rect 29376 65852 29440 65856
rect 29376 65796 29380 65852
rect 29380 65796 29436 65852
rect 29436 65796 29440 65852
rect 29376 65792 29440 65796
rect 29456 65852 29520 65856
rect 29456 65796 29460 65852
rect 29460 65796 29516 65852
rect 29516 65796 29520 65852
rect 29456 65792 29520 65796
rect 39216 65852 39280 65856
rect 39216 65796 39220 65852
rect 39220 65796 39276 65852
rect 39276 65796 39280 65852
rect 39216 65792 39280 65796
rect 39296 65852 39360 65856
rect 39296 65796 39300 65852
rect 39300 65796 39356 65852
rect 39356 65796 39360 65852
rect 39296 65792 39360 65796
rect 39376 65852 39440 65856
rect 39376 65796 39380 65852
rect 39380 65796 39436 65852
rect 39436 65796 39440 65852
rect 39376 65792 39440 65796
rect 39456 65852 39520 65856
rect 39456 65796 39460 65852
rect 39460 65796 39516 65852
rect 39516 65796 39520 65852
rect 39456 65792 39520 65796
rect 49216 65852 49280 65856
rect 49216 65796 49220 65852
rect 49220 65796 49276 65852
rect 49276 65796 49280 65852
rect 49216 65792 49280 65796
rect 49296 65852 49360 65856
rect 49296 65796 49300 65852
rect 49300 65796 49356 65852
rect 49356 65796 49360 65852
rect 49296 65792 49360 65796
rect 49376 65852 49440 65856
rect 49376 65796 49380 65852
rect 49380 65796 49436 65852
rect 49436 65796 49440 65852
rect 49376 65792 49440 65796
rect 49456 65852 49520 65856
rect 49456 65796 49460 65852
rect 49460 65796 49516 65852
rect 49516 65796 49520 65852
rect 49456 65792 49520 65796
rect 59216 65852 59280 65856
rect 59216 65796 59220 65852
rect 59220 65796 59276 65852
rect 59276 65796 59280 65852
rect 59216 65792 59280 65796
rect 59296 65852 59360 65856
rect 59296 65796 59300 65852
rect 59300 65796 59356 65852
rect 59356 65796 59360 65852
rect 59296 65792 59360 65796
rect 59376 65852 59440 65856
rect 59376 65796 59380 65852
rect 59380 65796 59436 65852
rect 59436 65796 59440 65852
rect 59376 65792 59440 65796
rect 59456 65852 59520 65856
rect 59456 65796 59460 65852
rect 59460 65796 59516 65852
rect 59516 65796 59520 65852
rect 59456 65792 59520 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 14216 65308 14280 65312
rect 14216 65252 14220 65308
rect 14220 65252 14276 65308
rect 14276 65252 14280 65308
rect 14216 65248 14280 65252
rect 14296 65308 14360 65312
rect 14296 65252 14300 65308
rect 14300 65252 14356 65308
rect 14356 65252 14360 65308
rect 14296 65248 14360 65252
rect 14376 65308 14440 65312
rect 14376 65252 14380 65308
rect 14380 65252 14436 65308
rect 14436 65252 14440 65308
rect 14376 65248 14440 65252
rect 14456 65308 14520 65312
rect 14456 65252 14460 65308
rect 14460 65252 14516 65308
rect 14516 65252 14520 65308
rect 14456 65248 14520 65252
rect 24216 65308 24280 65312
rect 24216 65252 24220 65308
rect 24220 65252 24276 65308
rect 24276 65252 24280 65308
rect 24216 65248 24280 65252
rect 24296 65308 24360 65312
rect 24296 65252 24300 65308
rect 24300 65252 24356 65308
rect 24356 65252 24360 65308
rect 24296 65248 24360 65252
rect 24376 65308 24440 65312
rect 24376 65252 24380 65308
rect 24380 65252 24436 65308
rect 24436 65252 24440 65308
rect 24376 65248 24440 65252
rect 24456 65308 24520 65312
rect 24456 65252 24460 65308
rect 24460 65252 24516 65308
rect 24516 65252 24520 65308
rect 24456 65248 24520 65252
rect 34216 65308 34280 65312
rect 34216 65252 34220 65308
rect 34220 65252 34276 65308
rect 34276 65252 34280 65308
rect 34216 65248 34280 65252
rect 34296 65308 34360 65312
rect 34296 65252 34300 65308
rect 34300 65252 34356 65308
rect 34356 65252 34360 65308
rect 34296 65248 34360 65252
rect 34376 65308 34440 65312
rect 34376 65252 34380 65308
rect 34380 65252 34436 65308
rect 34436 65252 34440 65308
rect 34376 65248 34440 65252
rect 34456 65308 34520 65312
rect 34456 65252 34460 65308
rect 34460 65252 34516 65308
rect 34516 65252 34520 65308
rect 34456 65248 34520 65252
rect 44216 65308 44280 65312
rect 44216 65252 44220 65308
rect 44220 65252 44276 65308
rect 44276 65252 44280 65308
rect 44216 65248 44280 65252
rect 44296 65308 44360 65312
rect 44296 65252 44300 65308
rect 44300 65252 44356 65308
rect 44356 65252 44360 65308
rect 44296 65248 44360 65252
rect 44376 65308 44440 65312
rect 44376 65252 44380 65308
rect 44380 65252 44436 65308
rect 44436 65252 44440 65308
rect 44376 65248 44440 65252
rect 44456 65308 44520 65312
rect 44456 65252 44460 65308
rect 44460 65252 44516 65308
rect 44516 65252 44520 65308
rect 44456 65248 44520 65252
rect 54216 65308 54280 65312
rect 54216 65252 54220 65308
rect 54220 65252 54276 65308
rect 54276 65252 54280 65308
rect 54216 65248 54280 65252
rect 54296 65308 54360 65312
rect 54296 65252 54300 65308
rect 54300 65252 54356 65308
rect 54356 65252 54360 65308
rect 54296 65248 54360 65252
rect 54376 65308 54440 65312
rect 54376 65252 54380 65308
rect 54380 65252 54436 65308
rect 54436 65252 54440 65308
rect 54376 65248 54440 65252
rect 54456 65308 54520 65312
rect 54456 65252 54460 65308
rect 54460 65252 54516 65308
rect 54516 65252 54520 65308
rect 54456 65248 54520 65252
rect 64216 65308 64280 65312
rect 64216 65252 64220 65308
rect 64220 65252 64276 65308
rect 64276 65252 64280 65308
rect 64216 65248 64280 65252
rect 64296 65308 64360 65312
rect 64296 65252 64300 65308
rect 64300 65252 64356 65308
rect 64356 65252 64360 65308
rect 64296 65248 64360 65252
rect 64376 65308 64440 65312
rect 64376 65252 64380 65308
rect 64380 65252 64436 65308
rect 64436 65252 64440 65308
rect 64376 65248 64440 65252
rect 64456 65308 64520 65312
rect 64456 65252 64460 65308
rect 64460 65252 64516 65308
rect 64516 65252 64520 65308
rect 64456 65248 64520 65252
rect 9216 64764 9280 64768
rect 9216 64708 9220 64764
rect 9220 64708 9276 64764
rect 9276 64708 9280 64764
rect 9216 64704 9280 64708
rect 9296 64764 9360 64768
rect 9296 64708 9300 64764
rect 9300 64708 9356 64764
rect 9356 64708 9360 64764
rect 9296 64704 9360 64708
rect 9376 64764 9440 64768
rect 9376 64708 9380 64764
rect 9380 64708 9436 64764
rect 9436 64708 9440 64764
rect 9376 64704 9440 64708
rect 9456 64764 9520 64768
rect 9456 64708 9460 64764
rect 9460 64708 9516 64764
rect 9516 64708 9520 64764
rect 9456 64704 9520 64708
rect 19216 64764 19280 64768
rect 19216 64708 19220 64764
rect 19220 64708 19276 64764
rect 19276 64708 19280 64764
rect 19216 64704 19280 64708
rect 19296 64764 19360 64768
rect 19296 64708 19300 64764
rect 19300 64708 19356 64764
rect 19356 64708 19360 64764
rect 19296 64704 19360 64708
rect 19376 64764 19440 64768
rect 19376 64708 19380 64764
rect 19380 64708 19436 64764
rect 19436 64708 19440 64764
rect 19376 64704 19440 64708
rect 19456 64764 19520 64768
rect 19456 64708 19460 64764
rect 19460 64708 19516 64764
rect 19516 64708 19520 64764
rect 19456 64704 19520 64708
rect 29216 64764 29280 64768
rect 29216 64708 29220 64764
rect 29220 64708 29276 64764
rect 29276 64708 29280 64764
rect 29216 64704 29280 64708
rect 29296 64764 29360 64768
rect 29296 64708 29300 64764
rect 29300 64708 29356 64764
rect 29356 64708 29360 64764
rect 29296 64704 29360 64708
rect 29376 64764 29440 64768
rect 29376 64708 29380 64764
rect 29380 64708 29436 64764
rect 29436 64708 29440 64764
rect 29376 64704 29440 64708
rect 29456 64764 29520 64768
rect 29456 64708 29460 64764
rect 29460 64708 29516 64764
rect 29516 64708 29520 64764
rect 29456 64704 29520 64708
rect 39216 64764 39280 64768
rect 39216 64708 39220 64764
rect 39220 64708 39276 64764
rect 39276 64708 39280 64764
rect 39216 64704 39280 64708
rect 39296 64764 39360 64768
rect 39296 64708 39300 64764
rect 39300 64708 39356 64764
rect 39356 64708 39360 64764
rect 39296 64704 39360 64708
rect 39376 64764 39440 64768
rect 39376 64708 39380 64764
rect 39380 64708 39436 64764
rect 39436 64708 39440 64764
rect 39376 64704 39440 64708
rect 39456 64764 39520 64768
rect 39456 64708 39460 64764
rect 39460 64708 39516 64764
rect 39516 64708 39520 64764
rect 39456 64704 39520 64708
rect 49216 64764 49280 64768
rect 49216 64708 49220 64764
rect 49220 64708 49276 64764
rect 49276 64708 49280 64764
rect 49216 64704 49280 64708
rect 49296 64764 49360 64768
rect 49296 64708 49300 64764
rect 49300 64708 49356 64764
rect 49356 64708 49360 64764
rect 49296 64704 49360 64708
rect 49376 64764 49440 64768
rect 49376 64708 49380 64764
rect 49380 64708 49436 64764
rect 49436 64708 49440 64764
rect 49376 64704 49440 64708
rect 49456 64764 49520 64768
rect 49456 64708 49460 64764
rect 49460 64708 49516 64764
rect 49516 64708 49520 64764
rect 49456 64704 49520 64708
rect 59216 64764 59280 64768
rect 59216 64708 59220 64764
rect 59220 64708 59276 64764
rect 59276 64708 59280 64764
rect 59216 64704 59280 64708
rect 59296 64764 59360 64768
rect 59296 64708 59300 64764
rect 59300 64708 59356 64764
rect 59356 64708 59360 64764
rect 59296 64704 59360 64708
rect 59376 64764 59440 64768
rect 59376 64708 59380 64764
rect 59380 64708 59436 64764
rect 59436 64708 59440 64764
rect 59376 64704 59440 64708
rect 59456 64764 59520 64768
rect 59456 64708 59460 64764
rect 59460 64708 59516 64764
rect 59516 64708 59520 64764
rect 59456 64704 59520 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 14216 64220 14280 64224
rect 14216 64164 14220 64220
rect 14220 64164 14276 64220
rect 14276 64164 14280 64220
rect 14216 64160 14280 64164
rect 14296 64220 14360 64224
rect 14296 64164 14300 64220
rect 14300 64164 14356 64220
rect 14356 64164 14360 64220
rect 14296 64160 14360 64164
rect 14376 64220 14440 64224
rect 14376 64164 14380 64220
rect 14380 64164 14436 64220
rect 14436 64164 14440 64220
rect 14376 64160 14440 64164
rect 14456 64220 14520 64224
rect 14456 64164 14460 64220
rect 14460 64164 14516 64220
rect 14516 64164 14520 64220
rect 14456 64160 14520 64164
rect 24216 64220 24280 64224
rect 24216 64164 24220 64220
rect 24220 64164 24276 64220
rect 24276 64164 24280 64220
rect 24216 64160 24280 64164
rect 24296 64220 24360 64224
rect 24296 64164 24300 64220
rect 24300 64164 24356 64220
rect 24356 64164 24360 64220
rect 24296 64160 24360 64164
rect 24376 64220 24440 64224
rect 24376 64164 24380 64220
rect 24380 64164 24436 64220
rect 24436 64164 24440 64220
rect 24376 64160 24440 64164
rect 24456 64220 24520 64224
rect 24456 64164 24460 64220
rect 24460 64164 24516 64220
rect 24516 64164 24520 64220
rect 24456 64160 24520 64164
rect 34216 64220 34280 64224
rect 34216 64164 34220 64220
rect 34220 64164 34276 64220
rect 34276 64164 34280 64220
rect 34216 64160 34280 64164
rect 34296 64220 34360 64224
rect 34296 64164 34300 64220
rect 34300 64164 34356 64220
rect 34356 64164 34360 64220
rect 34296 64160 34360 64164
rect 34376 64220 34440 64224
rect 34376 64164 34380 64220
rect 34380 64164 34436 64220
rect 34436 64164 34440 64220
rect 34376 64160 34440 64164
rect 34456 64220 34520 64224
rect 34456 64164 34460 64220
rect 34460 64164 34516 64220
rect 34516 64164 34520 64220
rect 34456 64160 34520 64164
rect 44216 64220 44280 64224
rect 44216 64164 44220 64220
rect 44220 64164 44276 64220
rect 44276 64164 44280 64220
rect 44216 64160 44280 64164
rect 44296 64220 44360 64224
rect 44296 64164 44300 64220
rect 44300 64164 44356 64220
rect 44356 64164 44360 64220
rect 44296 64160 44360 64164
rect 44376 64220 44440 64224
rect 44376 64164 44380 64220
rect 44380 64164 44436 64220
rect 44436 64164 44440 64220
rect 44376 64160 44440 64164
rect 44456 64220 44520 64224
rect 44456 64164 44460 64220
rect 44460 64164 44516 64220
rect 44516 64164 44520 64220
rect 44456 64160 44520 64164
rect 54216 64220 54280 64224
rect 54216 64164 54220 64220
rect 54220 64164 54276 64220
rect 54276 64164 54280 64220
rect 54216 64160 54280 64164
rect 54296 64220 54360 64224
rect 54296 64164 54300 64220
rect 54300 64164 54356 64220
rect 54356 64164 54360 64220
rect 54296 64160 54360 64164
rect 54376 64220 54440 64224
rect 54376 64164 54380 64220
rect 54380 64164 54436 64220
rect 54436 64164 54440 64220
rect 54376 64160 54440 64164
rect 54456 64220 54520 64224
rect 54456 64164 54460 64220
rect 54460 64164 54516 64220
rect 54516 64164 54520 64220
rect 54456 64160 54520 64164
rect 64216 64220 64280 64224
rect 64216 64164 64220 64220
rect 64220 64164 64276 64220
rect 64276 64164 64280 64220
rect 64216 64160 64280 64164
rect 64296 64220 64360 64224
rect 64296 64164 64300 64220
rect 64300 64164 64356 64220
rect 64356 64164 64360 64220
rect 64296 64160 64360 64164
rect 64376 64220 64440 64224
rect 64376 64164 64380 64220
rect 64380 64164 64436 64220
rect 64436 64164 64440 64220
rect 64376 64160 64440 64164
rect 64456 64220 64520 64224
rect 64456 64164 64460 64220
rect 64460 64164 64516 64220
rect 64516 64164 64520 64220
rect 64456 64160 64520 64164
rect 9216 63676 9280 63680
rect 9216 63620 9220 63676
rect 9220 63620 9276 63676
rect 9276 63620 9280 63676
rect 9216 63616 9280 63620
rect 9296 63676 9360 63680
rect 9296 63620 9300 63676
rect 9300 63620 9356 63676
rect 9356 63620 9360 63676
rect 9296 63616 9360 63620
rect 9376 63676 9440 63680
rect 9376 63620 9380 63676
rect 9380 63620 9436 63676
rect 9436 63620 9440 63676
rect 9376 63616 9440 63620
rect 9456 63676 9520 63680
rect 9456 63620 9460 63676
rect 9460 63620 9516 63676
rect 9516 63620 9520 63676
rect 9456 63616 9520 63620
rect 19216 63676 19280 63680
rect 19216 63620 19220 63676
rect 19220 63620 19276 63676
rect 19276 63620 19280 63676
rect 19216 63616 19280 63620
rect 19296 63676 19360 63680
rect 19296 63620 19300 63676
rect 19300 63620 19356 63676
rect 19356 63620 19360 63676
rect 19296 63616 19360 63620
rect 19376 63676 19440 63680
rect 19376 63620 19380 63676
rect 19380 63620 19436 63676
rect 19436 63620 19440 63676
rect 19376 63616 19440 63620
rect 19456 63676 19520 63680
rect 19456 63620 19460 63676
rect 19460 63620 19516 63676
rect 19516 63620 19520 63676
rect 19456 63616 19520 63620
rect 29216 63676 29280 63680
rect 29216 63620 29220 63676
rect 29220 63620 29276 63676
rect 29276 63620 29280 63676
rect 29216 63616 29280 63620
rect 29296 63676 29360 63680
rect 29296 63620 29300 63676
rect 29300 63620 29356 63676
rect 29356 63620 29360 63676
rect 29296 63616 29360 63620
rect 29376 63676 29440 63680
rect 29376 63620 29380 63676
rect 29380 63620 29436 63676
rect 29436 63620 29440 63676
rect 29376 63616 29440 63620
rect 29456 63676 29520 63680
rect 29456 63620 29460 63676
rect 29460 63620 29516 63676
rect 29516 63620 29520 63676
rect 29456 63616 29520 63620
rect 39216 63676 39280 63680
rect 39216 63620 39220 63676
rect 39220 63620 39276 63676
rect 39276 63620 39280 63676
rect 39216 63616 39280 63620
rect 39296 63676 39360 63680
rect 39296 63620 39300 63676
rect 39300 63620 39356 63676
rect 39356 63620 39360 63676
rect 39296 63616 39360 63620
rect 39376 63676 39440 63680
rect 39376 63620 39380 63676
rect 39380 63620 39436 63676
rect 39436 63620 39440 63676
rect 39376 63616 39440 63620
rect 39456 63676 39520 63680
rect 39456 63620 39460 63676
rect 39460 63620 39516 63676
rect 39516 63620 39520 63676
rect 39456 63616 39520 63620
rect 49216 63676 49280 63680
rect 49216 63620 49220 63676
rect 49220 63620 49276 63676
rect 49276 63620 49280 63676
rect 49216 63616 49280 63620
rect 49296 63676 49360 63680
rect 49296 63620 49300 63676
rect 49300 63620 49356 63676
rect 49356 63620 49360 63676
rect 49296 63616 49360 63620
rect 49376 63676 49440 63680
rect 49376 63620 49380 63676
rect 49380 63620 49436 63676
rect 49436 63620 49440 63676
rect 49376 63616 49440 63620
rect 49456 63676 49520 63680
rect 49456 63620 49460 63676
rect 49460 63620 49516 63676
rect 49516 63620 49520 63676
rect 49456 63616 49520 63620
rect 59216 63676 59280 63680
rect 59216 63620 59220 63676
rect 59220 63620 59276 63676
rect 59276 63620 59280 63676
rect 59216 63616 59280 63620
rect 59296 63676 59360 63680
rect 59296 63620 59300 63676
rect 59300 63620 59356 63676
rect 59356 63620 59360 63676
rect 59296 63616 59360 63620
rect 59376 63676 59440 63680
rect 59376 63620 59380 63676
rect 59380 63620 59436 63676
rect 59436 63620 59440 63676
rect 59376 63616 59440 63620
rect 59456 63676 59520 63680
rect 59456 63620 59460 63676
rect 59460 63620 59516 63676
rect 59516 63620 59520 63676
rect 59456 63616 59520 63620
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 14216 63132 14280 63136
rect 14216 63076 14220 63132
rect 14220 63076 14276 63132
rect 14276 63076 14280 63132
rect 14216 63072 14280 63076
rect 14296 63132 14360 63136
rect 14296 63076 14300 63132
rect 14300 63076 14356 63132
rect 14356 63076 14360 63132
rect 14296 63072 14360 63076
rect 14376 63132 14440 63136
rect 14376 63076 14380 63132
rect 14380 63076 14436 63132
rect 14436 63076 14440 63132
rect 14376 63072 14440 63076
rect 14456 63132 14520 63136
rect 14456 63076 14460 63132
rect 14460 63076 14516 63132
rect 14516 63076 14520 63132
rect 14456 63072 14520 63076
rect 24216 63132 24280 63136
rect 24216 63076 24220 63132
rect 24220 63076 24276 63132
rect 24276 63076 24280 63132
rect 24216 63072 24280 63076
rect 24296 63132 24360 63136
rect 24296 63076 24300 63132
rect 24300 63076 24356 63132
rect 24356 63076 24360 63132
rect 24296 63072 24360 63076
rect 24376 63132 24440 63136
rect 24376 63076 24380 63132
rect 24380 63076 24436 63132
rect 24436 63076 24440 63132
rect 24376 63072 24440 63076
rect 24456 63132 24520 63136
rect 24456 63076 24460 63132
rect 24460 63076 24516 63132
rect 24516 63076 24520 63132
rect 24456 63072 24520 63076
rect 34216 63132 34280 63136
rect 34216 63076 34220 63132
rect 34220 63076 34276 63132
rect 34276 63076 34280 63132
rect 34216 63072 34280 63076
rect 34296 63132 34360 63136
rect 34296 63076 34300 63132
rect 34300 63076 34356 63132
rect 34356 63076 34360 63132
rect 34296 63072 34360 63076
rect 34376 63132 34440 63136
rect 34376 63076 34380 63132
rect 34380 63076 34436 63132
rect 34436 63076 34440 63132
rect 34376 63072 34440 63076
rect 34456 63132 34520 63136
rect 34456 63076 34460 63132
rect 34460 63076 34516 63132
rect 34516 63076 34520 63132
rect 34456 63072 34520 63076
rect 44216 63132 44280 63136
rect 44216 63076 44220 63132
rect 44220 63076 44276 63132
rect 44276 63076 44280 63132
rect 44216 63072 44280 63076
rect 44296 63132 44360 63136
rect 44296 63076 44300 63132
rect 44300 63076 44356 63132
rect 44356 63076 44360 63132
rect 44296 63072 44360 63076
rect 44376 63132 44440 63136
rect 44376 63076 44380 63132
rect 44380 63076 44436 63132
rect 44436 63076 44440 63132
rect 44376 63072 44440 63076
rect 44456 63132 44520 63136
rect 44456 63076 44460 63132
rect 44460 63076 44516 63132
rect 44516 63076 44520 63132
rect 44456 63072 44520 63076
rect 54216 63132 54280 63136
rect 54216 63076 54220 63132
rect 54220 63076 54276 63132
rect 54276 63076 54280 63132
rect 54216 63072 54280 63076
rect 54296 63132 54360 63136
rect 54296 63076 54300 63132
rect 54300 63076 54356 63132
rect 54356 63076 54360 63132
rect 54296 63072 54360 63076
rect 54376 63132 54440 63136
rect 54376 63076 54380 63132
rect 54380 63076 54436 63132
rect 54436 63076 54440 63132
rect 54376 63072 54440 63076
rect 54456 63132 54520 63136
rect 54456 63076 54460 63132
rect 54460 63076 54516 63132
rect 54516 63076 54520 63132
rect 54456 63072 54520 63076
rect 64216 63132 64280 63136
rect 64216 63076 64220 63132
rect 64220 63076 64276 63132
rect 64276 63076 64280 63132
rect 64216 63072 64280 63076
rect 64296 63132 64360 63136
rect 64296 63076 64300 63132
rect 64300 63076 64356 63132
rect 64356 63076 64360 63132
rect 64296 63072 64360 63076
rect 64376 63132 64440 63136
rect 64376 63076 64380 63132
rect 64380 63076 64436 63132
rect 64436 63076 64440 63132
rect 64376 63072 64440 63076
rect 64456 63132 64520 63136
rect 64456 63076 64460 63132
rect 64460 63076 64516 63132
rect 64516 63076 64520 63132
rect 64456 63072 64520 63076
rect 9216 62588 9280 62592
rect 9216 62532 9220 62588
rect 9220 62532 9276 62588
rect 9276 62532 9280 62588
rect 9216 62528 9280 62532
rect 9296 62588 9360 62592
rect 9296 62532 9300 62588
rect 9300 62532 9356 62588
rect 9356 62532 9360 62588
rect 9296 62528 9360 62532
rect 9376 62588 9440 62592
rect 9376 62532 9380 62588
rect 9380 62532 9436 62588
rect 9436 62532 9440 62588
rect 9376 62528 9440 62532
rect 9456 62588 9520 62592
rect 9456 62532 9460 62588
rect 9460 62532 9516 62588
rect 9516 62532 9520 62588
rect 9456 62528 9520 62532
rect 19216 62588 19280 62592
rect 19216 62532 19220 62588
rect 19220 62532 19276 62588
rect 19276 62532 19280 62588
rect 19216 62528 19280 62532
rect 19296 62588 19360 62592
rect 19296 62532 19300 62588
rect 19300 62532 19356 62588
rect 19356 62532 19360 62588
rect 19296 62528 19360 62532
rect 19376 62588 19440 62592
rect 19376 62532 19380 62588
rect 19380 62532 19436 62588
rect 19436 62532 19440 62588
rect 19376 62528 19440 62532
rect 19456 62588 19520 62592
rect 19456 62532 19460 62588
rect 19460 62532 19516 62588
rect 19516 62532 19520 62588
rect 19456 62528 19520 62532
rect 29216 62588 29280 62592
rect 29216 62532 29220 62588
rect 29220 62532 29276 62588
rect 29276 62532 29280 62588
rect 29216 62528 29280 62532
rect 29296 62588 29360 62592
rect 29296 62532 29300 62588
rect 29300 62532 29356 62588
rect 29356 62532 29360 62588
rect 29296 62528 29360 62532
rect 29376 62588 29440 62592
rect 29376 62532 29380 62588
rect 29380 62532 29436 62588
rect 29436 62532 29440 62588
rect 29376 62528 29440 62532
rect 29456 62588 29520 62592
rect 29456 62532 29460 62588
rect 29460 62532 29516 62588
rect 29516 62532 29520 62588
rect 29456 62528 29520 62532
rect 39216 62588 39280 62592
rect 39216 62532 39220 62588
rect 39220 62532 39276 62588
rect 39276 62532 39280 62588
rect 39216 62528 39280 62532
rect 39296 62588 39360 62592
rect 39296 62532 39300 62588
rect 39300 62532 39356 62588
rect 39356 62532 39360 62588
rect 39296 62528 39360 62532
rect 39376 62588 39440 62592
rect 39376 62532 39380 62588
rect 39380 62532 39436 62588
rect 39436 62532 39440 62588
rect 39376 62528 39440 62532
rect 39456 62588 39520 62592
rect 39456 62532 39460 62588
rect 39460 62532 39516 62588
rect 39516 62532 39520 62588
rect 39456 62528 39520 62532
rect 49216 62588 49280 62592
rect 49216 62532 49220 62588
rect 49220 62532 49276 62588
rect 49276 62532 49280 62588
rect 49216 62528 49280 62532
rect 49296 62588 49360 62592
rect 49296 62532 49300 62588
rect 49300 62532 49356 62588
rect 49356 62532 49360 62588
rect 49296 62528 49360 62532
rect 49376 62588 49440 62592
rect 49376 62532 49380 62588
rect 49380 62532 49436 62588
rect 49436 62532 49440 62588
rect 49376 62528 49440 62532
rect 49456 62588 49520 62592
rect 49456 62532 49460 62588
rect 49460 62532 49516 62588
rect 49516 62532 49520 62588
rect 49456 62528 49520 62532
rect 59216 62588 59280 62592
rect 59216 62532 59220 62588
rect 59220 62532 59276 62588
rect 59276 62532 59280 62588
rect 59216 62528 59280 62532
rect 59296 62588 59360 62592
rect 59296 62532 59300 62588
rect 59300 62532 59356 62588
rect 59356 62532 59360 62588
rect 59296 62528 59360 62532
rect 59376 62588 59440 62592
rect 59376 62532 59380 62588
rect 59380 62532 59436 62588
rect 59436 62532 59440 62588
rect 59376 62528 59440 62532
rect 59456 62588 59520 62592
rect 59456 62532 59460 62588
rect 59460 62532 59516 62588
rect 59516 62532 59520 62588
rect 59456 62528 59520 62532
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 14216 62044 14280 62048
rect 14216 61988 14220 62044
rect 14220 61988 14276 62044
rect 14276 61988 14280 62044
rect 14216 61984 14280 61988
rect 14296 62044 14360 62048
rect 14296 61988 14300 62044
rect 14300 61988 14356 62044
rect 14356 61988 14360 62044
rect 14296 61984 14360 61988
rect 14376 62044 14440 62048
rect 14376 61988 14380 62044
rect 14380 61988 14436 62044
rect 14436 61988 14440 62044
rect 14376 61984 14440 61988
rect 14456 62044 14520 62048
rect 14456 61988 14460 62044
rect 14460 61988 14516 62044
rect 14516 61988 14520 62044
rect 14456 61984 14520 61988
rect 24216 62044 24280 62048
rect 24216 61988 24220 62044
rect 24220 61988 24276 62044
rect 24276 61988 24280 62044
rect 24216 61984 24280 61988
rect 24296 62044 24360 62048
rect 24296 61988 24300 62044
rect 24300 61988 24356 62044
rect 24356 61988 24360 62044
rect 24296 61984 24360 61988
rect 24376 62044 24440 62048
rect 24376 61988 24380 62044
rect 24380 61988 24436 62044
rect 24436 61988 24440 62044
rect 24376 61984 24440 61988
rect 24456 62044 24520 62048
rect 24456 61988 24460 62044
rect 24460 61988 24516 62044
rect 24516 61988 24520 62044
rect 24456 61984 24520 61988
rect 34216 62044 34280 62048
rect 34216 61988 34220 62044
rect 34220 61988 34276 62044
rect 34276 61988 34280 62044
rect 34216 61984 34280 61988
rect 34296 62044 34360 62048
rect 34296 61988 34300 62044
rect 34300 61988 34356 62044
rect 34356 61988 34360 62044
rect 34296 61984 34360 61988
rect 34376 62044 34440 62048
rect 34376 61988 34380 62044
rect 34380 61988 34436 62044
rect 34436 61988 34440 62044
rect 34376 61984 34440 61988
rect 34456 62044 34520 62048
rect 34456 61988 34460 62044
rect 34460 61988 34516 62044
rect 34516 61988 34520 62044
rect 34456 61984 34520 61988
rect 44216 62044 44280 62048
rect 44216 61988 44220 62044
rect 44220 61988 44276 62044
rect 44276 61988 44280 62044
rect 44216 61984 44280 61988
rect 44296 62044 44360 62048
rect 44296 61988 44300 62044
rect 44300 61988 44356 62044
rect 44356 61988 44360 62044
rect 44296 61984 44360 61988
rect 44376 62044 44440 62048
rect 44376 61988 44380 62044
rect 44380 61988 44436 62044
rect 44436 61988 44440 62044
rect 44376 61984 44440 61988
rect 44456 62044 44520 62048
rect 44456 61988 44460 62044
rect 44460 61988 44516 62044
rect 44516 61988 44520 62044
rect 44456 61984 44520 61988
rect 54216 62044 54280 62048
rect 54216 61988 54220 62044
rect 54220 61988 54276 62044
rect 54276 61988 54280 62044
rect 54216 61984 54280 61988
rect 54296 62044 54360 62048
rect 54296 61988 54300 62044
rect 54300 61988 54356 62044
rect 54356 61988 54360 62044
rect 54296 61984 54360 61988
rect 54376 62044 54440 62048
rect 54376 61988 54380 62044
rect 54380 61988 54436 62044
rect 54436 61988 54440 62044
rect 54376 61984 54440 61988
rect 54456 62044 54520 62048
rect 54456 61988 54460 62044
rect 54460 61988 54516 62044
rect 54516 61988 54520 62044
rect 54456 61984 54520 61988
rect 64216 62044 64280 62048
rect 64216 61988 64220 62044
rect 64220 61988 64276 62044
rect 64276 61988 64280 62044
rect 64216 61984 64280 61988
rect 64296 62044 64360 62048
rect 64296 61988 64300 62044
rect 64300 61988 64356 62044
rect 64356 61988 64360 62044
rect 64296 61984 64360 61988
rect 64376 62044 64440 62048
rect 64376 61988 64380 62044
rect 64380 61988 64436 62044
rect 64436 61988 64440 62044
rect 64376 61984 64440 61988
rect 64456 62044 64520 62048
rect 64456 61988 64460 62044
rect 64460 61988 64516 62044
rect 64516 61988 64520 62044
rect 64456 61984 64520 61988
rect 9216 61500 9280 61504
rect 9216 61444 9220 61500
rect 9220 61444 9276 61500
rect 9276 61444 9280 61500
rect 9216 61440 9280 61444
rect 9296 61500 9360 61504
rect 9296 61444 9300 61500
rect 9300 61444 9356 61500
rect 9356 61444 9360 61500
rect 9296 61440 9360 61444
rect 9376 61500 9440 61504
rect 9376 61444 9380 61500
rect 9380 61444 9436 61500
rect 9436 61444 9440 61500
rect 9376 61440 9440 61444
rect 9456 61500 9520 61504
rect 9456 61444 9460 61500
rect 9460 61444 9516 61500
rect 9516 61444 9520 61500
rect 9456 61440 9520 61444
rect 19216 61500 19280 61504
rect 19216 61444 19220 61500
rect 19220 61444 19276 61500
rect 19276 61444 19280 61500
rect 19216 61440 19280 61444
rect 19296 61500 19360 61504
rect 19296 61444 19300 61500
rect 19300 61444 19356 61500
rect 19356 61444 19360 61500
rect 19296 61440 19360 61444
rect 19376 61500 19440 61504
rect 19376 61444 19380 61500
rect 19380 61444 19436 61500
rect 19436 61444 19440 61500
rect 19376 61440 19440 61444
rect 19456 61500 19520 61504
rect 19456 61444 19460 61500
rect 19460 61444 19516 61500
rect 19516 61444 19520 61500
rect 19456 61440 19520 61444
rect 29216 61500 29280 61504
rect 29216 61444 29220 61500
rect 29220 61444 29276 61500
rect 29276 61444 29280 61500
rect 29216 61440 29280 61444
rect 29296 61500 29360 61504
rect 29296 61444 29300 61500
rect 29300 61444 29356 61500
rect 29356 61444 29360 61500
rect 29296 61440 29360 61444
rect 29376 61500 29440 61504
rect 29376 61444 29380 61500
rect 29380 61444 29436 61500
rect 29436 61444 29440 61500
rect 29376 61440 29440 61444
rect 29456 61500 29520 61504
rect 29456 61444 29460 61500
rect 29460 61444 29516 61500
rect 29516 61444 29520 61500
rect 29456 61440 29520 61444
rect 39216 61500 39280 61504
rect 39216 61444 39220 61500
rect 39220 61444 39276 61500
rect 39276 61444 39280 61500
rect 39216 61440 39280 61444
rect 39296 61500 39360 61504
rect 39296 61444 39300 61500
rect 39300 61444 39356 61500
rect 39356 61444 39360 61500
rect 39296 61440 39360 61444
rect 39376 61500 39440 61504
rect 39376 61444 39380 61500
rect 39380 61444 39436 61500
rect 39436 61444 39440 61500
rect 39376 61440 39440 61444
rect 39456 61500 39520 61504
rect 39456 61444 39460 61500
rect 39460 61444 39516 61500
rect 39516 61444 39520 61500
rect 39456 61440 39520 61444
rect 49216 61500 49280 61504
rect 49216 61444 49220 61500
rect 49220 61444 49276 61500
rect 49276 61444 49280 61500
rect 49216 61440 49280 61444
rect 49296 61500 49360 61504
rect 49296 61444 49300 61500
rect 49300 61444 49356 61500
rect 49356 61444 49360 61500
rect 49296 61440 49360 61444
rect 49376 61500 49440 61504
rect 49376 61444 49380 61500
rect 49380 61444 49436 61500
rect 49436 61444 49440 61500
rect 49376 61440 49440 61444
rect 49456 61500 49520 61504
rect 49456 61444 49460 61500
rect 49460 61444 49516 61500
rect 49516 61444 49520 61500
rect 49456 61440 49520 61444
rect 59216 61500 59280 61504
rect 59216 61444 59220 61500
rect 59220 61444 59276 61500
rect 59276 61444 59280 61500
rect 59216 61440 59280 61444
rect 59296 61500 59360 61504
rect 59296 61444 59300 61500
rect 59300 61444 59356 61500
rect 59356 61444 59360 61500
rect 59296 61440 59360 61444
rect 59376 61500 59440 61504
rect 59376 61444 59380 61500
rect 59380 61444 59436 61500
rect 59436 61444 59440 61500
rect 59376 61440 59440 61444
rect 59456 61500 59520 61504
rect 59456 61444 59460 61500
rect 59460 61444 59516 61500
rect 59516 61444 59520 61500
rect 59456 61440 59520 61444
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 14216 60956 14280 60960
rect 14216 60900 14220 60956
rect 14220 60900 14276 60956
rect 14276 60900 14280 60956
rect 14216 60896 14280 60900
rect 14296 60956 14360 60960
rect 14296 60900 14300 60956
rect 14300 60900 14356 60956
rect 14356 60900 14360 60956
rect 14296 60896 14360 60900
rect 14376 60956 14440 60960
rect 14376 60900 14380 60956
rect 14380 60900 14436 60956
rect 14436 60900 14440 60956
rect 14376 60896 14440 60900
rect 14456 60956 14520 60960
rect 14456 60900 14460 60956
rect 14460 60900 14516 60956
rect 14516 60900 14520 60956
rect 14456 60896 14520 60900
rect 24216 60956 24280 60960
rect 24216 60900 24220 60956
rect 24220 60900 24276 60956
rect 24276 60900 24280 60956
rect 24216 60896 24280 60900
rect 24296 60956 24360 60960
rect 24296 60900 24300 60956
rect 24300 60900 24356 60956
rect 24356 60900 24360 60956
rect 24296 60896 24360 60900
rect 24376 60956 24440 60960
rect 24376 60900 24380 60956
rect 24380 60900 24436 60956
rect 24436 60900 24440 60956
rect 24376 60896 24440 60900
rect 24456 60956 24520 60960
rect 24456 60900 24460 60956
rect 24460 60900 24516 60956
rect 24516 60900 24520 60956
rect 24456 60896 24520 60900
rect 34216 60956 34280 60960
rect 34216 60900 34220 60956
rect 34220 60900 34276 60956
rect 34276 60900 34280 60956
rect 34216 60896 34280 60900
rect 34296 60956 34360 60960
rect 34296 60900 34300 60956
rect 34300 60900 34356 60956
rect 34356 60900 34360 60956
rect 34296 60896 34360 60900
rect 34376 60956 34440 60960
rect 34376 60900 34380 60956
rect 34380 60900 34436 60956
rect 34436 60900 34440 60956
rect 34376 60896 34440 60900
rect 34456 60956 34520 60960
rect 34456 60900 34460 60956
rect 34460 60900 34516 60956
rect 34516 60900 34520 60956
rect 34456 60896 34520 60900
rect 44216 60956 44280 60960
rect 44216 60900 44220 60956
rect 44220 60900 44276 60956
rect 44276 60900 44280 60956
rect 44216 60896 44280 60900
rect 44296 60956 44360 60960
rect 44296 60900 44300 60956
rect 44300 60900 44356 60956
rect 44356 60900 44360 60956
rect 44296 60896 44360 60900
rect 44376 60956 44440 60960
rect 44376 60900 44380 60956
rect 44380 60900 44436 60956
rect 44436 60900 44440 60956
rect 44376 60896 44440 60900
rect 44456 60956 44520 60960
rect 44456 60900 44460 60956
rect 44460 60900 44516 60956
rect 44516 60900 44520 60956
rect 44456 60896 44520 60900
rect 54216 60956 54280 60960
rect 54216 60900 54220 60956
rect 54220 60900 54276 60956
rect 54276 60900 54280 60956
rect 54216 60896 54280 60900
rect 54296 60956 54360 60960
rect 54296 60900 54300 60956
rect 54300 60900 54356 60956
rect 54356 60900 54360 60956
rect 54296 60896 54360 60900
rect 54376 60956 54440 60960
rect 54376 60900 54380 60956
rect 54380 60900 54436 60956
rect 54436 60900 54440 60956
rect 54376 60896 54440 60900
rect 54456 60956 54520 60960
rect 54456 60900 54460 60956
rect 54460 60900 54516 60956
rect 54516 60900 54520 60956
rect 54456 60896 54520 60900
rect 64216 60956 64280 60960
rect 64216 60900 64220 60956
rect 64220 60900 64276 60956
rect 64276 60900 64280 60956
rect 64216 60896 64280 60900
rect 64296 60956 64360 60960
rect 64296 60900 64300 60956
rect 64300 60900 64356 60956
rect 64356 60900 64360 60956
rect 64296 60896 64360 60900
rect 64376 60956 64440 60960
rect 64376 60900 64380 60956
rect 64380 60900 64436 60956
rect 64436 60900 64440 60956
rect 64376 60896 64440 60900
rect 64456 60956 64520 60960
rect 64456 60900 64460 60956
rect 64460 60900 64516 60956
rect 64516 60900 64520 60956
rect 64456 60896 64520 60900
rect 9216 60412 9280 60416
rect 9216 60356 9220 60412
rect 9220 60356 9276 60412
rect 9276 60356 9280 60412
rect 9216 60352 9280 60356
rect 9296 60412 9360 60416
rect 9296 60356 9300 60412
rect 9300 60356 9356 60412
rect 9356 60356 9360 60412
rect 9296 60352 9360 60356
rect 9376 60412 9440 60416
rect 9376 60356 9380 60412
rect 9380 60356 9436 60412
rect 9436 60356 9440 60412
rect 9376 60352 9440 60356
rect 9456 60412 9520 60416
rect 9456 60356 9460 60412
rect 9460 60356 9516 60412
rect 9516 60356 9520 60412
rect 9456 60352 9520 60356
rect 19216 60412 19280 60416
rect 19216 60356 19220 60412
rect 19220 60356 19276 60412
rect 19276 60356 19280 60412
rect 19216 60352 19280 60356
rect 19296 60412 19360 60416
rect 19296 60356 19300 60412
rect 19300 60356 19356 60412
rect 19356 60356 19360 60412
rect 19296 60352 19360 60356
rect 19376 60412 19440 60416
rect 19376 60356 19380 60412
rect 19380 60356 19436 60412
rect 19436 60356 19440 60412
rect 19376 60352 19440 60356
rect 19456 60412 19520 60416
rect 19456 60356 19460 60412
rect 19460 60356 19516 60412
rect 19516 60356 19520 60412
rect 19456 60352 19520 60356
rect 29216 60412 29280 60416
rect 29216 60356 29220 60412
rect 29220 60356 29276 60412
rect 29276 60356 29280 60412
rect 29216 60352 29280 60356
rect 29296 60412 29360 60416
rect 29296 60356 29300 60412
rect 29300 60356 29356 60412
rect 29356 60356 29360 60412
rect 29296 60352 29360 60356
rect 29376 60412 29440 60416
rect 29376 60356 29380 60412
rect 29380 60356 29436 60412
rect 29436 60356 29440 60412
rect 29376 60352 29440 60356
rect 29456 60412 29520 60416
rect 29456 60356 29460 60412
rect 29460 60356 29516 60412
rect 29516 60356 29520 60412
rect 29456 60352 29520 60356
rect 39216 60412 39280 60416
rect 39216 60356 39220 60412
rect 39220 60356 39276 60412
rect 39276 60356 39280 60412
rect 39216 60352 39280 60356
rect 39296 60412 39360 60416
rect 39296 60356 39300 60412
rect 39300 60356 39356 60412
rect 39356 60356 39360 60412
rect 39296 60352 39360 60356
rect 39376 60412 39440 60416
rect 39376 60356 39380 60412
rect 39380 60356 39436 60412
rect 39436 60356 39440 60412
rect 39376 60352 39440 60356
rect 39456 60412 39520 60416
rect 39456 60356 39460 60412
rect 39460 60356 39516 60412
rect 39516 60356 39520 60412
rect 39456 60352 39520 60356
rect 49216 60412 49280 60416
rect 49216 60356 49220 60412
rect 49220 60356 49276 60412
rect 49276 60356 49280 60412
rect 49216 60352 49280 60356
rect 49296 60412 49360 60416
rect 49296 60356 49300 60412
rect 49300 60356 49356 60412
rect 49356 60356 49360 60412
rect 49296 60352 49360 60356
rect 49376 60412 49440 60416
rect 49376 60356 49380 60412
rect 49380 60356 49436 60412
rect 49436 60356 49440 60412
rect 49376 60352 49440 60356
rect 49456 60412 49520 60416
rect 49456 60356 49460 60412
rect 49460 60356 49516 60412
rect 49516 60356 49520 60412
rect 49456 60352 49520 60356
rect 59216 60412 59280 60416
rect 59216 60356 59220 60412
rect 59220 60356 59276 60412
rect 59276 60356 59280 60412
rect 59216 60352 59280 60356
rect 59296 60412 59360 60416
rect 59296 60356 59300 60412
rect 59300 60356 59356 60412
rect 59356 60356 59360 60412
rect 59296 60352 59360 60356
rect 59376 60412 59440 60416
rect 59376 60356 59380 60412
rect 59380 60356 59436 60412
rect 59436 60356 59440 60412
rect 59376 60352 59440 60356
rect 59456 60412 59520 60416
rect 59456 60356 59460 60412
rect 59460 60356 59516 60412
rect 59516 60356 59520 60412
rect 59456 60352 59520 60356
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 14216 59868 14280 59872
rect 14216 59812 14220 59868
rect 14220 59812 14276 59868
rect 14276 59812 14280 59868
rect 14216 59808 14280 59812
rect 14296 59868 14360 59872
rect 14296 59812 14300 59868
rect 14300 59812 14356 59868
rect 14356 59812 14360 59868
rect 14296 59808 14360 59812
rect 14376 59868 14440 59872
rect 14376 59812 14380 59868
rect 14380 59812 14436 59868
rect 14436 59812 14440 59868
rect 14376 59808 14440 59812
rect 14456 59868 14520 59872
rect 14456 59812 14460 59868
rect 14460 59812 14516 59868
rect 14516 59812 14520 59868
rect 14456 59808 14520 59812
rect 24216 59868 24280 59872
rect 24216 59812 24220 59868
rect 24220 59812 24276 59868
rect 24276 59812 24280 59868
rect 24216 59808 24280 59812
rect 24296 59868 24360 59872
rect 24296 59812 24300 59868
rect 24300 59812 24356 59868
rect 24356 59812 24360 59868
rect 24296 59808 24360 59812
rect 24376 59868 24440 59872
rect 24376 59812 24380 59868
rect 24380 59812 24436 59868
rect 24436 59812 24440 59868
rect 24376 59808 24440 59812
rect 24456 59868 24520 59872
rect 24456 59812 24460 59868
rect 24460 59812 24516 59868
rect 24516 59812 24520 59868
rect 24456 59808 24520 59812
rect 34216 59868 34280 59872
rect 34216 59812 34220 59868
rect 34220 59812 34276 59868
rect 34276 59812 34280 59868
rect 34216 59808 34280 59812
rect 34296 59868 34360 59872
rect 34296 59812 34300 59868
rect 34300 59812 34356 59868
rect 34356 59812 34360 59868
rect 34296 59808 34360 59812
rect 34376 59868 34440 59872
rect 34376 59812 34380 59868
rect 34380 59812 34436 59868
rect 34436 59812 34440 59868
rect 34376 59808 34440 59812
rect 34456 59868 34520 59872
rect 34456 59812 34460 59868
rect 34460 59812 34516 59868
rect 34516 59812 34520 59868
rect 34456 59808 34520 59812
rect 44216 59868 44280 59872
rect 44216 59812 44220 59868
rect 44220 59812 44276 59868
rect 44276 59812 44280 59868
rect 44216 59808 44280 59812
rect 44296 59868 44360 59872
rect 44296 59812 44300 59868
rect 44300 59812 44356 59868
rect 44356 59812 44360 59868
rect 44296 59808 44360 59812
rect 44376 59868 44440 59872
rect 44376 59812 44380 59868
rect 44380 59812 44436 59868
rect 44436 59812 44440 59868
rect 44376 59808 44440 59812
rect 44456 59868 44520 59872
rect 44456 59812 44460 59868
rect 44460 59812 44516 59868
rect 44516 59812 44520 59868
rect 44456 59808 44520 59812
rect 54216 59868 54280 59872
rect 54216 59812 54220 59868
rect 54220 59812 54276 59868
rect 54276 59812 54280 59868
rect 54216 59808 54280 59812
rect 54296 59868 54360 59872
rect 54296 59812 54300 59868
rect 54300 59812 54356 59868
rect 54356 59812 54360 59868
rect 54296 59808 54360 59812
rect 54376 59868 54440 59872
rect 54376 59812 54380 59868
rect 54380 59812 54436 59868
rect 54436 59812 54440 59868
rect 54376 59808 54440 59812
rect 54456 59868 54520 59872
rect 54456 59812 54460 59868
rect 54460 59812 54516 59868
rect 54516 59812 54520 59868
rect 54456 59808 54520 59812
rect 64216 59868 64280 59872
rect 64216 59812 64220 59868
rect 64220 59812 64276 59868
rect 64276 59812 64280 59868
rect 64216 59808 64280 59812
rect 64296 59868 64360 59872
rect 64296 59812 64300 59868
rect 64300 59812 64356 59868
rect 64356 59812 64360 59868
rect 64296 59808 64360 59812
rect 64376 59868 64440 59872
rect 64376 59812 64380 59868
rect 64380 59812 64436 59868
rect 64436 59812 64440 59868
rect 64376 59808 64440 59812
rect 64456 59868 64520 59872
rect 64456 59812 64460 59868
rect 64460 59812 64516 59868
rect 64516 59812 64520 59868
rect 64456 59808 64520 59812
rect 9216 59324 9280 59328
rect 9216 59268 9220 59324
rect 9220 59268 9276 59324
rect 9276 59268 9280 59324
rect 9216 59264 9280 59268
rect 9296 59324 9360 59328
rect 9296 59268 9300 59324
rect 9300 59268 9356 59324
rect 9356 59268 9360 59324
rect 9296 59264 9360 59268
rect 9376 59324 9440 59328
rect 9376 59268 9380 59324
rect 9380 59268 9436 59324
rect 9436 59268 9440 59324
rect 9376 59264 9440 59268
rect 9456 59324 9520 59328
rect 9456 59268 9460 59324
rect 9460 59268 9516 59324
rect 9516 59268 9520 59324
rect 9456 59264 9520 59268
rect 19216 59324 19280 59328
rect 19216 59268 19220 59324
rect 19220 59268 19276 59324
rect 19276 59268 19280 59324
rect 19216 59264 19280 59268
rect 19296 59324 19360 59328
rect 19296 59268 19300 59324
rect 19300 59268 19356 59324
rect 19356 59268 19360 59324
rect 19296 59264 19360 59268
rect 19376 59324 19440 59328
rect 19376 59268 19380 59324
rect 19380 59268 19436 59324
rect 19436 59268 19440 59324
rect 19376 59264 19440 59268
rect 19456 59324 19520 59328
rect 19456 59268 19460 59324
rect 19460 59268 19516 59324
rect 19516 59268 19520 59324
rect 19456 59264 19520 59268
rect 29216 59324 29280 59328
rect 29216 59268 29220 59324
rect 29220 59268 29276 59324
rect 29276 59268 29280 59324
rect 29216 59264 29280 59268
rect 29296 59324 29360 59328
rect 29296 59268 29300 59324
rect 29300 59268 29356 59324
rect 29356 59268 29360 59324
rect 29296 59264 29360 59268
rect 29376 59324 29440 59328
rect 29376 59268 29380 59324
rect 29380 59268 29436 59324
rect 29436 59268 29440 59324
rect 29376 59264 29440 59268
rect 29456 59324 29520 59328
rect 29456 59268 29460 59324
rect 29460 59268 29516 59324
rect 29516 59268 29520 59324
rect 29456 59264 29520 59268
rect 39216 59324 39280 59328
rect 39216 59268 39220 59324
rect 39220 59268 39276 59324
rect 39276 59268 39280 59324
rect 39216 59264 39280 59268
rect 39296 59324 39360 59328
rect 39296 59268 39300 59324
rect 39300 59268 39356 59324
rect 39356 59268 39360 59324
rect 39296 59264 39360 59268
rect 39376 59324 39440 59328
rect 39376 59268 39380 59324
rect 39380 59268 39436 59324
rect 39436 59268 39440 59324
rect 39376 59264 39440 59268
rect 39456 59324 39520 59328
rect 39456 59268 39460 59324
rect 39460 59268 39516 59324
rect 39516 59268 39520 59324
rect 39456 59264 39520 59268
rect 49216 59324 49280 59328
rect 49216 59268 49220 59324
rect 49220 59268 49276 59324
rect 49276 59268 49280 59324
rect 49216 59264 49280 59268
rect 49296 59324 49360 59328
rect 49296 59268 49300 59324
rect 49300 59268 49356 59324
rect 49356 59268 49360 59324
rect 49296 59264 49360 59268
rect 49376 59324 49440 59328
rect 49376 59268 49380 59324
rect 49380 59268 49436 59324
rect 49436 59268 49440 59324
rect 49376 59264 49440 59268
rect 49456 59324 49520 59328
rect 49456 59268 49460 59324
rect 49460 59268 49516 59324
rect 49516 59268 49520 59324
rect 49456 59264 49520 59268
rect 59216 59324 59280 59328
rect 59216 59268 59220 59324
rect 59220 59268 59276 59324
rect 59276 59268 59280 59324
rect 59216 59264 59280 59268
rect 59296 59324 59360 59328
rect 59296 59268 59300 59324
rect 59300 59268 59356 59324
rect 59356 59268 59360 59324
rect 59296 59264 59360 59268
rect 59376 59324 59440 59328
rect 59376 59268 59380 59324
rect 59380 59268 59436 59324
rect 59436 59268 59440 59324
rect 59376 59264 59440 59268
rect 59456 59324 59520 59328
rect 59456 59268 59460 59324
rect 59460 59268 59516 59324
rect 59516 59268 59520 59324
rect 59456 59264 59520 59268
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 14216 58780 14280 58784
rect 14216 58724 14220 58780
rect 14220 58724 14276 58780
rect 14276 58724 14280 58780
rect 14216 58720 14280 58724
rect 14296 58780 14360 58784
rect 14296 58724 14300 58780
rect 14300 58724 14356 58780
rect 14356 58724 14360 58780
rect 14296 58720 14360 58724
rect 14376 58780 14440 58784
rect 14376 58724 14380 58780
rect 14380 58724 14436 58780
rect 14436 58724 14440 58780
rect 14376 58720 14440 58724
rect 14456 58780 14520 58784
rect 14456 58724 14460 58780
rect 14460 58724 14516 58780
rect 14516 58724 14520 58780
rect 14456 58720 14520 58724
rect 24216 58780 24280 58784
rect 24216 58724 24220 58780
rect 24220 58724 24276 58780
rect 24276 58724 24280 58780
rect 24216 58720 24280 58724
rect 24296 58780 24360 58784
rect 24296 58724 24300 58780
rect 24300 58724 24356 58780
rect 24356 58724 24360 58780
rect 24296 58720 24360 58724
rect 24376 58780 24440 58784
rect 24376 58724 24380 58780
rect 24380 58724 24436 58780
rect 24436 58724 24440 58780
rect 24376 58720 24440 58724
rect 24456 58780 24520 58784
rect 24456 58724 24460 58780
rect 24460 58724 24516 58780
rect 24516 58724 24520 58780
rect 24456 58720 24520 58724
rect 34216 58780 34280 58784
rect 34216 58724 34220 58780
rect 34220 58724 34276 58780
rect 34276 58724 34280 58780
rect 34216 58720 34280 58724
rect 34296 58780 34360 58784
rect 34296 58724 34300 58780
rect 34300 58724 34356 58780
rect 34356 58724 34360 58780
rect 34296 58720 34360 58724
rect 34376 58780 34440 58784
rect 34376 58724 34380 58780
rect 34380 58724 34436 58780
rect 34436 58724 34440 58780
rect 34376 58720 34440 58724
rect 34456 58780 34520 58784
rect 34456 58724 34460 58780
rect 34460 58724 34516 58780
rect 34516 58724 34520 58780
rect 34456 58720 34520 58724
rect 44216 58780 44280 58784
rect 44216 58724 44220 58780
rect 44220 58724 44276 58780
rect 44276 58724 44280 58780
rect 44216 58720 44280 58724
rect 44296 58780 44360 58784
rect 44296 58724 44300 58780
rect 44300 58724 44356 58780
rect 44356 58724 44360 58780
rect 44296 58720 44360 58724
rect 44376 58780 44440 58784
rect 44376 58724 44380 58780
rect 44380 58724 44436 58780
rect 44436 58724 44440 58780
rect 44376 58720 44440 58724
rect 44456 58780 44520 58784
rect 44456 58724 44460 58780
rect 44460 58724 44516 58780
rect 44516 58724 44520 58780
rect 44456 58720 44520 58724
rect 54216 58780 54280 58784
rect 54216 58724 54220 58780
rect 54220 58724 54276 58780
rect 54276 58724 54280 58780
rect 54216 58720 54280 58724
rect 54296 58780 54360 58784
rect 54296 58724 54300 58780
rect 54300 58724 54356 58780
rect 54356 58724 54360 58780
rect 54296 58720 54360 58724
rect 54376 58780 54440 58784
rect 54376 58724 54380 58780
rect 54380 58724 54436 58780
rect 54436 58724 54440 58780
rect 54376 58720 54440 58724
rect 54456 58780 54520 58784
rect 54456 58724 54460 58780
rect 54460 58724 54516 58780
rect 54516 58724 54520 58780
rect 54456 58720 54520 58724
rect 64216 58780 64280 58784
rect 64216 58724 64220 58780
rect 64220 58724 64276 58780
rect 64276 58724 64280 58780
rect 64216 58720 64280 58724
rect 64296 58780 64360 58784
rect 64296 58724 64300 58780
rect 64300 58724 64356 58780
rect 64356 58724 64360 58780
rect 64296 58720 64360 58724
rect 64376 58780 64440 58784
rect 64376 58724 64380 58780
rect 64380 58724 64436 58780
rect 64436 58724 64440 58780
rect 64376 58720 64440 58724
rect 64456 58780 64520 58784
rect 64456 58724 64460 58780
rect 64460 58724 64516 58780
rect 64516 58724 64520 58780
rect 64456 58720 64520 58724
rect 9216 58236 9280 58240
rect 9216 58180 9220 58236
rect 9220 58180 9276 58236
rect 9276 58180 9280 58236
rect 9216 58176 9280 58180
rect 9296 58236 9360 58240
rect 9296 58180 9300 58236
rect 9300 58180 9356 58236
rect 9356 58180 9360 58236
rect 9296 58176 9360 58180
rect 9376 58236 9440 58240
rect 9376 58180 9380 58236
rect 9380 58180 9436 58236
rect 9436 58180 9440 58236
rect 9376 58176 9440 58180
rect 9456 58236 9520 58240
rect 9456 58180 9460 58236
rect 9460 58180 9516 58236
rect 9516 58180 9520 58236
rect 9456 58176 9520 58180
rect 19216 58236 19280 58240
rect 19216 58180 19220 58236
rect 19220 58180 19276 58236
rect 19276 58180 19280 58236
rect 19216 58176 19280 58180
rect 19296 58236 19360 58240
rect 19296 58180 19300 58236
rect 19300 58180 19356 58236
rect 19356 58180 19360 58236
rect 19296 58176 19360 58180
rect 19376 58236 19440 58240
rect 19376 58180 19380 58236
rect 19380 58180 19436 58236
rect 19436 58180 19440 58236
rect 19376 58176 19440 58180
rect 19456 58236 19520 58240
rect 19456 58180 19460 58236
rect 19460 58180 19516 58236
rect 19516 58180 19520 58236
rect 19456 58176 19520 58180
rect 29216 58236 29280 58240
rect 29216 58180 29220 58236
rect 29220 58180 29276 58236
rect 29276 58180 29280 58236
rect 29216 58176 29280 58180
rect 29296 58236 29360 58240
rect 29296 58180 29300 58236
rect 29300 58180 29356 58236
rect 29356 58180 29360 58236
rect 29296 58176 29360 58180
rect 29376 58236 29440 58240
rect 29376 58180 29380 58236
rect 29380 58180 29436 58236
rect 29436 58180 29440 58236
rect 29376 58176 29440 58180
rect 29456 58236 29520 58240
rect 29456 58180 29460 58236
rect 29460 58180 29516 58236
rect 29516 58180 29520 58236
rect 29456 58176 29520 58180
rect 39216 58236 39280 58240
rect 39216 58180 39220 58236
rect 39220 58180 39276 58236
rect 39276 58180 39280 58236
rect 39216 58176 39280 58180
rect 39296 58236 39360 58240
rect 39296 58180 39300 58236
rect 39300 58180 39356 58236
rect 39356 58180 39360 58236
rect 39296 58176 39360 58180
rect 39376 58236 39440 58240
rect 39376 58180 39380 58236
rect 39380 58180 39436 58236
rect 39436 58180 39440 58236
rect 39376 58176 39440 58180
rect 39456 58236 39520 58240
rect 39456 58180 39460 58236
rect 39460 58180 39516 58236
rect 39516 58180 39520 58236
rect 39456 58176 39520 58180
rect 49216 58236 49280 58240
rect 49216 58180 49220 58236
rect 49220 58180 49276 58236
rect 49276 58180 49280 58236
rect 49216 58176 49280 58180
rect 49296 58236 49360 58240
rect 49296 58180 49300 58236
rect 49300 58180 49356 58236
rect 49356 58180 49360 58236
rect 49296 58176 49360 58180
rect 49376 58236 49440 58240
rect 49376 58180 49380 58236
rect 49380 58180 49436 58236
rect 49436 58180 49440 58236
rect 49376 58176 49440 58180
rect 49456 58236 49520 58240
rect 49456 58180 49460 58236
rect 49460 58180 49516 58236
rect 49516 58180 49520 58236
rect 49456 58176 49520 58180
rect 59216 58236 59280 58240
rect 59216 58180 59220 58236
rect 59220 58180 59276 58236
rect 59276 58180 59280 58236
rect 59216 58176 59280 58180
rect 59296 58236 59360 58240
rect 59296 58180 59300 58236
rect 59300 58180 59356 58236
rect 59356 58180 59360 58236
rect 59296 58176 59360 58180
rect 59376 58236 59440 58240
rect 59376 58180 59380 58236
rect 59380 58180 59436 58236
rect 59436 58180 59440 58236
rect 59376 58176 59440 58180
rect 59456 58236 59520 58240
rect 59456 58180 59460 58236
rect 59460 58180 59516 58236
rect 59516 58180 59520 58236
rect 59456 58176 59520 58180
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 14216 57692 14280 57696
rect 14216 57636 14220 57692
rect 14220 57636 14276 57692
rect 14276 57636 14280 57692
rect 14216 57632 14280 57636
rect 14296 57692 14360 57696
rect 14296 57636 14300 57692
rect 14300 57636 14356 57692
rect 14356 57636 14360 57692
rect 14296 57632 14360 57636
rect 14376 57692 14440 57696
rect 14376 57636 14380 57692
rect 14380 57636 14436 57692
rect 14436 57636 14440 57692
rect 14376 57632 14440 57636
rect 14456 57692 14520 57696
rect 14456 57636 14460 57692
rect 14460 57636 14516 57692
rect 14516 57636 14520 57692
rect 14456 57632 14520 57636
rect 24216 57692 24280 57696
rect 24216 57636 24220 57692
rect 24220 57636 24276 57692
rect 24276 57636 24280 57692
rect 24216 57632 24280 57636
rect 24296 57692 24360 57696
rect 24296 57636 24300 57692
rect 24300 57636 24356 57692
rect 24356 57636 24360 57692
rect 24296 57632 24360 57636
rect 24376 57692 24440 57696
rect 24376 57636 24380 57692
rect 24380 57636 24436 57692
rect 24436 57636 24440 57692
rect 24376 57632 24440 57636
rect 24456 57692 24520 57696
rect 24456 57636 24460 57692
rect 24460 57636 24516 57692
rect 24516 57636 24520 57692
rect 24456 57632 24520 57636
rect 34216 57692 34280 57696
rect 34216 57636 34220 57692
rect 34220 57636 34276 57692
rect 34276 57636 34280 57692
rect 34216 57632 34280 57636
rect 34296 57692 34360 57696
rect 34296 57636 34300 57692
rect 34300 57636 34356 57692
rect 34356 57636 34360 57692
rect 34296 57632 34360 57636
rect 34376 57692 34440 57696
rect 34376 57636 34380 57692
rect 34380 57636 34436 57692
rect 34436 57636 34440 57692
rect 34376 57632 34440 57636
rect 34456 57692 34520 57696
rect 34456 57636 34460 57692
rect 34460 57636 34516 57692
rect 34516 57636 34520 57692
rect 34456 57632 34520 57636
rect 44216 57692 44280 57696
rect 44216 57636 44220 57692
rect 44220 57636 44276 57692
rect 44276 57636 44280 57692
rect 44216 57632 44280 57636
rect 44296 57692 44360 57696
rect 44296 57636 44300 57692
rect 44300 57636 44356 57692
rect 44356 57636 44360 57692
rect 44296 57632 44360 57636
rect 44376 57692 44440 57696
rect 44376 57636 44380 57692
rect 44380 57636 44436 57692
rect 44436 57636 44440 57692
rect 44376 57632 44440 57636
rect 44456 57692 44520 57696
rect 44456 57636 44460 57692
rect 44460 57636 44516 57692
rect 44516 57636 44520 57692
rect 44456 57632 44520 57636
rect 54216 57692 54280 57696
rect 54216 57636 54220 57692
rect 54220 57636 54276 57692
rect 54276 57636 54280 57692
rect 54216 57632 54280 57636
rect 54296 57692 54360 57696
rect 54296 57636 54300 57692
rect 54300 57636 54356 57692
rect 54356 57636 54360 57692
rect 54296 57632 54360 57636
rect 54376 57692 54440 57696
rect 54376 57636 54380 57692
rect 54380 57636 54436 57692
rect 54436 57636 54440 57692
rect 54376 57632 54440 57636
rect 54456 57692 54520 57696
rect 54456 57636 54460 57692
rect 54460 57636 54516 57692
rect 54516 57636 54520 57692
rect 54456 57632 54520 57636
rect 64216 57692 64280 57696
rect 64216 57636 64220 57692
rect 64220 57636 64276 57692
rect 64276 57636 64280 57692
rect 64216 57632 64280 57636
rect 64296 57692 64360 57696
rect 64296 57636 64300 57692
rect 64300 57636 64356 57692
rect 64356 57636 64360 57692
rect 64296 57632 64360 57636
rect 64376 57692 64440 57696
rect 64376 57636 64380 57692
rect 64380 57636 64436 57692
rect 64436 57636 64440 57692
rect 64376 57632 64440 57636
rect 64456 57692 64520 57696
rect 64456 57636 64460 57692
rect 64460 57636 64516 57692
rect 64516 57636 64520 57692
rect 64456 57632 64520 57636
rect 9216 57148 9280 57152
rect 9216 57092 9220 57148
rect 9220 57092 9276 57148
rect 9276 57092 9280 57148
rect 9216 57088 9280 57092
rect 9296 57148 9360 57152
rect 9296 57092 9300 57148
rect 9300 57092 9356 57148
rect 9356 57092 9360 57148
rect 9296 57088 9360 57092
rect 9376 57148 9440 57152
rect 9376 57092 9380 57148
rect 9380 57092 9436 57148
rect 9436 57092 9440 57148
rect 9376 57088 9440 57092
rect 9456 57148 9520 57152
rect 9456 57092 9460 57148
rect 9460 57092 9516 57148
rect 9516 57092 9520 57148
rect 9456 57088 9520 57092
rect 19216 57148 19280 57152
rect 19216 57092 19220 57148
rect 19220 57092 19276 57148
rect 19276 57092 19280 57148
rect 19216 57088 19280 57092
rect 19296 57148 19360 57152
rect 19296 57092 19300 57148
rect 19300 57092 19356 57148
rect 19356 57092 19360 57148
rect 19296 57088 19360 57092
rect 19376 57148 19440 57152
rect 19376 57092 19380 57148
rect 19380 57092 19436 57148
rect 19436 57092 19440 57148
rect 19376 57088 19440 57092
rect 19456 57148 19520 57152
rect 19456 57092 19460 57148
rect 19460 57092 19516 57148
rect 19516 57092 19520 57148
rect 19456 57088 19520 57092
rect 29216 57148 29280 57152
rect 29216 57092 29220 57148
rect 29220 57092 29276 57148
rect 29276 57092 29280 57148
rect 29216 57088 29280 57092
rect 29296 57148 29360 57152
rect 29296 57092 29300 57148
rect 29300 57092 29356 57148
rect 29356 57092 29360 57148
rect 29296 57088 29360 57092
rect 29376 57148 29440 57152
rect 29376 57092 29380 57148
rect 29380 57092 29436 57148
rect 29436 57092 29440 57148
rect 29376 57088 29440 57092
rect 29456 57148 29520 57152
rect 29456 57092 29460 57148
rect 29460 57092 29516 57148
rect 29516 57092 29520 57148
rect 29456 57088 29520 57092
rect 39216 57148 39280 57152
rect 39216 57092 39220 57148
rect 39220 57092 39276 57148
rect 39276 57092 39280 57148
rect 39216 57088 39280 57092
rect 39296 57148 39360 57152
rect 39296 57092 39300 57148
rect 39300 57092 39356 57148
rect 39356 57092 39360 57148
rect 39296 57088 39360 57092
rect 39376 57148 39440 57152
rect 39376 57092 39380 57148
rect 39380 57092 39436 57148
rect 39436 57092 39440 57148
rect 39376 57088 39440 57092
rect 39456 57148 39520 57152
rect 39456 57092 39460 57148
rect 39460 57092 39516 57148
rect 39516 57092 39520 57148
rect 39456 57088 39520 57092
rect 49216 57148 49280 57152
rect 49216 57092 49220 57148
rect 49220 57092 49276 57148
rect 49276 57092 49280 57148
rect 49216 57088 49280 57092
rect 49296 57148 49360 57152
rect 49296 57092 49300 57148
rect 49300 57092 49356 57148
rect 49356 57092 49360 57148
rect 49296 57088 49360 57092
rect 49376 57148 49440 57152
rect 49376 57092 49380 57148
rect 49380 57092 49436 57148
rect 49436 57092 49440 57148
rect 49376 57088 49440 57092
rect 49456 57148 49520 57152
rect 49456 57092 49460 57148
rect 49460 57092 49516 57148
rect 49516 57092 49520 57148
rect 49456 57088 49520 57092
rect 59216 57148 59280 57152
rect 59216 57092 59220 57148
rect 59220 57092 59276 57148
rect 59276 57092 59280 57148
rect 59216 57088 59280 57092
rect 59296 57148 59360 57152
rect 59296 57092 59300 57148
rect 59300 57092 59356 57148
rect 59356 57092 59360 57148
rect 59296 57088 59360 57092
rect 59376 57148 59440 57152
rect 59376 57092 59380 57148
rect 59380 57092 59436 57148
rect 59436 57092 59440 57148
rect 59376 57088 59440 57092
rect 59456 57148 59520 57152
rect 59456 57092 59460 57148
rect 59460 57092 59516 57148
rect 59516 57092 59520 57148
rect 59456 57088 59520 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 14216 56604 14280 56608
rect 14216 56548 14220 56604
rect 14220 56548 14276 56604
rect 14276 56548 14280 56604
rect 14216 56544 14280 56548
rect 14296 56604 14360 56608
rect 14296 56548 14300 56604
rect 14300 56548 14356 56604
rect 14356 56548 14360 56604
rect 14296 56544 14360 56548
rect 14376 56604 14440 56608
rect 14376 56548 14380 56604
rect 14380 56548 14436 56604
rect 14436 56548 14440 56604
rect 14376 56544 14440 56548
rect 14456 56604 14520 56608
rect 14456 56548 14460 56604
rect 14460 56548 14516 56604
rect 14516 56548 14520 56604
rect 14456 56544 14520 56548
rect 24216 56604 24280 56608
rect 24216 56548 24220 56604
rect 24220 56548 24276 56604
rect 24276 56548 24280 56604
rect 24216 56544 24280 56548
rect 24296 56604 24360 56608
rect 24296 56548 24300 56604
rect 24300 56548 24356 56604
rect 24356 56548 24360 56604
rect 24296 56544 24360 56548
rect 24376 56604 24440 56608
rect 24376 56548 24380 56604
rect 24380 56548 24436 56604
rect 24436 56548 24440 56604
rect 24376 56544 24440 56548
rect 24456 56604 24520 56608
rect 24456 56548 24460 56604
rect 24460 56548 24516 56604
rect 24516 56548 24520 56604
rect 24456 56544 24520 56548
rect 34216 56604 34280 56608
rect 34216 56548 34220 56604
rect 34220 56548 34276 56604
rect 34276 56548 34280 56604
rect 34216 56544 34280 56548
rect 34296 56604 34360 56608
rect 34296 56548 34300 56604
rect 34300 56548 34356 56604
rect 34356 56548 34360 56604
rect 34296 56544 34360 56548
rect 34376 56604 34440 56608
rect 34376 56548 34380 56604
rect 34380 56548 34436 56604
rect 34436 56548 34440 56604
rect 34376 56544 34440 56548
rect 34456 56604 34520 56608
rect 34456 56548 34460 56604
rect 34460 56548 34516 56604
rect 34516 56548 34520 56604
rect 34456 56544 34520 56548
rect 44216 56604 44280 56608
rect 44216 56548 44220 56604
rect 44220 56548 44276 56604
rect 44276 56548 44280 56604
rect 44216 56544 44280 56548
rect 44296 56604 44360 56608
rect 44296 56548 44300 56604
rect 44300 56548 44356 56604
rect 44356 56548 44360 56604
rect 44296 56544 44360 56548
rect 44376 56604 44440 56608
rect 44376 56548 44380 56604
rect 44380 56548 44436 56604
rect 44436 56548 44440 56604
rect 44376 56544 44440 56548
rect 44456 56604 44520 56608
rect 44456 56548 44460 56604
rect 44460 56548 44516 56604
rect 44516 56548 44520 56604
rect 44456 56544 44520 56548
rect 54216 56604 54280 56608
rect 54216 56548 54220 56604
rect 54220 56548 54276 56604
rect 54276 56548 54280 56604
rect 54216 56544 54280 56548
rect 54296 56604 54360 56608
rect 54296 56548 54300 56604
rect 54300 56548 54356 56604
rect 54356 56548 54360 56604
rect 54296 56544 54360 56548
rect 54376 56604 54440 56608
rect 54376 56548 54380 56604
rect 54380 56548 54436 56604
rect 54436 56548 54440 56604
rect 54376 56544 54440 56548
rect 54456 56604 54520 56608
rect 54456 56548 54460 56604
rect 54460 56548 54516 56604
rect 54516 56548 54520 56604
rect 54456 56544 54520 56548
rect 64216 56604 64280 56608
rect 64216 56548 64220 56604
rect 64220 56548 64276 56604
rect 64276 56548 64280 56604
rect 64216 56544 64280 56548
rect 64296 56604 64360 56608
rect 64296 56548 64300 56604
rect 64300 56548 64356 56604
rect 64356 56548 64360 56604
rect 64296 56544 64360 56548
rect 64376 56604 64440 56608
rect 64376 56548 64380 56604
rect 64380 56548 64436 56604
rect 64436 56548 64440 56604
rect 64376 56544 64440 56548
rect 64456 56604 64520 56608
rect 64456 56548 64460 56604
rect 64460 56548 64516 56604
rect 64516 56548 64520 56604
rect 64456 56544 64520 56548
rect 9216 56060 9280 56064
rect 9216 56004 9220 56060
rect 9220 56004 9276 56060
rect 9276 56004 9280 56060
rect 9216 56000 9280 56004
rect 9296 56060 9360 56064
rect 9296 56004 9300 56060
rect 9300 56004 9356 56060
rect 9356 56004 9360 56060
rect 9296 56000 9360 56004
rect 9376 56060 9440 56064
rect 9376 56004 9380 56060
rect 9380 56004 9436 56060
rect 9436 56004 9440 56060
rect 9376 56000 9440 56004
rect 9456 56060 9520 56064
rect 9456 56004 9460 56060
rect 9460 56004 9516 56060
rect 9516 56004 9520 56060
rect 9456 56000 9520 56004
rect 19216 56060 19280 56064
rect 19216 56004 19220 56060
rect 19220 56004 19276 56060
rect 19276 56004 19280 56060
rect 19216 56000 19280 56004
rect 19296 56060 19360 56064
rect 19296 56004 19300 56060
rect 19300 56004 19356 56060
rect 19356 56004 19360 56060
rect 19296 56000 19360 56004
rect 19376 56060 19440 56064
rect 19376 56004 19380 56060
rect 19380 56004 19436 56060
rect 19436 56004 19440 56060
rect 19376 56000 19440 56004
rect 19456 56060 19520 56064
rect 19456 56004 19460 56060
rect 19460 56004 19516 56060
rect 19516 56004 19520 56060
rect 19456 56000 19520 56004
rect 29216 56060 29280 56064
rect 29216 56004 29220 56060
rect 29220 56004 29276 56060
rect 29276 56004 29280 56060
rect 29216 56000 29280 56004
rect 29296 56060 29360 56064
rect 29296 56004 29300 56060
rect 29300 56004 29356 56060
rect 29356 56004 29360 56060
rect 29296 56000 29360 56004
rect 29376 56060 29440 56064
rect 29376 56004 29380 56060
rect 29380 56004 29436 56060
rect 29436 56004 29440 56060
rect 29376 56000 29440 56004
rect 29456 56060 29520 56064
rect 29456 56004 29460 56060
rect 29460 56004 29516 56060
rect 29516 56004 29520 56060
rect 29456 56000 29520 56004
rect 39216 56060 39280 56064
rect 39216 56004 39220 56060
rect 39220 56004 39276 56060
rect 39276 56004 39280 56060
rect 39216 56000 39280 56004
rect 39296 56060 39360 56064
rect 39296 56004 39300 56060
rect 39300 56004 39356 56060
rect 39356 56004 39360 56060
rect 39296 56000 39360 56004
rect 39376 56060 39440 56064
rect 39376 56004 39380 56060
rect 39380 56004 39436 56060
rect 39436 56004 39440 56060
rect 39376 56000 39440 56004
rect 39456 56060 39520 56064
rect 39456 56004 39460 56060
rect 39460 56004 39516 56060
rect 39516 56004 39520 56060
rect 39456 56000 39520 56004
rect 49216 56060 49280 56064
rect 49216 56004 49220 56060
rect 49220 56004 49276 56060
rect 49276 56004 49280 56060
rect 49216 56000 49280 56004
rect 49296 56060 49360 56064
rect 49296 56004 49300 56060
rect 49300 56004 49356 56060
rect 49356 56004 49360 56060
rect 49296 56000 49360 56004
rect 49376 56060 49440 56064
rect 49376 56004 49380 56060
rect 49380 56004 49436 56060
rect 49436 56004 49440 56060
rect 49376 56000 49440 56004
rect 49456 56060 49520 56064
rect 49456 56004 49460 56060
rect 49460 56004 49516 56060
rect 49516 56004 49520 56060
rect 49456 56000 49520 56004
rect 59216 56060 59280 56064
rect 59216 56004 59220 56060
rect 59220 56004 59276 56060
rect 59276 56004 59280 56060
rect 59216 56000 59280 56004
rect 59296 56060 59360 56064
rect 59296 56004 59300 56060
rect 59300 56004 59356 56060
rect 59356 56004 59360 56060
rect 59296 56000 59360 56004
rect 59376 56060 59440 56064
rect 59376 56004 59380 56060
rect 59380 56004 59436 56060
rect 59436 56004 59440 56060
rect 59376 56000 59440 56004
rect 59456 56060 59520 56064
rect 59456 56004 59460 56060
rect 59460 56004 59516 56060
rect 59516 56004 59520 56060
rect 59456 56000 59520 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 14216 55516 14280 55520
rect 14216 55460 14220 55516
rect 14220 55460 14276 55516
rect 14276 55460 14280 55516
rect 14216 55456 14280 55460
rect 14296 55516 14360 55520
rect 14296 55460 14300 55516
rect 14300 55460 14356 55516
rect 14356 55460 14360 55516
rect 14296 55456 14360 55460
rect 14376 55516 14440 55520
rect 14376 55460 14380 55516
rect 14380 55460 14436 55516
rect 14436 55460 14440 55516
rect 14376 55456 14440 55460
rect 14456 55516 14520 55520
rect 14456 55460 14460 55516
rect 14460 55460 14516 55516
rect 14516 55460 14520 55516
rect 14456 55456 14520 55460
rect 24216 55516 24280 55520
rect 24216 55460 24220 55516
rect 24220 55460 24276 55516
rect 24276 55460 24280 55516
rect 24216 55456 24280 55460
rect 24296 55516 24360 55520
rect 24296 55460 24300 55516
rect 24300 55460 24356 55516
rect 24356 55460 24360 55516
rect 24296 55456 24360 55460
rect 24376 55516 24440 55520
rect 24376 55460 24380 55516
rect 24380 55460 24436 55516
rect 24436 55460 24440 55516
rect 24376 55456 24440 55460
rect 24456 55516 24520 55520
rect 24456 55460 24460 55516
rect 24460 55460 24516 55516
rect 24516 55460 24520 55516
rect 24456 55456 24520 55460
rect 34216 55516 34280 55520
rect 34216 55460 34220 55516
rect 34220 55460 34276 55516
rect 34276 55460 34280 55516
rect 34216 55456 34280 55460
rect 34296 55516 34360 55520
rect 34296 55460 34300 55516
rect 34300 55460 34356 55516
rect 34356 55460 34360 55516
rect 34296 55456 34360 55460
rect 34376 55516 34440 55520
rect 34376 55460 34380 55516
rect 34380 55460 34436 55516
rect 34436 55460 34440 55516
rect 34376 55456 34440 55460
rect 34456 55516 34520 55520
rect 34456 55460 34460 55516
rect 34460 55460 34516 55516
rect 34516 55460 34520 55516
rect 34456 55456 34520 55460
rect 44216 55516 44280 55520
rect 44216 55460 44220 55516
rect 44220 55460 44276 55516
rect 44276 55460 44280 55516
rect 44216 55456 44280 55460
rect 44296 55516 44360 55520
rect 44296 55460 44300 55516
rect 44300 55460 44356 55516
rect 44356 55460 44360 55516
rect 44296 55456 44360 55460
rect 44376 55516 44440 55520
rect 44376 55460 44380 55516
rect 44380 55460 44436 55516
rect 44436 55460 44440 55516
rect 44376 55456 44440 55460
rect 44456 55516 44520 55520
rect 44456 55460 44460 55516
rect 44460 55460 44516 55516
rect 44516 55460 44520 55516
rect 44456 55456 44520 55460
rect 54216 55516 54280 55520
rect 54216 55460 54220 55516
rect 54220 55460 54276 55516
rect 54276 55460 54280 55516
rect 54216 55456 54280 55460
rect 54296 55516 54360 55520
rect 54296 55460 54300 55516
rect 54300 55460 54356 55516
rect 54356 55460 54360 55516
rect 54296 55456 54360 55460
rect 54376 55516 54440 55520
rect 54376 55460 54380 55516
rect 54380 55460 54436 55516
rect 54436 55460 54440 55516
rect 54376 55456 54440 55460
rect 54456 55516 54520 55520
rect 54456 55460 54460 55516
rect 54460 55460 54516 55516
rect 54516 55460 54520 55516
rect 54456 55456 54520 55460
rect 64216 55516 64280 55520
rect 64216 55460 64220 55516
rect 64220 55460 64276 55516
rect 64276 55460 64280 55516
rect 64216 55456 64280 55460
rect 64296 55516 64360 55520
rect 64296 55460 64300 55516
rect 64300 55460 64356 55516
rect 64356 55460 64360 55516
rect 64296 55456 64360 55460
rect 64376 55516 64440 55520
rect 64376 55460 64380 55516
rect 64380 55460 64436 55516
rect 64436 55460 64440 55516
rect 64376 55456 64440 55460
rect 64456 55516 64520 55520
rect 64456 55460 64460 55516
rect 64460 55460 64516 55516
rect 64516 55460 64520 55516
rect 64456 55456 64520 55460
rect 9216 54972 9280 54976
rect 9216 54916 9220 54972
rect 9220 54916 9276 54972
rect 9276 54916 9280 54972
rect 9216 54912 9280 54916
rect 9296 54972 9360 54976
rect 9296 54916 9300 54972
rect 9300 54916 9356 54972
rect 9356 54916 9360 54972
rect 9296 54912 9360 54916
rect 9376 54972 9440 54976
rect 9376 54916 9380 54972
rect 9380 54916 9436 54972
rect 9436 54916 9440 54972
rect 9376 54912 9440 54916
rect 9456 54972 9520 54976
rect 9456 54916 9460 54972
rect 9460 54916 9516 54972
rect 9516 54916 9520 54972
rect 9456 54912 9520 54916
rect 19216 54972 19280 54976
rect 19216 54916 19220 54972
rect 19220 54916 19276 54972
rect 19276 54916 19280 54972
rect 19216 54912 19280 54916
rect 19296 54972 19360 54976
rect 19296 54916 19300 54972
rect 19300 54916 19356 54972
rect 19356 54916 19360 54972
rect 19296 54912 19360 54916
rect 19376 54972 19440 54976
rect 19376 54916 19380 54972
rect 19380 54916 19436 54972
rect 19436 54916 19440 54972
rect 19376 54912 19440 54916
rect 19456 54972 19520 54976
rect 19456 54916 19460 54972
rect 19460 54916 19516 54972
rect 19516 54916 19520 54972
rect 19456 54912 19520 54916
rect 29216 54972 29280 54976
rect 29216 54916 29220 54972
rect 29220 54916 29276 54972
rect 29276 54916 29280 54972
rect 29216 54912 29280 54916
rect 29296 54972 29360 54976
rect 29296 54916 29300 54972
rect 29300 54916 29356 54972
rect 29356 54916 29360 54972
rect 29296 54912 29360 54916
rect 29376 54972 29440 54976
rect 29376 54916 29380 54972
rect 29380 54916 29436 54972
rect 29436 54916 29440 54972
rect 29376 54912 29440 54916
rect 29456 54972 29520 54976
rect 29456 54916 29460 54972
rect 29460 54916 29516 54972
rect 29516 54916 29520 54972
rect 29456 54912 29520 54916
rect 39216 54972 39280 54976
rect 39216 54916 39220 54972
rect 39220 54916 39276 54972
rect 39276 54916 39280 54972
rect 39216 54912 39280 54916
rect 39296 54972 39360 54976
rect 39296 54916 39300 54972
rect 39300 54916 39356 54972
rect 39356 54916 39360 54972
rect 39296 54912 39360 54916
rect 39376 54972 39440 54976
rect 39376 54916 39380 54972
rect 39380 54916 39436 54972
rect 39436 54916 39440 54972
rect 39376 54912 39440 54916
rect 39456 54972 39520 54976
rect 39456 54916 39460 54972
rect 39460 54916 39516 54972
rect 39516 54916 39520 54972
rect 39456 54912 39520 54916
rect 49216 54972 49280 54976
rect 49216 54916 49220 54972
rect 49220 54916 49276 54972
rect 49276 54916 49280 54972
rect 49216 54912 49280 54916
rect 49296 54972 49360 54976
rect 49296 54916 49300 54972
rect 49300 54916 49356 54972
rect 49356 54916 49360 54972
rect 49296 54912 49360 54916
rect 49376 54972 49440 54976
rect 49376 54916 49380 54972
rect 49380 54916 49436 54972
rect 49436 54916 49440 54972
rect 49376 54912 49440 54916
rect 49456 54972 49520 54976
rect 49456 54916 49460 54972
rect 49460 54916 49516 54972
rect 49516 54916 49520 54972
rect 49456 54912 49520 54916
rect 59216 54972 59280 54976
rect 59216 54916 59220 54972
rect 59220 54916 59276 54972
rect 59276 54916 59280 54972
rect 59216 54912 59280 54916
rect 59296 54972 59360 54976
rect 59296 54916 59300 54972
rect 59300 54916 59356 54972
rect 59356 54916 59360 54972
rect 59296 54912 59360 54916
rect 59376 54972 59440 54976
rect 59376 54916 59380 54972
rect 59380 54916 59436 54972
rect 59436 54916 59440 54972
rect 59376 54912 59440 54916
rect 59456 54972 59520 54976
rect 59456 54916 59460 54972
rect 59460 54916 59516 54972
rect 59516 54916 59520 54972
rect 59456 54912 59520 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 14216 54428 14280 54432
rect 14216 54372 14220 54428
rect 14220 54372 14276 54428
rect 14276 54372 14280 54428
rect 14216 54368 14280 54372
rect 14296 54428 14360 54432
rect 14296 54372 14300 54428
rect 14300 54372 14356 54428
rect 14356 54372 14360 54428
rect 14296 54368 14360 54372
rect 14376 54428 14440 54432
rect 14376 54372 14380 54428
rect 14380 54372 14436 54428
rect 14436 54372 14440 54428
rect 14376 54368 14440 54372
rect 14456 54428 14520 54432
rect 14456 54372 14460 54428
rect 14460 54372 14516 54428
rect 14516 54372 14520 54428
rect 14456 54368 14520 54372
rect 24216 54428 24280 54432
rect 24216 54372 24220 54428
rect 24220 54372 24276 54428
rect 24276 54372 24280 54428
rect 24216 54368 24280 54372
rect 24296 54428 24360 54432
rect 24296 54372 24300 54428
rect 24300 54372 24356 54428
rect 24356 54372 24360 54428
rect 24296 54368 24360 54372
rect 24376 54428 24440 54432
rect 24376 54372 24380 54428
rect 24380 54372 24436 54428
rect 24436 54372 24440 54428
rect 24376 54368 24440 54372
rect 24456 54428 24520 54432
rect 24456 54372 24460 54428
rect 24460 54372 24516 54428
rect 24516 54372 24520 54428
rect 24456 54368 24520 54372
rect 34216 54428 34280 54432
rect 34216 54372 34220 54428
rect 34220 54372 34276 54428
rect 34276 54372 34280 54428
rect 34216 54368 34280 54372
rect 34296 54428 34360 54432
rect 34296 54372 34300 54428
rect 34300 54372 34356 54428
rect 34356 54372 34360 54428
rect 34296 54368 34360 54372
rect 34376 54428 34440 54432
rect 34376 54372 34380 54428
rect 34380 54372 34436 54428
rect 34436 54372 34440 54428
rect 34376 54368 34440 54372
rect 34456 54428 34520 54432
rect 34456 54372 34460 54428
rect 34460 54372 34516 54428
rect 34516 54372 34520 54428
rect 34456 54368 34520 54372
rect 44216 54428 44280 54432
rect 44216 54372 44220 54428
rect 44220 54372 44276 54428
rect 44276 54372 44280 54428
rect 44216 54368 44280 54372
rect 44296 54428 44360 54432
rect 44296 54372 44300 54428
rect 44300 54372 44356 54428
rect 44356 54372 44360 54428
rect 44296 54368 44360 54372
rect 44376 54428 44440 54432
rect 44376 54372 44380 54428
rect 44380 54372 44436 54428
rect 44436 54372 44440 54428
rect 44376 54368 44440 54372
rect 44456 54428 44520 54432
rect 44456 54372 44460 54428
rect 44460 54372 44516 54428
rect 44516 54372 44520 54428
rect 44456 54368 44520 54372
rect 54216 54428 54280 54432
rect 54216 54372 54220 54428
rect 54220 54372 54276 54428
rect 54276 54372 54280 54428
rect 54216 54368 54280 54372
rect 54296 54428 54360 54432
rect 54296 54372 54300 54428
rect 54300 54372 54356 54428
rect 54356 54372 54360 54428
rect 54296 54368 54360 54372
rect 54376 54428 54440 54432
rect 54376 54372 54380 54428
rect 54380 54372 54436 54428
rect 54436 54372 54440 54428
rect 54376 54368 54440 54372
rect 54456 54428 54520 54432
rect 54456 54372 54460 54428
rect 54460 54372 54516 54428
rect 54516 54372 54520 54428
rect 54456 54368 54520 54372
rect 64216 54428 64280 54432
rect 64216 54372 64220 54428
rect 64220 54372 64276 54428
rect 64276 54372 64280 54428
rect 64216 54368 64280 54372
rect 64296 54428 64360 54432
rect 64296 54372 64300 54428
rect 64300 54372 64356 54428
rect 64356 54372 64360 54428
rect 64296 54368 64360 54372
rect 64376 54428 64440 54432
rect 64376 54372 64380 54428
rect 64380 54372 64436 54428
rect 64436 54372 64440 54428
rect 64376 54368 64440 54372
rect 64456 54428 64520 54432
rect 64456 54372 64460 54428
rect 64460 54372 64516 54428
rect 64516 54372 64520 54428
rect 64456 54368 64520 54372
rect 9216 53884 9280 53888
rect 9216 53828 9220 53884
rect 9220 53828 9276 53884
rect 9276 53828 9280 53884
rect 9216 53824 9280 53828
rect 9296 53884 9360 53888
rect 9296 53828 9300 53884
rect 9300 53828 9356 53884
rect 9356 53828 9360 53884
rect 9296 53824 9360 53828
rect 9376 53884 9440 53888
rect 9376 53828 9380 53884
rect 9380 53828 9436 53884
rect 9436 53828 9440 53884
rect 9376 53824 9440 53828
rect 9456 53884 9520 53888
rect 9456 53828 9460 53884
rect 9460 53828 9516 53884
rect 9516 53828 9520 53884
rect 9456 53824 9520 53828
rect 19216 53884 19280 53888
rect 19216 53828 19220 53884
rect 19220 53828 19276 53884
rect 19276 53828 19280 53884
rect 19216 53824 19280 53828
rect 19296 53884 19360 53888
rect 19296 53828 19300 53884
rect 19300 53828 19356 53884
rect 19356 53828 19360 53884
rect 19296 53824 19360 53828
rect 19376 53884 19440 53888
rect 19376 53828 19380 53884
rect 19380 53828 19436 53884
rect 19436 53828 19440 53884
rect 19376 53824 19440 53828
rect 19456 53884 19520 53888
rect 19456 53828 19460 53884
rect 19460 53828 19516 53884
rect 19516 53828 19520 53884
rect 19456 53824 19520 53828
rect 29216 53884 29280 53888
rect 29216 53828 29220 53884
rect 29220 53828 29276 53884
rect 29276 53828 29280 53884
rect 29216 53824 29280 53828
rect 29296 53884 29360 53888
rect 29296 53828 29300 53884
rect 29300 53828 29356 53884
rect 29356 53828 29360 53884
rect 29296 53824 29360 53828
rect 29376 53884 29440 53888
rect 29376 53828 29380 53884
rect 29380 53828 29436 53884
rect 29436 53828 29440 53884
rect 29376 53824 29440 53828
rect 29456 53884 29520 53888
rect 29456 53828 29460 53884
rect 29460 53828 29516 53884
rect 29516 53828 29520 53884
rect 29456 53824 29520 53828
rect 39216 53884 39280 53888
rect 39216 53828 39220 53884
rect 39220 53828 39276 53884
rect 39276 53828 39280 53884
rect 39216 53824 39280 53828
rect 39296 53884 39360 53888
rect 39296 53828 39300 53884
rect 39300 53828 39356 53884
rect 39356 53828 39360 53884
rect 39296 53824 39360 53828
rect 39376 53884 39440 53888
rect 39376 53828 39380 53884
rect 39380 53828 39436 53884
rect 39436 53828 39440 53884
rect 39376 53824 39440 53828
rect 39456 53884 39520 53888
rect 39456 53828 39460 53884
rect 39460 53828 39516 53884
rect 39516 53828 39520 53884
rect 39456 53824 39520 53828
rect 49216 53884 49280 53888
rect 49216 53828 49220 53884
rect 49220 53828 49276 53884
rect 49276 53828 49280 53884
rect 49216 53824 49280 53828
rect 49296 53884 49360 53888
rect 49296 53828 49300 53884
rect 49300 53828 49356 53884
rect 49356 53828 49360 53884
rect 49296 53824 49360 53828
rect 49376 53884 49440 53888
rect 49376 53828 49380 53884
rect 49380 53828 49436 53884
rect 49436 53828 49440 53884
rect 49376 53824 49440 53828
rect 49456 53884 49520 53888
rect 49456 53828 49460 53884
rect 49460 53828 49516 53884
rect 49516 53828 49520 53884
rect 49456 53824 49520 53828
rect 59216 53884 59280 53888
rect 59216 53828 59220 53884
rect 59220 53828 59276 53884
rect 59276 53828 59280 53884
rect 59216 53824 59280 53828
rect 59296 53884 59360 53888
rect 59296 53828 59300 53884
rect 59300 53828 59356 53884
rect 59356 53828 59360 53884
rect 59296 53824 59360 53828
rect 59376 53884 59440 53888
rect 59376 53828 59380 53884
rect 59380 53828 59436 53884
rect 59436 53828 59440 53884
rect 59376 53824 59440 53828
rect 59456 53884 59520 53888
rect 59456 53828 59460 53884
rect 59460 53828 59516 53884
rect 59516 53828 59520 53884
rect 59456 53824 59520 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 14216 53340 14280 53344
rect 14216 53284 14220 53340
rect 14220 53284 14276 53340
rect 14276 53284 14280 53340
rect 14216 53280 14280 53284
rect 14296 53340 14360 53344
rect 14296 53284 14300 53340
rect 14300 53284 14356 53340
rect 14356 53284 14360 53340
rect 14296 53280 14360 53284
rect 14376 53340 14440 53344
rect 14376 53284 14380 53340
rect 14380 53284 14436 53340
rect 14436 53284 14440 53340
rect 14376 53280 14440 53284
rect 14456 53340 14520 53344
rect 14456 53284 14460 53340
rect 14460 53284 14516 53340
rect 14516 53284 14520 53340
rect 14456 53280 14520 53284
rect 24216 53340 24280 53344
rect 24216 53284 24220 53340
rect 24220 53284 24276 53340
rect 24276 53284 24280 53340
rect 24216 53280 24280 53284
rect 24296 53340 24360 53344
rect 24296 53284 24300 53340
rect 24300 53284 24356 53340
rect 24356 53284 24360 53340
rect 24296 53280 24360 53284
rect 24376 53340 24440 53344
rect 24376 53284 24380 53340
rect 24380 53284 24436 53340
rect 24436 53284 24440 53340
rect 24376 53280 24440 53284
rect 24456 53340 24520 53344
rect 24456 53284 24460 53340
rect 24460 53284 24516 53340
rect 24516 53284 24520 53340
rect 24456 53280 24520 53284
rect 34216 53340 34280 53344
rect 34216 53284 34220 53340
rect 34220 53284 34276 53340
rect 34276 53284 34280 53340
rect 34216 53280 34280 53284
rect 34296 53340 34360 53344
rect 34296 53284 34300 53340
rect 34300 53284 34356 53340
rect 34356 53284 34360 53340
rect 34296 53280 34360 53284
rect 34376 53340 34440 53344
rect 34376 53284 34380 53340
rect 34380 53284 34436 53340
rect 34436 53284 34440 53340
rect 34376 53280 34440 53284
rect 34456 53340 34520 53344
rect 34456 53284 34460 53340
rect 34460 53284 34516 53340
rect 34516 53284 34520 53340
rect 34456 53280 34520 53284
rect 44216 53340 44280 53344
rect 44216 53284 44220 53340
rect 44220 53284 44276 53340
rect 44276 53284 44280 53340
rect 44216 53280 44280 53284
rect 44296 53340 44360 53344
rect 44296 53284 44300 53340
rect 44300 53284 44356 53340
rect 44356 53284 44360 53340
rect 44296 53280 44360 53284
rect 44376 53340 44440 53344
rect 44376 53284 44380 53340
rect 44380 53284 44436 53340
rect 44436 53284 44440 53340
rect 44376 53280 44440 53284
rect 44456 53340 44520 53344
rect 44456 53284 44460 53340
rect 44460 53284 44516 53340
rect 44516 53284 44520 53340
rect 44456 53280 44520 53284
rect 54216 53340 54280 53344
rect 54216 53284 54220 53340
rect 54220 53284 54276 53340
rect 54276 53284 54280 53340
rect 54216 53280 54280 53284
rect 54296 53340 54360 53344
rect 54296 53284 54300 53340
rect 54300 53284 54356 53340
rect 54356 53284 54360 53340
rect 54296 53280 54360 53284
rect 54376 53340 54440 53344
rect 54376 53284 54380 53340
rect 54380 53284 54436 53340
rect 54436 53284 54440 53340
rect 54376 53280 54440 53284
rect 54456 53340 54520 53344
rect 54456 53284 54460 53340
rect 54460 53284 54516 53340
rect 54516 53284 54520 53340
rect 54456 53280 54520 53284
rect 64216 53340 64280 53344
rect 64216 53284 64220 53340
rect 64220 53284 64276 53340
rect 64276 53284 64280 53340
rect 64216 53280 64280 53284
rect 64296 53340 64360 53344
rect 64296 53284 64300 53340
rect 64300 53284 64356 53340
rect 64356 53284 64360 53340
rect 64296 53280 64360 53284
rect 64376 53340 64440 53344
rect 64376 53284 64380 53340
rect 64380 53284 64436 53340
rect 64436 53284 64440 53340
rect 64376 53280 64440 53284
rect 64456 53340 64520 53344
rect 64456 53284 64460 53340
rect 64460 53284 64516 53340
rect 64516 53284 64520 53340
rect 64456 53280 64520 53284
rect 9216 52796 9280 52800
rect 9216 52740 9220 52796
rect 9220 52740 9276 52796
rect 9276 52740 9280 52796
rect 9216 52736 9280 52740
rect 9296 52796 9360 52800
rect 9296 52740 9300 52796
rect 9300 52740 9356 52796
rect 9356 52740 9360 52796
rect 9296 52736 9360 52740
rect 9376 52796 9440 52800
rect 9376 52740 9380 52796
rect 9380 52740 9436 52796
rect 9436 52740 9440 52796
rect 9376 52736 9440 52740
rect 9456 52796 9520 52800
rect 9456 52740 9460 52796
rect 9460 52740 9516 52796
rect 9516 52740 9520 52796
rect 9456 52736 9520 52740
rect 19216 52796 19280 52800
rect 19216 52740 19220 52796
rect 19220 52740 19276 52796
rect 19276 52740 19280 52796
rect 19216 52736 19280 52740
rect 19296 52796 19360 52800
rect 19296 52740 19300 52796
rect 19300 52740 19356 52796
rect 19356 52740 19360 52796
rect 19296 52736 19360 52740
rect 19376 52796 19440 52800
rect 19376 52740 19380 52796
rect 19380 52740 19436 52796
rect 19436 52740 19440 52796
rect 19376 52736 19440 52740
rect 19456 52796 19520 52800
rect 19456 52740 19460 52796
rect 19460 52740 19516 52796
rect 19516 52740 19520 52796
rect 19456 52736 19520 52740
rect 29216 52796 29280 52800
rect 29216 52740 29220 52796
rect 29220 52740 29276 52796
rect 29276 52740 29280 52796
rect 29216 52736 29280 52740
rect 29296 52796 29360 52800
rect 29296 52740 29300 52796
rect 29300 52740 29356 52796
rect 29356 52740 29360 52796
rect 29296 52736 29360 52740
rect 29376 52796 29440 52800
rect 29376 52740 29380 52796
rect 29380 52740 29436 52796
rect 29436 52740 29440 52796
rect 29376 52736 29440 52740
rect 29456 52796 29520 52800
rect 29456 52740 29460 52796
rect 29460 52740 29516 52796
rect 29516 52740 29520 52796
rect 29456 52736 29520 52740
rect 39216 52796 39280 52800
rect 39216 52740 39220 52796
rect 39220 52740 39276 52796
rect 39276 52740 39280 52796
rect 39216 52736 39280 52740
rect 39296 52796 39360 52800
rect 39296 52740 39300 52796
rect 39300 52740 39356 52796
rect 39356 52740 39360 52796
rect 39296 52736 39360 52740
rect 39376 52796 39440 52800
rect 39376 52740 39380 52796
rect 39380 52740 39436 52796
rect 39436 52740 39440 52796
rect 39376 52736 39440 52740
rect 39456 52796 39520 52800
rect 39456 52740 39460 52796
rect 39460 52740 39516 52796
rect 39516 52740 39520 52796
rect 39456 52736 39520 52740
rect 49216 52796 49280 52800
rect 49216 52740 49220 52796
rect 49220 52740 49276 52796
rect 49276 52740 49280 52796
rect 49216 52736 49280 52740
rect 49296 52796 49360 52800
rect 49296 52740 49300 52796
rect 49300 52740 49356 52796
rect 49356 52740 49360 52796
rect 49296 52736 49360 52740
rect 49376 52796 49440 52800
rect 49376 52740 49380 52796
rect 49380 52740 49436 52796
rect 49436 52740 49440 52796
rect 49376 52736 49440 52740
rect 49456 52796 49520 52800
rect 49456 52740 49460 52796
rect 49460 52740 49516 52796
rect 49516 52740 49520 52796
rect 49456 52736 49520 52740
rect 59216 52796 59280 52800
rect 59216 52740 59220 52796
rect 59220 52740 59276 52796
rect 59276 52740 59280 52796
rect 59216 52736 59280 52740
rect 59296 52796 59360 52800
rect 59296 52740 59300 52796
rect 59300 52740 59356 52796
rect 59356 52740 59360 52796
rect 59296 52736 59360 52740
rect 59376 52796 59440 52800
rect 59376 52740 59380 52796
rect 59380 52740 59436 52796
rect 59436 52740 59440 52796
rect 59376 52736 59440 52740
rect 59456 52796 59520 52800
rect 59456 52740 59460 52796
rect 59460 52740 59516 52796
rect 59516 52740 59520 52796
rect 59456 52736 59520 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 14216 52252 14280 52256
rect 14216 52196 14220 52252
rect 14220 52196 14276 52252
rect 14276 52196 14280 52252
rect 14216 52192 14280 52196
rect 14296 52252 14360 52256
rect 14296 52196 14300 52252
rect 14300 52196 14356 52252
rect 14356 52196 14360 52252
rect 14296 52192 14360 52196
rect 14376 52252 14440 52256
rect 14376 52196 14380 52252
rect 14380 52196 14436 52252
rect 14436 52196 14440 52252
rect 14376 52192 14440 52196
rect 14456 52252 14520 52256
rect 14456 52196 14460 52252
rect 14460 52196 14516 52252
rect 14516 52196 14520 52252
rect 14456 52192 14520 52196
rect 24216 52252 24280 52256
rect 24216 52196 24220 52252
rect 24220 52196 24276 52252
rect 24276 52196 24280 52252
rect 24216 52192 24280 52196
rect 24296 52252 24360 52256
rect 24296 52196 24300 52252
rect 24300 52196 24356 52252
rect 24356 52196 24360 52252
rect 24296 52192 24360 52196
rect 24376 52252 24440 52256
rect 24376 52196 24380 52252
rect 24380 52196 24436 52252
rect 24436 52196 24440 52252
rect 24376 52192 24440 52196
rect 24456 52252 24520 52256
rect 24456 52196 24460 52252
rect 24460 52196 24516 52252
rect 24516 52196 24520 52252
rect 24456 52192 24520 52196
rect 34216 52252 34280 52256
rect 34216 52196 34220 52252
rect 34220 52196 34276 52252
rect 34276 52196 34280 52252
rect 34216 52192 34280 52196
rect 34296 52252 34360 52256
rect 34296 52196 34300 52252
rect 34300 52196 34356 52252
rect 34356 52196 34360 52252
rect 34296 52192 34360 52196
rect 34376 52252 34440 52256
rect 34376 52196 34380 52252
rect 34380 52196 34436 52252
rect 34436 52196 34440 52252
rect 34376 52192 34440 52196
rect 34456 52252 34520 52256
rect 34456 52196 34460 52252
rect 34460 52196 34516 52252
rect 34516 52196 34520 52252
rect 34456 52192 34520 52196
rect 44216 52252 44280 52256
rect 44216 52196 44220 52252
rect 44220 52196 44276 52252
rect 44276 52196 44280 52252
rect 44216 52192 44280 52196
rect 44296 52252 44360 52256
rect 44296 52196 44300 52252
rect 44300 52196 44356 52252
rect 44356 52196 44360 52252
rect 44296 52192 44360 52196
rect 44376 52252 44440 52256
rect 44376 52196 44380 52252
rect 44380 52196 44436 52252
rect 44436 52196 44440 52252
rect 44376 52192 44440 52196
rect 44456 52252 44520 52256
rect 44456 52196 44460 52252
rect 44460 52196 44516 52252
rect 44516 52196 44520 52252
rect 44456 52192 44520 52196
rect 54216 52252 54280 52256
rect 54216 52196 54220 52252
rect 54220 52196 54276 52252
rect 54276 52196 54280 52252
rect 54216 52192 54280 52196
rect 54296 52252 54360 52256
rect 54296 52196 54300 52252
rect 54300 52196 54356 52252
rect 54356 52196 54360 52252
rect 54296 52192 54360 52196
rect 54376 52252 54440 52256
rect 54376 52196 54380 52252
rect 54380 52196 54436 52252
rect 54436 52196 54440 52252
rect 54376 52192 54440 52196
rect 54456 52252 54520 52256
rect 54456 52196 54460 52252
rect 54460 52196 54516 52252
rect 54516 52196 54520 52252
rect 54456 52192 54520 52196
rect 64216 52252 64280 52256
rect 64216 52196 64220 52252
rect 64220 52196 64276 52252
rect 64276 52196 64280 52252
rect 64216 52192 64280 52196
rect 64296 52252 64360 52256
rect 64296 52196 64300 52252
rect 64300 52196 64356 52252
rect 64356 52196 64360 52252
rect 64296 52192 64360 52196
rect 64376 52252 64440 52256
rect 64376 52196 64380 52252
rect 64380 52196 64436 52252
rect 64436 52196 64440 52252
rect 64376 52192 64440 52196
rect 64456 52252 64520 52256
rect 64456 52196 64460 52252
rect 64460 52196 64516 52252
rect 64516 52196 64520 52252
rect 64456 52192 64520 52196
rect 9216 51708 9280 51712
rect 9216 51652 9220 51708
rect 9220 51652 9276 51708
rect 9276 51652 9280 51708
rect 9216 51648 9280 51652
rect 9296 51708 9360 51712
rect 9296 51652 9300 51708
rect 9300 51652 9356 51708
rect 9356 51652 9360 51708
rect 9296 51648 9360 51652
rect 9376 51708 9440 51712
rect 9376 51652 9380 51708
rect 9380 51652 9436 51708
rect 9436 51652 9440 51708
rect 9376 51648 9440 51652
rect 9456 51708 9520 51712
rect 9456 51652 9460 51708
rect 9460 51652 9516 51708
rect 9516 51652 9520 51708
rect 9456 51648 9520 51652
rect 19216 51708 19280 51712
rect 19216 51652 19220 51708
rect 19220 51652 19276 51708
rect 19276 51652 19280 51708
rect 19216 51648 19280 51652
rect 19296 51708 19360 51712
rect 19296 51652 19300 51708
rect 19300 51652 19356 51708
rect 19356 51652 19360 51708
rect 19296 51648 19360 51652
rect 19376 51708 19440 51712
rect 19376 51652 19380 51708
rect 19380 51652 19436 51708
rect 19436 51652 19440 51708
rect 19376 51648 19440 51652
rect 19456 51708 19520 51712
rect 19456 51652 19460 51708
rect 19460 51652 19516 51708
rect 19516 51652 19520 51708
rect 19456 51648 19520 51652
rect 29216 51708 29280 51712
rect 29216 51652 29220 51708
rect 29220 51652 29276 51708
rect 29276 51652 29280 51708
rect 29216 51648 29280 51652
rect 29296 51708 29360 51712
rect 29296 51652 29300 51708
rect 29300 51652 29356 51708
rect 29356 51652 29360 51708
rect 29296 51648 29360 51652
rect 29376 51708 29440 51712
rect 29376 51652 29380 51708
rect 29380 51652 29436 51708
rect 29436 51652 29440 51708
rect 29376 51648 29440 51652
rect 29456 51708 29520 51712
rect 29456 51652 29460 51708
rect 29460 51652 29516 51708
rect 29516 51652 29520 51708
rect 29456 51648 29520 51652
rect 39216 51708 39280 51712
rect 39216 51652 39220 51708
rect 39220 51652 39276 51708
rect 39276 51652 39280 51708
rect 39216 51648 39280 51652
rect 39296 51708 39360 51712
rect 39296 51652 39300 51708
rect 39300 51652 39356 51708
rect 39356 51652 39360 51708
rect 39296 51648 39360 51652
rect 39376 51708 39440 51712
rect 39376 51652 39380 51708
rect 39380 51652 39436 51708
rect 39436 51652 39440 51708
rect 39376 51648 39440 51652
rect 39456 51708 39520 51712
rect 39456 51652 39460 51708
rect 39460 51652 39516 51708
rect 39516 51652 39520 51708
rect 39456 51648 39520 51652
rect 49216 51708 49280 51712
rect 49216 51652 49220 51708
rect 49220 51652 49276 51708
rect 49276 51652 49280 51708
rect 49216 51648 49280 51652
rect 49296 51708 49360 51712
rect 49296 51652 49300 51708
rect 49300 51652 49356 51708
rect 49356 51652 49360 51708
rect 49296 51648 49360 51652
rect 49376 51708 49440 51712
rect 49376 51652 49380 51708
rect 49380 51652 49436 51708
rect 49436 51652 49440 51708
rect 49376 51648 49440 51652
rect 49456 51708 49520 51712
rect 49456 51652 49460 51708
rect 49460 51652 49516 51708
rect 49516 51652 49520 51708
rect 49456 51648 49520 51652
rect 59216 51708 59280 51712
rect 59216 51652 59220 51708
rect 59220 51652 59276 51708
rect 59276 51652 59280 51708
rect 59216 51648 59280 51652
rect 59296 51708 59360 51712
rect 59296 51652 59300 51708
rect 59300 51652 59356 51708
rect 59356 51652 59360 51708
rect 59296 51648 59360 51652
rect 59376 51708 59440 51712
rect 59376 51652 59380 51708
rect 59380 51652 59436 51708
rect 59436 51652 59440 51708
rect 59376 51648 59440 51652
rect 59456 51708 59520 51712
rect 59456 51652 59460 51708
rect 59460 51652 59516 51708
rect 59516 51652 59520 51708
rect 59456 51648 59520 51652
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 14216 51164 14280 51168
rect 14216 51108 14220 51164
rect 14220 51108 14276 51164
rect 14276 51108 14280 51164
rect 14216 51104 14280 51108
rect 14296 51164 14360 51168
rect 14296 51108 14300 51164
rect 14300 51108 14356 51164
rect 14356 51108 14360 51164
rect 14296 51104 14360 51108
rect 14376 51164 14440 51168
rect 14376 51108 14380 51164
rect 14380 51108 14436 51164
rect 14436 51108 14440 51164
rect 14376 51104 14440 51108
rect 14456 51164 14520 51168
rect 14456 51108 14460 51164
rect 14460 51108 14516 51164
rect 14516 51108 14520 51164
rect 14456 51104 14520 51108
rect 24216 51164 24280 51168
rect 24216 51108 24220 51164
rect 24220 51108 24276 51164
rect 24276 51108 24280 51164
rect 24216 51104 24280 51108
rect 24296 51164 24360 51168
rect 24296 51108 24300 51164
rect 24300 51108 24356 51164
rect 24356 51108 24360 51164
rect 24296 51104 24360 51108
rect 24376 51164 24440 51168
rect 24376 51108 24380 51164
rect 24380 51108 24436 51164
rect 24436 51108 24440 51164
rect 24376 51104 24440 51108
rect 24456 51164 24520 51168
rect 24456 51108 24460 51164
rect 24460 51108 24516 51164
rect 24516 51108 24520 51164
rect 24456 51104 24520 51108
rect 34216 51164 34280 51168
rect 34216 51108 34220 51164
rect 34220 51108 34276 51164
rect 34276 51108 34280 51164
rect 34216 51104 34280 51108
rect 34296 51164 34360 51168
rect 34296 51108 34300 51164
rect 34300 51108 34356 51164
rect 34356 51108 34360 51164
rect 34296 51104 34360 51108
rect 34376 51164 34440 51168
rect 34376 51108 34380 51164
rect 34380 51108 34436 51164
rect 34436 51108 34440 51164
rect 34376 51104 34440 51108
rect 34456 51164 34520 51168
rect 34456 51108 34460 51164
rect 34460 51108 34516 51164
rect 34516 51108 34520 51164
rect 34456 51104 34520 51108
rect 44216 51164 44280 51168
rect 44216 51108 44220 51164
rect 44220 51108 44276 51164
rect 44276 51108 44280 51164
rect 44216 51104 44280 51108
rect 44296 51164 44360 51168
rect 44296 51108 44300 51164
rect 44300 51108 44356 51164
rect 44356 51108 44360 51164
rect 44296 51104 44360 51108
rect 44376 51164 44440 51168
rect 44376 51108 44380 51164
rect 44380 51108 44436 51164
rect 44436 51108 44440 51164
rect 44376 51104 44440 51108
rect 44456 51164 44520 51168
rect 44456 51108 44460 51164
rect 44460 51108 44516 51164
rect 44516 51108 44520 51164
rect 44456 51104 44520 51108
rect 54216 51164 54280 51168
rect 54216 51108 54220 51164
rect 54220 51108 54276 51164
rect 54276 51108 54280 51164
rect 54216 51104 54280 51108
rect 54296 51164 54360 51168
rect 54296 51108 54300 51164
rect 54300 51108 54356 51164
rect 54356 51108 54360 51164
rect 54296 51104 54360 51108
rect 54376 51164 54440 51168
rect 54376 51108 54380 51164
rect 54380 51108 54436 51164
rect 54436 51108 54440 51164
rect 54376 51104 54440 51108
rect 54456 51164 54520 51168
rect 54456 51108 54460 51164
rect 54460 51108 54516 51164
rect 54516 51108 54520 51164
rect 54456 51104 54520 51108
rect 64216 51164 64280 51168
rect 64216 51108 64220 51164
rect 64220 51108 64276 51164
rect 64276 51108 64280 51164
rect 64216 51104 64280 51108
rect 64296 51164 64360 51168
rect 64296 51108 64300 51164
rect 64300 51108 64356 51164
rect 64356 51108 64360 51164
rect 64296 51104 64360 51108
rect 64376 51164 64440 51168
rect 64376 51108 64380 51164
rect 64380 51108 64436 51164
rect 64436 51108 64440 51164
rect 64376 51104 64440 51108
rect 64456 51164 64520 51168
rect 64456 51108 64460 51164
rect 64460 51108 64516 51164
rect 64516 51108 64520 51164
rect 64456 51104 64520 51108
rect 9216 50620 9280 50624
rect 9216 50564 9220 50620
rect 9220 50564 9276 50620
rect 9276 50564 9280 50620
rect 9216 50560 9280 50564
rect 9296 50620 9360 50624
rect 9296 50564 9300 50620
rect 9300 50564 9356 50620
rect 9356 50564 9360 50620
rect 9296 50560 9360 50564
rect 9376 50620 9440 50624
rect 9376 50564 9380 50620
rect 9380 50564 9436 50620
rect 9436 50564 9440 50620
rect 9376 50560 9440 50564
rect 9456 50620 9520 50624
rect 9456 50564 9460 50620
rect 9460 50564 9516 50620
rect 9516 50564 9520 50620
rect 9456 50560 9520 50564
rect 19216 50620 19280 50624
rect 19216 50564 19220 50620
rect 19220 50564 19276 50620
rect 19276 50564 19280 50620
rect 19216 50560 19280 50564
rect 19296 50620 19360 50624
rect 19296 50564 19300 50620
rect 19300 50564 19356 50620
rect 19356 50564 19360 50620
rect 19296 50560 19360 50564
rect 19376 50620 19440 50624
rect 19376 50564 19380 50620
rect 19380 50564 19436 50620
rect 19436 50564 19440 50620
rect 19376 50560 19440 50564
rect 19456 50620 19520 50624
rect 19456 50564 19460 50620
rect 19460 50564 19516 50620
rect 19516 50564 19520 50620
rect 19456 50560 19520 50564
rect 29216 50620 29280 50624
rect 29216 50564 29220 50620
rect 29220 50564 29276 50620
rect 29276 50564 29280 50620
rect 29216 50560 29280 50564
rect 29296 50620 29360 50624
rect 29296 50564 29300 50620
rect 29300 50564 29356 50620
rect 29356 50564 29360 50620
rect 29296 50560 29360 50564
rect 29376 50620 29440 50624
rect 29376 50564 29380 50620
rect 29380 50564 29436 50620
rect 29436 50564 29440 50620
rect 29376 50560 29440 50564
rect 29456 50620 29520 50624
rect 29456 50564 29460 50620
rect 29460 50564 29516 50620
rect 29516 50564 29520 50620
rect 29456 50560 29520 50564
rect 39216 50620 39280 50624
rect 39216 50564 39220 50620
rect 39220 50564 39276 50620
rect 39276 50564 39280 50620
rect 39216 50560 39280 50564
rect 39296 50620 39360 50624
rect 39296 50564 39300 50620
rect 39300 50564 39356 50620
rect 39356 50564 39360 50620
rect 39296 50560 39360 50564
rect 39376 50620 39440 50624
rect 39376 50564 39380 50620
rect 39380 50564 39436 50620
rect 39436 50564 39440 50620
rect 39376 50560 39440 50564
rect 39456 50620 39520 50624
rect 39456 50564 39460 50620
rect 39460 50564 39516 50620
rect 39516 50564 39520 50620
rect 39456 50560 39520 50564
rect 49216 50620 49280 50624
rect 49216 50564 49220 50620
rect 49220 50564 49276 50620
rect 49276 50564 49280 50620
rect 49216 50560 49280 50564
rect 49296 50620 49360 50624
rect 49296 50564 49300 50620
rect 49300 50564 49356 50620
rect 49356 50564 49360 50620
rect 49296 50560 49360 50564
rect 49376 50620 49440 50624
rect 49376 50564 49380 50620
rect 49380 50564 49436 50620
rect 49436 50564 49440 50620
rect 49376 50560 49440 50564
rect 49456 50620 49520 50624
rect 49456 50564 49460 50620
rect 49460 50564 49516 50620
rect 49516 50564 49520 50620
rect 49456 50560 49520 50564
rect 59216 50620 59280 50624
rect 59216 50564 59220 50620
rect 59220 50564 59276 50620
rect 59276 50564 59280 50620
rect 59216 50560 59280 50564
rect 59296 50620 59360 50624
rect 59296 50564 59300 50620
rect 59300 50564 59356 50620
rect 59356 50564 59360 50620
rect 59296 50560 59360 50564
rect 59376 50620 59440 50624
rect 59376 50564 59380 50620
rect 59380 50564 59436 50620
rect 59436 50564 59440 50620
rect 59376 50560 59440 50564
rect 59456 50620 59520 50624
rect 59456 50564 59460 50620
rect 59460 50564 59516 50620
rect 59516 50564 59520 50620
rect 59456 50560 59520 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 14216 50076 14280 50080
rect 14216 50020 14220 50076
rect 14220 50020 14276 50076
rect 14276 50020 14280 50076
rect 14216 50016 14280 50020
rect 14296 50076 14360 50080
rect 14296 50020 14300 50076
rect 14300 50020 14356 50076
rect 14356 50020 14360 50076
rect 14296 50016 14360 50020
rect 14376 50076 14440 50080
rect 14376 50020 14380 50076
rect 14380 50020 14436 50076
rect 14436 50020 14440 50076
rect 14376 50016 14440 50020
rect 14456 50076 14520 50080
rect 14456 50020 14460 50076
rect 14460 50020 14516 50076
rect 14516 50020 14520 50076
rect 14456 50016 14520 50020
rect 24216 50076 24280 50080
rect 24216 50020 24220 50076
rect 24220 50020 24276 50076
rect 24276 50020 24280 50076
rect 24216 50016 24280 50020
rect 24296 50076 24360 50080
rect 24296 50020 24300 50076
rect 24300 50020 24356 50076
rect 24356 50020 24360 50076
rect 24296 50016 24360 50020
rect 24376 50076 24440 50080
rect 24376 50020 24380 50076
rect 24380 50020 24436 50076
rect 24436 50020 24440 50076
rect 24376 50016 24440 50020
rect 24456 50076 24520 50080
rect 24456 50020 24460 50076
rect 24460 50020 24516 50076
rect 24516 50020 24520 50076
rect 24456 50016 24520 50020
rect 34216 50076 34280 50080
rect 34216 50020 34220 50076
rect 34220 50020 34276 50076
rect 34276 50020 34280 50076
rect 34216 50016 34280 50020
rect 34296 50076 34360 50080
rect 34296 50020 34300 50076
rect 34300 50020 34356 50076
rect 34356 50020 34360 50076
rect 34296 50016 34360 50020
rect 34376 50076 34440 50080
rect 34376 50020 34380 50076
rect 34380 50020 34436 50076
rect 34436 50020 34440 50076
rect 34376 50016 34440 50020
rect 34456 50076 34520 50080
rect 34456 50020 34460 50076
rect 34460 50020 34516 50076
rect 34516 50020 34520 50076
rect 34456 50016 34520 50020
rect 44216 50076 44280 50080
rect 44216 50020 44220 50076
rect 44220 50020 44276 50076
rect 44276 50020 44280 50076
rect 44216 50016 44280 50020
rect 44296 50076 44360 50080
rect 44296 50020 44300 50076
rect 44300 50020 44356 50076
rect 44356 50020 44360 50076
rect 44296 50016 44360 50020
rect 44376 50076 44440 50080
rect 44376 50020 44380 50076
rect 44380 50020 44436 50076
rect 44436 50020 44440 50076
rect 44376 50016 44440 50020
rect 44456 50076 44520 50080
rect 44456 50020 44460 50076
rect 44460 50020 44516 50076
rect 44516 50020 44520 50076
rect 44456 50016 44520 50020
rect 54216 50076 54280 50080
rect 54216 50020 54220 50076
rect 54220 50020 54276 50076
rect 54276 50020 54280 50076
rect 54216 50016 54280 50020
rect 54296 50076 54360 50080
rect 54296 50020 54300 50076
rect 54300 50020 54356 50076
rect 54356 50020 54360 50076
rect 54296 50016 54360 50020
rect 54376 50076 54440 50080
rect 54376 50020 54380 50076
rect 54380 50020 54436 50076
rect 54436 50020 54440 50076
rect 54376 50016 54440 50020
rect 54456 50076 54520 50080
rect 54456 50020 54460 50076
rect 54460 50020 54516 50076
rect 54516 50020 54520 50076
rect 54456 50016 54520 50020
rect 64216 50076 64280 50080
rect 64216 50020 64220 50076
rect 64220 50020 64276 50076
rect 64276 50020 64280 50076
rect 64216 50016 64280 50020
rect 64296 50076 64360 50080
rect 64296 50020 64300 50076
rect 64300 50020 64356 50076
rect 64356 50020 64360 50076
rect 64296 50016 64360 50020
rect 64376 50076 64440 50080
rect 64376 50020 64380 50076
rect 64380 50020 64436 50076
rect 64436 50020 64440 50076
rect 64376 50016 64440 50020
rect 64456 50076 64520 50080
rect 64456 50020 64460 50076
rect 64460 50020 64516 50076
rect 64516 50020 64520 50076
rect 64456 50016 64520 50020
rect 9216 49532 9280 49536
rect 9216 49476 9220 49532
rect 9220 49476 9276 49532
rect 9276 49476 9280 49532
rect 9216 49472 9280 49476
rect 9296 49532 9360 49536
rect 9296 49476 9300 49532
rect 9300 49476 9356 49532
rect 9356 49476 9360 49532
rect 9296 49472 9360 49476
rect 9376 49532 9440 49536
rect 9376 49476 9380 49532
rect 9380 49476 9436 49532
rect 9436 49476 9440 49532
rect 9376 49472 9440 49476
rect 9456 49532 9520 49536
rect 9456 49476 9460 49532
rect 9460 49476 9516 49532
rect 9516 49476 9520 49532
rect 9456 49472 9520 49476
rect 19216 49532 19280 49536
rect 19216 49476 19220 49532
rect 19220 49476 19276 49532
rect 19276 49476 19280 49532
rect 19216 49472 19280 49476
rect 19296 49532 19360 49536
rect 19296 49476 19300 49532
rect 19300 49476 19356 49532
rect 19356 49476 19360 49532
rect 19296 49472 19360 49476
rect 19376 49532 19440 49536
rect 19376 49476 19380 49532
rect 19380 49476 19436 49532
rect 19436 49476 19440 49532
rect 19376 49472 19440 49476
rect 19456 49532 19520 49536
rect 19456 49476 19460 49532
rect 19460 49476 19516 49532
rect 19516 49476 19520 49532
rect 19456 49472 19520 49476
rect 29216 49532 29280 49536
rect 29216 49476 29220 49532
rect 29220 49476 29276 49532
rect 29276 49476 29280 49532
rect 29216 49472 29280 49476
rect 29296 49532 29360 49536
rect 29296 49476 29300 49532
rect 29300 49476 29356 49532
rect 29356 49476 29360 49532
rect 29296 49472 29360 49476
rect 29376 49532 29440 49536
rect 29376 49476 29380 49532
rect 29380 49476 29436 49532
rect 29436 49476 29440 49532
rect 29376 49472 29440 49476
rect 29456 49532 29520 49536
rect 29456 49476 29460 49532
rect 29460 49476 29516 49532
rect 29516 49476 29520 49532
rect 29456 49472 29520 49476
rect 39216 49532 39280 49536
rect 39216 49476 39220 49532
rect 39220 49476 39276 49532
rect 39276 49476 39280 49532
rect 39216 49472 39280 49476
rect 39296 49532 39360 49536
rect 39296 49476 39300 49532
rect 39300 49476 39356 49532
rect 39356 49476 39360 49532
rect 39296 49472 39360 49476
rect 39376 49532 39440 49536
rect 39376 49476 39380 49532
rect 39380 49476 39436 49532
rect 39436 49476 39440 49532
rect 39376 49472 39440 49476
rect 39456 49532 39520 49536
rect 39456 49476 39460 49532
rect 39460 49476 39516 49532
rect 39516 49476 39520 49532
rect 39456 49472 39520 49476
rect 49216 49532 49280 49536
rect 49216 49476 49220 49532
rect 49220 49476 49276 49532
rect 49276 49476 49280 49532
rect 49216 49472 49280 49476
rect 49296 49532 49360 49536
rect 49296 49476 49300 49532
rect 49300 49476 49356 49532
rect 49356 49476 49360 49532
rect 49296 49472 49360 49476
rect 49376 49532 49440 49536
rect 49376 49476 49380 49532
rect 49380 49476 49436 49532
rect 49436 49476 49440 49532
rect 49376 49472 49440 49476
rect 49456 49532 49520 49536
rect 49456 49476 49460 49532
rect 49460 49476 49516 49532
rect 49516 49476 49520 49532
rect 49456 49472 49520 49476
rect 59216 49532 59280 49536
rect 59216 49476 59220 49532
rect 59220 49476 59276 49532
rect 59276 49476 59280 49532
rect 59216 49472 59280 49476
rect 59296 49532 59360 49536
rect 59296 49476 59300 49532
rect 59300 49476 59356 49532
rect 59356 49476 59360 49532
rect 59296 49472 59360 49476
rect 59376 49532 59440 49536
rect 59376 49476 59380 49532
rect 59380 49476 59436 49532
rect 59436 49476 59440 49532
rect 59376 49472 59440 49476
rect 59456 49532 59520 49536
rect 59456 49476 59460 49532
rect 59460 49476 59516 49532
rect 59516 49476 59520 49532
rect 59456 49472 59520 49476
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 14216 48988 14280 48992
rect 14216 48932 14220 48988
rect 14220 48932 14276 48988
rect 14276 48932 14280 48988
rect 14216 48928 14280 48932
rect 14296 48988 14360 48992
rect 14296 48932 14300 48988
rect 14300 48932 14356 48988
rect 14356 48932 14360 48988
rect 14296 48928 14360 48932
rect 14376 48988 14440 48992
rect 14376 48932 14380 48988
rect 14380 48932 14436 48988
rect 14436 48932 14440 48988
rect 14376 48928 14440 48932
rect 14456 48988 14520 48992
rect 14456 48932 14460 48988
rect 14460 48932 14516 48988
rect 14516 48932 14520 48988
rect 14456 48928 14520 48932
rect 24216 48988 24280 48992
rect 24216 48932 24220 48988
rect 24220 48932 24276 48988
rect 24276 48932 24280 48988
rect 24216 48928 24280 48932
rect 24296 48988 24360 48992
rect 24296 48932 24300 48988
rect 24300 48932 24356 48988
rect 24356 48932 24360 48988
rect 24296 48928 24360 48932
rect 24376 48988 24440 48992
rect 24376 48932 24380 48988
rect 24380 48932 24436 48988
rect 24436 48932 24440 48988
rect 24376 48928 24440 48932
rect 24456 48988 24520 48992
rect 24456 48932 24460 48988
rect 24460 48932 24516 48988
rect 24516 48932 24520 48988
rect 24456 48928 24520 48932
rect 34216 48988 34280 48992
rect 34216 48932 34220 48988
rect 34220 48932 34276 48988
rect 34276 48932 34280 48988
rect 34216 48928 34280 48932
rect 34296 48988 34360 48992
rect 34296 48932 34300 48988
rect 34300 48932 34356 48988
rect 34356 48932 34360 48988
rect 34296 48928 34360 48932
rect 34376 48988 34440 48992
rect 34376 48932 34380 48988
rect 34380 48932 34436 48988
rect 34436 48932 34440 48988
rect 34376 48928 34440 48932
rect 34456 48988 34520 48992
rect 34456 48932 34460 48988
rect 34460 48932 34516 48988
rect 34516 48932 34520 48988
rect 34456 48928 34520 48932
rect 44216 48988 44280 48992
rect 44216 48932 44220 48988
rect 44220 48932 44276 48988
rect 44276 48932 44280 48988
rect 44216 48928 44280 48932
rect 44296 48988 44360 48992
rect 44296 48932 44300 48988
rect 44300 48932 44356 48988
rect 44356 48932 44360 48988
rect 44296 48928 44360 48932
rect 44376 48988 44440 48992
rect 44376 48932 44380 48988
rect 44380 48932 44436 48988
rect 44436 48932 44440 48988
rect 44376 48928 44440 48932
rect 44456 48988 44520 48992
rect 44456 48932 44460 48988
rect 44460 48932 44516 48988
rect 44516 48932 44520 48988
rect 44456 48928 44520 48932
rect 54216 48988 54280 48992
rect 54216 48932 54220 48988
rect 54220 48932 54276 48988
rect 54276 48932 54280 48988
rect 54216 48928 54280 48932
rect 54296 48988 54360 48992
rect 54296 48932 54300 48988
rect 54300 48932 54356 48988
rect 54356 48932 54360 48988
rect 54296 48928 54360 48932
rect 54376 48988 54440 48992
rect 54376 48932 54380 48988
rect 54380 48932 54436 48988
rect 54436 48932 54440 48988
rect 54376 48928 54440 48932
rect 54456 48988 54520 48992
rect 54456 48932 54460 48988
rect 54460 48932 54516 48988
rect 54516 48932 54520 48988
rect 54456 48928 54520 48932
rect 64216 48988 64280 48992
rect 64216 48932 64220 48988
rect 64220 48932 64276 48988
rect 64276 48932 64280 48988
rect 64216 48928 64280 48932
rect 64296 48988 64360 48992
rect 64296 48932 64300 48988
rect 64300 48932 64356 48988
rect 64356 48932 64360 48988
rect 64296 48928 64360 48932
rect 64376 48988 64440 48992
rect 64376 48932 64380 48988
rect 64380 48932 64436 48988
rect 64436 48932 64440 48988
rect 64376 48928 64440 48932
rect 64456 48988 64520 48992
rect 64456 48932 64460 48988
rect 64460 48932 64516 48988
rect 64516 48932 64520 48988
rect 64456 48928 64520 48932
rect 9216 48444 9280 48448
rect 9216 48388 9220 48444
rect 9220 48388 9276 48444
rect 9276 48388 9280 48444
rect 9216 48384 9280 48388
rect 9296 48444 9360 48448
rect 9296 48388 9300 48444
rect 9300 48388 9356 48444
rect 9356 48388 9360 48444
rect 9296 48384 9360 48388
rect 9376 48444 9440 48448
rect 9376 48388 9380 48444
rect 9380 48388 9436 48444
rect 9436 48388 9440 48444
rect 9376 48384 9440 48388
rect 9456 48444 9520 48448
rect 9456 48388 9460 48444
rect 9460 48388 9516 48444
rect 9516 48388 9520 48444
rect 9456 48384 9520 48388
rect 19216 48444 19280 48448
rect 19216 48388 19220 48444
rect 19220 48388 19276 48444
rect 19276 48388 19280 48444
rect 19216 48384 19280 48388
rect 19296 48444 19360 48448
rect 19296 48388 19300 48444
rect 19300 48388 19356 48444
rect 19356 48388 19360 48444
rect 19296 48384 19360 48388
rect 19376 48444 19440 48448
rect 19376 48388 19380 48444
rect 19380 48388 19436 48444
rect 19436 48388 19440 48444
rect 19376 48384 19440 48388
rect 19456 48444 19520 48448
rect 19456 48388 19460 48444
rect 19460 48388 19516 48444
rect 19516 48388 19520 48444
rect 19456 48384 19520 48388
rect 29216 48444 29280 48448
rect 29216 48388 29220 48444
rect 29220 48388 29276 48444
rect 29276 48388 29280 48444
rect 29216 48384 29280 48388
rect 29296 48444 29360 48448
rect 29296 48388 29300 48444
rect 29300 48388 29356 48444
rect 29356 48388 29360 48444
rect 29296 48384 29360 48388
rect 29376 48444 29440 48448
rect 29376 48388 29380 48444
rect 29380 48388 29436 48444
rect 29436 48388 29440 48444
rect 29376 48384 29440 48388
rect 29456 48444 29520 48448
rect 29456 48388 29460 48444
rect 29460 48388 29516 48444
rect 29516 48388 29520 48444
rect 29456 48384 29520 48388
rect 39216 48444 39280 48448
rect 39216 48388 39220 48444
rect 39220 48388 39276 48444
rect 39276 48388 39280 48444
rect 39216 48384 39280 48388
rect 39296 48444 39360 48448
rect 39296 48388 39300 48444
rect 39300 48388 39356 48444
rect 39356 48388 39360 48444
rect 39296 48384 39360 48388
rect 39376 48444 39440 48448
rect 39376 48388 39380 48444
rect 39380 48388 39436 48444
rect 39436 48388 39440 48444
rect 39376 48384 39440 48388
rect 39456 48444 39520 48448
rect 39456 48388 39460 48444
rect 39460 48388 39516 48444
rect 39516 48388 39520 48444
rect 39456 48384 39520 48388
rect 49216 48444 49280 48448
rect 49216 48388 49220 48444
rect 49220 48388 49276 48444
rect 49276 48388 49280 48444
rect 49216 48384 49280 48388
rect 49296 48444 49360 48448
rect 49296 48388 49300 48444
rect 49300 48388 49356 48444
rect 49356 48388 49360 48444
rect 49296 48384 49360 48388
rect 49376 48444 49440 48448
rect 49376 48388 49380 48444
rect 49380 48388 49436 48444
rect 49436 48388 49440 48444
rect 49376 48384 49440 48388
rect 49456 48444 49520 48448
rect 49456 48388 49460 48444
rect 49460 48388 49516 48444
rect 49516 48388 49520 48444
rect 49456 48384 49520 48388
rect 59216 48444 59280 48448
rect 59216 48388 59220 48444
rect 59220 48388 59276 48444
rect 59276 48388 59280 48444
rect 59216 48384 59280 48388
rect 59296 48444 59360 48448
rect 59296 48388 59300 48444
rect 59300 48388 59356 48444
rect 59356 48388 59360 48444
rect 59296 48384 59360 48388
rect 59376 48444 59440 48448
rect 59376 48388 59380 48444
rect 59380 48388 59436 48444
rect 59436 48388 59440 48444
rect 59376 48384 59440 48388
rect 59456 48444 59520 48448
rect 59456 48388 59460 48444
rect 59460 48388 59516 48444
rect 59516 48388 59520 48444
rect 59456 48384 59520 48388
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 14216 47900 14280 47904
rect 14216 47844 14220 47900
rect 14220 47844 14276 47900
rect 14276 47844 14280 47900
rect 14216 47840 14280 47844
rect 14296 47900 14360 47904
rect 14296 47844 14300 47900
rect 14300 47844 14356 47900
rect 14356 47844 14360 47900
rect 14296 47840 14360 47844
rect 14376 47900 14440 47904
rect 14376 47844 14380 47900
rect 14380 47844 14436 47900
rect 14436 47844 14440 47900
rect 14376 47840 14440 47844
rect 14456 47900 14520 47904
rect 14456 47844 14460 47900
rect 14460 47844 14516 47900
rect 14516 47844 14520 47900
rect 14456 47840 14520 47844
rect 24216 47900 24280 47904
rect 24216 47844 24220 47900
rect 24220 47844 24276 47900
rect 24276 47844 24280 47900
rect 24216 47840 24280 47844
rect 24296 47900 24360 47904
rect 24296 47844 24300 47900
rect 24300 47844 24356 47900
rect 24356 47844 24360 47900
rect 24296 47840 24360 47844
rect 24376 47900 24440 47904
rect 24376 47844 24380 47900
rect 24380 47844 24436 47900
rect 24436 47844 24440 47900
rect 24376 47840 24440 47844
rect 24456 47900 24520 47904
rect 24456 47844 24460 47900
rect 24460 47844 24516 47900
rect 24516 47844 24520 47900
rect 24456 47840 24520 47844
rect 34216 47900 34280 47904
rect 34216 47844 34220 47900
rect 34220 47844 34276 47900
rect 34276 47844 34280 47900
rect 34216 47840 34280 47844
rect 34296 47900 34360 47904
rect 34296 47844 34300 47900
rect 34300 47844 34356 47900
rect 34356 47844 34360 47900
rect 34296 47840 34360 47844
rect 34376 47900 34440 47904
rect 34376 47844 34380 47900
rect 34380 47844 34436 47900
rect 34436 47844 34440 47900
rect 34376 47840 34440 47844
rect 34456 47900 34520 47904
rect 34456 47844 34460 47900
rect 34460 47844 34516 47900
rect 34516 47844 34520 47900
rect 34456 47840 34520 47844
rect 44216 47900 44280 47904
rect 44216 47844 44220 47900
rect 44220 47844 44276 47900
rect 44276 47844 44280 47900
rect 44216 47840 44280 47844
rect 44296 47900 44360 47904
rect 44296 47844 44300 47900
rect 44300 47844 44356 47900
rect 44356 47844 44360 47900
rect 44296 47840 44360 47844
rect 44376 47900 44440 47904
rect 44376 47844 44380 47900
rect 44380 47844 44436 47900
rect 44436 47844 44440 47900
rect 44376 47840 44440 47844
rect 44456 47900 44520 47904
rect 44456 47844 44460 47900
rect 44460 47844 44516 47900
rect 44516 47844 44520 47900
rect 44456 47840 44520 47844
rect 54216 47900 54280 47904
rect 54216 47844 54220 47900
rect 54220 47844 54276 47900
rect 54276 47844 54280 47900
rect 54216 47840 54280 47844
rect 54296 47900 54360 47904
rect 54296 47844 54300 47900
rect 54300 47844 54356 47900
rect 54356 47844 54360 47900
rect 54296 47840 54360 47844
rect 54376 47900 54440 47904
rect 54376 47844 54380 47900
rect 54380 47844 54436 47900
rect 54436 47844 54440 47900
rect 54376 47840 54440 47844
rect 54456 47900 54520 47904
rect 54456 47844 54460 47900
rect 54460 47844 54516 47900
rect 54516 47844 54520 47900
rect 54456 47840 54520 47844
rect 64216 47900 64280 47904
rect 64216 47844 64220 47900
rect 64220 47844 64276 47900
rect 64276 47844 64280 47900
rect 64216 47840 64280 47844
rect 64296 47900 64360 47904
rect 64296 47844 64300 47900
rect 64300 47844 64356 47900
rect 64356 47844 64360 47900
rect 64296 47840 64360 47844
rect 64376 47900 64440 47904
rect 64376 47844 64380 47900
rect 64380 47844 64436 47900
rect 64436 47844 64440 47900
rect 64376 47840 64440 47844
rect 64456 47900 64520 47904
rect 64456 47844 64460 47900
rect 64460 47844 64516 47900
rect 64516 47844 64520 47900
rect 64456 47840 64520 47844
rect 9216 47356 9280 47360
rect 9216 47300 9220 47356
rect 9220 47300 9276 47356
rect 9276 47300 9280 47356
rect 9216 47296 9280 47300
rect 9296 47356 9360 47360
rect 9296 47300 9300 47356
rect 9300 47300 9356 47356
rect 9356 47300 9360 47356
rect 9296 47296 9360 47300
rect 9376 47356 9440 47360
rect 9376 47300 9380 47356
rect 9380 47300 9436 47356
rect 9436 47300 9440 47356
rect 9376 47296 9440 47300
rect 9456 47356 9520 47360
rect 9456 47300 9460 47356
rect 9460 47300 9516 47356
rect 9516 47300 9520 47356
rect 9456 47296 9520 47300
rect 19216 47356 19280 47360
rect 19216 47300 19220 47356
rect 19220 47300 19276 47356
rect 19276 47300 19280 47356
rect 19216 47296 19280 47300
rect 19296 47356 19360 47360
rect 19296 47300 19300 47356
rect 19300 47300 19356 47356
rect 19356 47300 19360 47356
rect 19296 47296 19360 47300
rect 19376 47356 19440 47360
rect 19376 47300 19380 47356
rect 19380 47300 19436 47356
rect 19436 47300 19440 47356
rect 19376 47296 19440 47300
rect 19456 47356 19520 47360
rect 19456 47300 19460 47356
rect 19460 47300 19516 47356
rect 19516 47300 19520 47356
rect 19456 47296 19520 47300
rect 29216 47356 29280 47360
rect 29216 47300 29220 47356
rect 29220 47300 29276 47356
rect 29276 47300 29280 47356
rect 29216 47296 29280 47300
rect 29296 47356 29360 47360
rect 29296 47300 29300 47356
rect 29300 47300 29356 47356
rect 29356 47300 29360 47356
rect 29296 47296 29360 47300
rect 29376 47356 29440 47360
rect 29376 47300 29380 47356
rect 29380 47300 29436 47356
rect 29436 47300 29440 47356
rect 29376 47296 29440 47300
rect 29456 47356 29520 47360
rect 29456 47300 29460 47356
rect 29460 47300 29516 47356
rect 29516 47300 29520 47356
rect 29456 47296 29520 47300
rect 39216 47356 39280 47360
rect 39216 47300 39220 47356
rect 39220 47300 39276 47356
rect 39276 47300 39280 47356
rect 39216 47296 39280 47300
rect 39296 47356 39360 47360
rect 39296 47300 39300 47356
rect 39300 47300 39356 47356
rect 39356 47300 39360 47356
rect 39296 47296 39360 47300
rect 39376 47356 39440 47360
rect 39376 47300 39380 47356
rect 39380 47300 39436 47356
rect 39436 47300 39440 47356
rect 39376 47296 39440 47300
rect 39456 47356 39520 47360
rect 39456 47300 39460 47356
rect 39460 47300 39516 47356
rect 39516 47300 39520 47356
rect 39456 47296 39520 47300
rect 49216 47356 49280 47360
rect 49216 47300 49220 47356
rect 49220 47300 49276 47356
rect 49276 47300 49280 47356
rect 49216 47296 49280 47300
rect 49296 47356 49360 47360
rect 49296 47300 49300 47356
rect 49300 47300 49356 47356
rect 49356 47300 49360 47356
rect 49296 47296 49360 47300
rect 49376 47356 49440 47360
rect 49376 47300 49380 47356
rect 49380 47300 49436 47356
rect 49436 47300 49440 47356
rect 49376 47296 49440 47300
rect 49456 47356 49520 47360
rect 49456 47300 49460 47356
rect 49460 47300 49516 47356
rect 49516 47300 49520 47356
rect 49456 47296 49520 47300
rect 59216 47356 59280 47360
rect 59216 47300 59220 47356
rect 59220 47300 59276 47356
rect 59276 47300 59280 47356
rect 59216 47296 59280 47300
rect 59296 47356 59360 47360
rect 59296 47300 59300 47356
rect 59300 47300 59356 47356
rect 59356 47300 59360 47356
rect 59296 47296 59360 47300
rect 59376 47356 59440 47360
rect 59376 47300 59380 47356
rect 59380 47300 59436 47356
rect 59436 47300 59440 47356
rect 59376 47296 59440 47300
rect 59456 47356 59520 47360
rect 59456 47300 59460 47356
rect 59460 47300 59516 47356
rect 59516 47300 59520 47356
rect 59456 47296 59520 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 14216 46812 14280 46816
rect 14216 46756 14220 46812
rect 14220 46756 14276 46812
rect 14276 46756 14280 46812
rect 14216 46752 14280 46756
rect 14296 46812 14360 46816
rect 14296 46756 14300 46812
rect 14300 46756 14356 46812
rect 14356 46756 14360 46812
rect 14296 46752 14360 46756
rect 14376 46812 14440 46816
rect 14376 46756 14380 46812
rect 14380 46756 14436 46812
rect 14436 46756 14440 46812
rect 14376 46752 14440 46756
rect 14456 46812 14520 46816
rect 14456 46756 14460 46812
rect 14460 46756 14516 46812
rect 14516 46756 14520 46812
rect 14456 46752 14520 46756
rect 24216 46812 24280 46816
rect 24216 46756 24220 46812
rect 24220 46756 24276 46812
rect 24276 46756 24280 46812
rect 24216 46752 24280 46756
rect 24296 46812 24360 46816
rect 24296 46756 24300 46812
rect 24300 46756 24356 46812
rect 24356 46756 24360 46812
rect 24296 46752 24360 46756
rect 24376 46812 24440 46816
rect 24376 46756 24380 46812
rect 24380 46756 24436 46812
rect 24436 46756 24440 46812
rect 24376 46752 24440 46756
rect 24456 46812 24520 46816
rect 24456 46756 24460 46812
rect 24460 46756 24516 46812
rect 24516 46756 24520 46812
rect 24456 46752 24520 46756
rect 34216 46812 34280 46816
rect 34216 46756 34220 46812
rect 34220 46756 34276 46812
rect 34276 46756 34280 46812
rect 34216 46752 34280 46756
rect 34296 46812 34360 46816
rect 34296 46756 34300 46812
rect 34300 46756 34356 46812
rect 34356 46756 34360 46812
rect 34296 46752 34360 46756
rect 34376 46812 34440 46816
rect 34376 46756 34380 46812
rect 34380 46756 34436 46812
rect 34436 46756 34440 46812
rect 34376 46752 34440 46756
rect 34456 46812 34520 46816
rect 34456 46756 34460 46812
rect 34460 46756 34516 46812
rect 34516 46756 34520 46812
rect 34456 46752 34520 46756
rect 44216 46812 44280 46816
rect 44216 46756 44220 46812
rect 44220 46756 44276 46812
rect 44276 46756 44280 46812
rect 44216 46752 44280 46756
rect 44296 46812 44360 46816
rect 44296 46756 44300 46812
rect 44300 46756 44356 46812
rect 44356 46756 44360 46812
rect 44296 46752 44360 46756
rect 44376 46812 44440 46816
rect 44376 46756 44380 46812
rect 44380 46756 44436 46812
rect 44436 46756 44440 46812
rect 44376 46752 44440 46756
rect 44456 46812 44520 46816
rect 44456 46756 44460 46812
rect 44460 46756 44516 46812
rect 44516 46756 44520 46812
rect 44456 46752 44520 46756
rect 54216 46812 54280 46816
rect 54216 46756 54220 46812
rect 54220 46756 54276 46812
rect 54276 46756 54280 46812
rect 54216 46752 54280 46756
rect 54296 46812 54360 46816
rect 54296 46756 54300 46812
rect 54300 46756 54356 46812
rect 54356 46756 54360 46812
rect 54296 46752 54360 46756
rect 54376 46812 54440 46816
rect 54376 46756 54380 46812
rect 54380 46756 54436 46812
rect 54436 46756 54440 46812
rect 54376 46752 54440 46756
rect 54456 46812 54520 46816
rect 54456 46756 54460 46812
rect 54460 46756 54516 46812
rect 54516 46756 54520 46812
rect 54456 46752 54520 46756
rect 64216 46812 64280 46816
rect 64216 46756 64220 46812
rect 64220 46756 64276 46812
rect 64276 46756 64280 46812
rect 64216 46752 64280 46756
rect 64296 46812 64360 46816
rect 64296 46756 64300 46812
rect 64300 46756 64356 46812
rect 64356 46756 64360 46812
rect 64296 46752 64360 46756
rect 64376 46812 64440 46816
rect 64376 46756 64380 46812
rect 64380 46756 64436 46812
rect 64436 46756 64440 46812
rect 64376 46752 64440 46756
rect 64456 46812 64520 46816
rect 64456 46756 64460 46812
rect 64460 46756 64516 46812
rect 64516 46756 64520 46812
rect 64456 46752 64520 46756
rect 9216 46268 9280 46272
rect 9216 46212 9220 46268
rect 9220 46212 9276 46268
rect 9276 46212 9280 46268
rect 9216 46208 9280 46212
rect 9296 46268 9360 46272
rect 9296 46212 9300 46268
rect 9300 46212 9356 46268
rect 9356 46212 9360 46268
rect 9296 46208 9360 46212
rect 9376 46268 9440 46272
rect 9376 46212 9380 46268
rect 9380 46212 9436 46268
rect 9436 46212 9440 46268
rect 9376 46208 9440 46212
rect 9456 46268 9520 46272
rect 9456 46212 9460 46268
rect 9460 46212 9516 46268
rect 9516 46212 9520 46268
rect 9456 46208 9520 46212
rect 19216 46268 19280 46272
rect 19216 46212 19220 46268
rect 19220 46212 19276 46268
rect 19276 46212 19280 46268
rect 19216 46208 19280 46212
rect 19296 46268 19360 46272
rect 19296 46212 19300 46268
rect 19300 46212 19356 46268
rect 19356 46212 19360 46268
rect 19296 46208 19360 46212
rect 19376 46268 19440 46272
rect 19376 46212 19380 46268
rect 19380 46212 19436 46268
rect 19436 46212 19440 46268
rect 19376 46208 19440 46212
rect 19456 46268 19520 46272
rect 19456 46212 19460 46268
rect 19460 46212 19516 46268
rect 19516 46212 19520 46268
rect 19456 46208 19520 46212
rect 29216 46268 29280 46272
rect 29216 46212 29220 46268
rect 29220 46212 29276 46268
rect 29276 46212 29280 46268
rect 29216 46208 29280 46212
rect 29296 46268 29360 46272
rect 29296 46212 29300 46268
rect 29300 46212 29356 46268
rect 29356 46212 29360 46268
rect 29296 46208 29360 46212
rect 29376 46268 29440 46272
rect 29376 46212 29380 46268
rect 29380 46212 29436 46268
rect 29436 46212 29440 46268
rect 29376 46208 29440 46212
rect 29456 46268 29520 46272
rect 29456 46212 29460 46268
rect 29460 46212 29516 46268
rect 29516 46212 29520 46268
rect 29456 46208 29520 46212
rect 39216 46268 39280 46272
rect 39216 46212 39220 46268
rect 39220 46212 39276 46268
rect 39276 46212 39280 46268
rect 39216 46208 39280 46212
rect 39296 46268 39360 46272
rect 39296 46212 39300 46268
rect 39300 46212 39356 46268
rect 39356 46212 39360 46268
rect 39296 46208 39360 46212
rect 39376 46268 39440 46272
rect 39376 46212 39380 46268
rect 39380 46212 39436 46268
rect 39436 46212 39440 46268
rect 39376 46208 39440 46212
rect 39456 46268 39520 46272
rect 39456 46212 39460 46268
rect 39460 46212 39516 46268
rect 39516 46212 39520 46268
rect 39456 46208 39520 46212
rect 49216 46268 49280 46272
rect 49216 46212 49220 46268
rect 49220 46212 49276 46268
rect 49276 46212 49280 46268
rect 49216 46208 49280 46212
rect 49296 46268 49360 46272
rect 49296 46212 49300 46268
rect 49300 46212 49356 46268
rect 49356 46212 49360 46268
rect 49296 46208 49360 46212
rect 49376 46268 49440 46272
rect 49376 46212 49380 46268
rect 49380 46212 49436 46268
rect 49436 46212 49440 46268
rect 49376 46208 49440 46212
rect 49456 46268 49520 46272
rect 49456 46212 49460 46268
rect 49460 46212 49516 46268
rect 49516 46212 49520 46268
rect 49456 46208 49520 46212
rect 59216 46268 59280 46272
rect 59216 46212 59220 46268
rect 59220 46212 59276 46268
rect 59276 46212 59280 46268
rect 59216 46208 59280 46212
rect 59296 46268 59360 46272
rect 59296 46212 59300 46268
rect 59300 46212 59356 46268
rect 59356 46212 59360 46268
rect 59296 46208 59360 46212
rect 59376 46268 59440 46272
rect 59376 46212 59380 46268
rect 59380 46212 59436 46268
rect 59436 46212 59440 46268
rect 59376 46208 59440 46212
rect 59456 46268 59520 46272
rect 59456 46212 59460 46268
rect 59460 46212 59516 46268
rect 59516 46212 59520 46268
rect 59456 46208 59520 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 14216 45724 14280 45728
rect 14216 45668 14220 45724
rect 14220 45668 14276 45724
rect 14276 45668 14280 45724
rect 14216 45664 14280 45668
rect 14296 45724 14360 45728
rect 14296 45668 14300 45724
rect 14300 45668 14356 45724
rect 14356 45668 14360 45724
rect 14296 45664 14360 45668
rect 14376 45724 14440 45728
rect 14376 45668 14380 45724
rect 14380 45668 14436 45724
rect 14436 45668 14440 45724
rect 14376 45664 14440 45668
rect 14456 45724 14520 45728
rect 14456 45668 14460 45724
rect 14460 45668 14516 45724
rect 14516 45668 14520 45724
rect 14456 45664 14520 45668
rect 24216 45724 24280 45728
rect 24216 45668 24220 45724
rect 24220 45668 24276 45724
rect 24276 45668 24280 45724
rect 24216 45664 24280 45668
rect 24296 45724 24360 45728
rect 24296 45668 24300 45724
rect 24300 45668 24356 45724
rect 24356 45668 24360 45724
rect 24296 45664 24360 45668
rect 24376 45724 24440 45728
rect 24376 45668 24380 45724
rect 24380 45668 24436 45724
rect 24436 45668 24440 45724
rect 24376 45664 24440 45668
rect 24456 45724 24520 45728
rect 24456 45668 24460 45724
rect 24460 45668 24516 45724
rect 24516 45668 24520 45724
rect 24456 45664 24520 45668
rect 34216 45724 34280 45728
rect 34216 45668 34220 45724
rect 34220 45668 34276 45724
rect 34276 45668 34280 45724
rect 34216 45664 34280 45668
rect 34296 45724 34360 45728
rect 34296 45668 34300 45724
rect 34300 45668 34356 45724
rect 34356 45668 34360 45724
rect 34296 45664 34360 45668
rect 34376 45724 34440 45728
rect 34376 45668 34380 45724
rect 34380 45668 34436 45724
rect 34436 45668 34440 45724
rect 34376 45664 34440 45668
rect 34456 45724 34520 45728
rect 34456 45668 34460 45724
rect 34460 45668 34516 45724
rect 34516 45668 34520 45724
rect 34456 45664 34520 45668
rect 44216 45724 44280 45728
rect 44216 45668 44220 45724
rect 44220 45668 44276 45724
rect 44276 45668 44280 45724
rect 44216 45664 44280 45668
rect 44296 45724 44360 45728
rect 44296 45668 44300 45724
rect 44300 45668 44356 45724
rect 44356 45668 44360 45724
rect 44296 45664 44360 45668
rect 44376 45724 44440 45728
rect 44376 45668 44380 45724
rect 44380 45668 44436 45724
rect 44436 45668 44440 45724
rect 44376 45664 44440 45668
rect 44456 45724 44520 45728
rect 44456 45668 44460 45724
rect 44460 45668 44516 45724
rect 44516 45668 44520 45724
rect 44456 45664 44520 45668
rect 54216 45724 54280 45728
rect 54216 45668 54220 45724
rect 54220 45668 54276 45724
rect 54276 45668 54280 45724
rect 54216 45664 54280 45668
rect 54296 45724 54360 45728
rect 54296 45668 54300 45724
rect 54300 45668 54356 45724
rect 54356 45668 54360 45724
rect 54296 45664 54360 45668
rect 54376 45724 54440 45728
rect 54376 45668 54380 45724
rect 54380 45668 54436 45724
rect 54436 45668 54440 45724
rect 54376 45664 54440 45668
rect 54456 45724 54520 45728
rect 54456 45668 54460 45724
rect 54460 45668 54516 45724
rect 54516 45668 54520 45724
rect 54456 45664 54520 45668
rect 64216 45724 64280 45728
rect 64216 45668 64220 45724
rect 64220 45668 64276 45724
rect 64276 45668 64280 45724
rect 64216 45664 64280 45668
rect 64296 45724 64360 45728
rect 64296 45668 64300 45724
rect 64300 45668 64356 45724
rect 64356 45668 64360 45724
rect 64296 45664 64360 45668
rect 64376 45724 64440 45728
rect 64376 45668 64380 45724
rect 64380 45668 64436 45724
rect 64436 45668 64440 45724
rect 64376 45664 64440 45668
rect 64456 45724 64520 45728
rect 64456 45668 64460 45724
rect 64460 45668 64516 45724
rect 64516 45668 64520 45724
rect 64456 45664 64520 45668
rect 9216 45180 9280 45184
rect 9216 45124 9220 45180
rect 9220 45124 9276 45180
rect 9276 45124 9280 45180
rect 9216 45120 9280 45124
rect 9296 45180 9360 45184
rect 9296 45124 9300 45180
rect 9300 45124 9356 45180
rect 9356 45124 9360 45180
rect 9296 45120 9360 45124
rect 9376 45180 9440 45184
rect 9376 45124 9380 45180
rect 9380 45124 9436 45180
rect 9436 45124 9440 45180
rect 9376 45120 9440 45124
rect 9456 45180 9520 45184
rect 9456 45124 9460 45180
rect 9460 45124 9516 45180
rect 9516 45124 9520 45180
rect 9456 45120 9520 45124
rect 19216 45180 19280 45184
rect 19216 45124 19220 45180
rect 19220 45124 19276 45180
rect 19276 45124 19280 45180
rect 19216 45120 19280 45124
rect 19296 45180 19360 45184
rect 19296 45124 19300 45180
rect 19300 45124 19356 45180
rect 19356 45124 19360 45180
rect 19296 45120 19360 45124
rect 19376 45180 19440 45184
rect 19376 45124 19380 45180
rect 19380 45124 19436 45180
rect 19436 45124 19440 45180
rect 19376 45120 19440 45124
rect 19456 45180 19520 45184
rect 19456 45124 19460 45180
rect 19460 45124 19516 45180
rect 19516 45124 19520 45180
rect 19456 45120 19520 45124
rect 29216 45180 29280 45184
rect 29216 45124 29220 45180
rect 29220 45124 29276 45180
rect 29276 45124 29280 45180
rect 29216 45120 29280 45124
rect 29296 45180 29360 45184
rect 29296 45124 29300 45180
rect 29300 45124 29356 45180
rect 29356 45124 29360 45180
rect 29296 45120 29360 45124
rect 29376 45180 29440 45184
rect 29376 45124 29380 45180
rect 29380 45124 29436 45180
rect 29436 45124 29440 45180
rect 29376 45120 29440 45124
rect 29456 45180 29520 45184
rect 29456 45124 29460 45180
rect 29460 45124 29516 45180
rect 29516 45124 29520 45180
rect 29456 45120 29520 45124
rect 39216 45180 39280 45184
rect 39216 45124 39220 45180
rect 39220 45124 39276 45180
rect 39276 45124 39280 45180
rect 39216 45120 39280 45124
rect 39296 45180 39360 45184
rect 39296 45124 39300 45180
rect 39300 45124 39356 45180
rect 39356 45124 39360 45180
rect 39296 45120 39360 45124
rect 39376 45180 39440 45184
rect 39376 45124 39380 45180
rect 39380 45124 39436 45180
rect 39436 45124 39440 45180
rect 39376 45120 39440 45124
rect 39456 45180 39520 45184
rect 39456 45124 39460 45180
rect 39460 45124 39516 45180
rect 39516 45124 39520 45180
rect 39456 45120 39520 45124
rect 49216 45180 49280 45184
rect 49216 45124 49220 45180
rect 49220 45124 49276 45180
rect 49276 45124 49280 45180
rect 49216 45120 49280 45124
rect 49296 45180 49360 45184
rect 49296 45124 49300 45180
rect 49300 45124 49356 45180
rect 49356 45124 49360 45180
rect 49296 45120 49360 45124
rect 49376 45180 49440 45184
rect 49376 45124 49380 45180
rect 49380 45124 49436 45180
rect 49436 45124 49440 45180
rect 49376 45120 49440 45124
rect 49456 45180 49520 45184
rect 49456 45124 49460 45180
rect 49460 45124 49516 45180
rect 49516 45124 49520 45180
rect 49456 45120 49520 45124
rect 59216 45180 59280 45184
rect 59216 45124 59220 45180
rect 59220 45124 59276 45180
rect 59276 45124 59280 45180
rect 59216 45120 59280 45124
rect 59296 45180 59360 45184
rect 59296 45124 59300 45180
rect 59300 45124 59356 45180
rect 59356 45124 59360 45180
rect 59296 45120 59360 45124
rect 59376 45180 59440 45184
rect 59376 45124 59380 45180
rect 59380 45124 59436 45180
rect 59436 45124 59440 45180
rect 59376 45120 59440 45124
rect 59456 45180 59520 45184
rect 59456 45124 59460 45180
rect 59460 45124 59516 45180
rect 59516 45124 59520 45180
rect 59456 45120 59520 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 14216 44636 14280 44640
rect 14216 44580 14220 44636
rect 14220 44580 14276 44636
rect 14276 44580 14280 44636
rect 14216 44576 14280 44580
rect 14296 44636 14360 44640
rect 14296 44580 14300 44636
rect 14300 44580 14356 44636
rect 14356 44580 14360 44636
rect 14296 44576 14360 44580
rect 14376 44636 14440 44640
rect 14376 44580 14380 44636
rect 14380 44580 14436 44636
rect 14436 44580 14440 44636
rect 14376 44576 14440 44580
rect 14456 44636 14520 44640
rect 14456 44580 14460 44636
rect 14460 44580 14516 44636
rect 14516 44580 14520 44636
rect 14456 44576 14520 44580
rect 24216 44636 24280 44640
rect 24216 44580 24220 44636
rect 24220 44580 24276 44636
rect 24276 44580 24280 44636
rect 24216 44576 24280 44580
rect 24296 44636 24360 44640
rect 24296 44580 24300 44636
rect 24300 44580 24356 44636
rect 24356 44580 24360 44636
rect 24296 44576 24360 44580
rect 24376 44636 24440 44640
rect 24376 44580 24380 44636
rect 24380 44580 24436 44636
rect 24436 44580 24440 44636
rect 24376 44576 24440 44580
rect 24456 44636 24520 44640
rect 24456 44580 24460 44636
rect 24460 44580 24516 44636
rect 24516 44580 24520 44636
rect 24456 44576 24520 44580
rect 34216 44636 34280 44640
rect 34216 44580 34220 44636
rect 34220 44580 34276 44636
rect 34276 44580 34280 44636
rect 34216 44576 34280 44580
rect 34296 44636 34360 44640
rect 34296 44580 34300 44636
rect 34300 44580 34356 44636
rect 34356 44580 34360 44636
rect 34296 44576 34360 44580
rect 34376 44636 34440 44640
rect 34376 44580 34380 44636
rect 34380 44580 34436 44636
rect 34436 44580 34440 44636
rect 34376 44576 34440 44580
rect 34456 44636 34520 44640
rect 34456 44580 34460 44636
rect 34460 44580 34516 44636
rect 34516 44580 34520 44636
rect 34456 44576 34520 44580
rect 44216 44636 44280 44640
rect 44216 44580 44220 44636
rect 44220 44580 44276 44636
rect 44276 44580 44280 44636
rect 44216 44576 44280 44580
rect 44296 44636 44360 44640
rect 44296 44580 44300 44636
rect 44300 44580 44356 44636
rect 44356 44580 44360 44636
rect 44296 44576 44360 44580
rect 44376 44636 44440 44640
rect 44376 44580 44380 44636
rect 44380 44580 44436 44636
rect 44436 44580 44440 44636
rect 44376 44576 44440 44580
rect 44456 44636 44520 44640
rect 44456 44580 44460 44636
rect 44460 44580 44516 44636
rect 44516 44580 44520 44636
rect 44456 44576 44520 44580
rect 54216 44636 54280 44640
rect 54216 44580 54220 44636
rect 54220 44580 54276 44636
rect 54276 44580 54280 44636
rect 54216 44576 54280 44580
rect 54296 44636 54360 44640
rect 54296 44580 54300 44636
rect 54300 44580 54356 44636
rect 54356 44580 54360 44636
rect 54296 44576 54360 44580
rect 54376 44636 54440 44640
rect 54376 44580 54380 44636
rect 54380 44580 54436 44636
rect 54436 44580 54440 44636
rect 54376 44576 54440 44580
rect 54456 44636 54520 44640
rect 54456 44580 54460 44636
rect 54460 44580 54516 44636
rect 54516 44580 54520 44636
rect 54456 44576 54520 44580
rect 64216 44636 64280 44640
rect 64216 44580 64220 44636
rect 64220 44580 64276 44636
rect 64276 44580 64280 44636
rect 64216 44576 64280 44580
rect 64296 44636 64360 44640
rect 64296 44580 64300 44636
rect 64300 44580 64356 44636
rect 64356 44580 64360 44636
rect 64296 44576 64360 44580
rect 64376 44636 64440 44640
rect 64376 44580 64380 44636
rect 64380 44580 64436 44636
rect 64436 44580 64440 44636
rect 64376 44576 64440 44580
rect 64456 44636 64520 44640
rect 64456 44580 64460 44636
rect 64460 44580 64516 44636
rect 64516 44580 64520 44636
rect 64456 44576 64520 44580
rect 9216 44092 9280 44096
rect 9216 44036 9220 44092
rect 9220 44036 9276 44092
rect 9276 44036 9280 44092
rect 9216 44032 9280 44036
rect 9296 44092 9360 44096
rect 9296 44036 9300 44092
rect 9300 44036 9356 44092
rect 9356 44036 9360 44092
rect 9296 44032 9360 44036
rect 9376 44092 9440 44096
rect 9376 44036 9380 44092
rect 9380 44036 9436 44092
rect 9436 44036 9440 44092
rect 9376 44032 9440 44036
rect 9456 44092 9520 44096
rect 9456 44036 9460 44092
rect 9460 44036 9516 44092
rect 9516 44036 9520 44092
rect 9456 44032 9520 44036
rect 19216 44092 19280 44096
rect 19216 44036 19220 44092
rect 19220 44036 19276 44092
rect 19276 44036 19280 44092
rect 19216 44032 19280 44036
rect 19296 44092 19360 44096
rect 19296 44036 19300 44092
rect 19300 44036 19356 44092
rect 19356 44036 19360 44092
rect 19296 44032 19360 44036
rect 19376 44092 19440 44096
rect 19376 44036 19380 44092
rect 19380 44036 19436 44092
rect 19436 44036 19440 44092
rect 19376 44032 19440 44036
rect 19456 44092 19520 44096
rect 19456 44036 19460 44092
rect 19460 44036 19516 44092
rect 19516 44036 19520 44092
rect 19456 44032 19520 44036
rect 29216 44092 29280 44096
rect 29216 44036 29220 44092
rect 29220 44036 29276 44092
rect 29276 44036 29280 44092
rect 29216 44032 29280 44036
rect 29296 44092 29360 44096
rect 29296 44036 29300 44092
rect 29300 44036 29356 44092
rect 29356 44036 29360 44092
rect 29296 44032 29360 44036
rect 29376 44092 29440 44096
rect 29376 44036 29380 44092
rect 29380 44036 29436 44092
rect 29436 44036 29440 44092
rect 29376 44032 29440 44036
rect 29456 44092 29520 44096
rect 29456 44036 29460 44092
rect 29460 44036 29516 44092
rect 29516 44036 29520 44092
rect 29456 44032 29520 44036
rect 39216 44092 39280 44096
rect 39216 44036 39220 44092
rect 39220 44036 39276 44092
rect 39276 44036 39280 44092
rect 39216 44032 39280 44036
rect 39296 44092 39360 44096
rect 39296 44036 39300 44092
rect 39300 44036 39356 44092
rect 39356 44036 39360 44092
rect 39296 44032 39360 44036
rect 39376 44092 39440 44096
rect 39376 44036 39380 44092
rect 39380 44036 39436 44092
rect 39436 44036 39440 44092
rect 39376 44032 39440 44036
rect 39456 44092 39520 44096
rect 39456 44036 39460 44092
rect 39460 44036 39516 44092
rect 39516 44036 39520 44092
rect 39456 44032 39520 44036
rect 49216 44092 49280 44096
rect 49216 44036 49220 44092
rect 49220 44036 49276 44092
rect 49276 44036 49280 44092
rect 49216 44032 49280 44036
rect 49296 44092 49360 44096
rect 49296 44036 49300 44092
rect 49300 44036 49356 44092
rect 49356 44036 49360 44092
rect 49296 44032 49360 44036
rect 49376 44092 49440 44096
rect 49376 44036 49380 44092
rect 49380 44036 49436 44092
rect 49436 44036 49440 44092
rect 49376 44032 49440 44036
rect 49456 44092 49520 44096
rect 49456 44036 49460 44092
rect 49460 44036 49516 44092
rect 49516 44036 49520 44092
rect 49456 44032 49520 44036
rect 59216 44092 59280 44096
rect 59216 44036 59220 44092
rect 59220 44036 59276 44092
rect 59276 44036 59280 44092
rect 59216 44032 59280 44036
rect 59296 44092 59360 44096
rect 59296 44036 59300 44092
rect 59300 44036 59356 44092
rect 59356 44036 59360 44092
rect 59296 44032 59360 44036
rect 59376 44092 59440 44096
rect 59376 44036 59380 44092
rect 59380 44036 59436 44092
rect 59436 44036 59440 44092
rect 59376 44032 59440 44036
rect 59456 44092 59520 44096
rect 59456 44036 59460 44092
rect 59460 44036 59516 44092
rect 59516 44036 59520 44092
rect 59456 44032 59520 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 14216 43548 14280 43552
rect 14216 43492 14220 43548
rect 14220 43492 14276 43548
rect 14276 43492 14280 43548
rect 14216 43488 14280 43492
rect 14296 43548 14360 43552
rect 14296 43492 14300 43548
rect 14300 43492 14356 43548
rect 14356 43492 14360 43548
rect 14296 43488 14360 43492
rect 14376 43548 14440 43552
rect 14376 43492 14380 43548
rect 14380 43492 14436 43548
rect 14436 43492 14440 43548
rect 14376 43488 14440 43492
rect 14456 43548 14520 43552
rect 14456 43492 14460 43548
rect 14460 43492 14516 43548
rect 14516 43492 14520 43548
rect 14456 43488 14520 43492
rect 24216 43548 24280 43552
rect 24216 43492 24220 43548
rect 24220 43492 24276 43548
rect 24276 43492 24280 43548
rect 24216 43488 24280 43492
rect 24296 43548 24360 43552
rect 24296 43492 24300 43548
rect 24300 43492 24356 43548
rect 24356 43492 24360 43548
rect 24296 43488 24360 43492
rect 24376 43548 24440 43552
rect 24376 43492 24380 43548
rect 24380 43492 24436 43548
rect 24436 43492 24440 43548
rect 24376 43488 24440 43492
rect 24456 43548 24520 43552
rect 24456 43492 24460 43548
rect 24460 43492 24516 43548
rect 24516 43492 24520 43548
rect 24456 43488 24520 43492
rect 34216 43548 34280 43552
rect 34216 43492 34220 43548
rect 34220 43492 34276 43548
rect 34276 43492 34280 43548
rect 34216 43488 34280 43492
rect 34296 43548 34360 43552
rect 34296 43492 34300 43548
rect 34300 43492 34356 43548
rect 34356 43492 34360 43548
rect 34296 43488 34360 43492
rect 34376 43548 34440 43552
rect 34376 43492 34380 43548
rect 34380 43492 34436 43548
rect 34436 43492 34440 43548
rect 34376 43488 34440 43492
rect 34456 43548 34520 43552
rect 34456 43492 34460 43548
rect 34460 43492 34516 43548
rect 34516 43492 34520 43548
rect 34456 43488 34520 43492
rect 44216 43548 44280 43552
rect 44216 43492 44220 43548
rect 44220 43492 44276 43548
rect 44276 43492 44280 43548
rect 44216 43488 44280 43492
rect 44296 43548 44360 43552
rect 44296 43492 44300 43548
rect 44300 43492 44356 43548
rect 44356 43492 44360 43548
rect 44296 43488 44360 43492
rect 44376 43548 44440 43552
rect 44376 43492 44380 43548
rect 44380 43492 44436 43548
rect 44436 43492 44440 43548
rect 44376 43488 44440 43492
rect 44456 43548 44520 43552
rect 44456 43492 44460 43548
rect 44460 43492 44516 43548
rect 44516 43492 44520 43548
rect 44456 43488 44520 43492
rect 54216 43548 54280 43552
rect 54216 43492 54220 43548
rect 54220 43492 54276 43548
rect 54276 43492 54280 43548
rect 54216 43488 54280 43492
rect 54296 43548 54360 43552
rect 54296 43492 54300 43548
rect 54300 43492 54356 43548
rect 54356 43492 54360 43548
rect 54296 43488 54360 43492
rect 54376 43548 54440 43552
rect 54376 43492 54380 43548
rect 54380 43492 54436 43548
rect 54436 43492 54440 43548
rect 54376 43488 54440 43492
rect 54456 43548 54520 43552
rect 54456 43492 54460 43548
rect 54460 43492 54516 43548
rect 54516 43492 54520 43548
rect 54456 43488 54520 43492
rect 64216 43548 64280 43552
rect 64216 43492 64220 43548
rect 64220 43492 64276 43548
rect 64276 43492 64280 43548
rect 64216 43488 64280 43492
rect 64296 43548 64360 43552
rect 64296 43492 64300 43548
rect 64300 43492 64356 43548
rect 64356 43492 64360 43548
rect 64296 43488 64360 43492
rect 64376 43548 64440 43552
rect 64376 43492 64380 43548
rect 64380 43492 64436 43548
rect 64436 43492 64440 43548
rect 64376 43488 64440 43492
rect 64456 43548 64520 43552
rect 64456 43492 64460 43548
rect 64460 43492 64516 43548
rect 64516 43492 64520 43548
rect 64456 43488 64520 43492
rect 9216 43004 9280 43008
rect 9216 42948 9220 43004
rect 9220 42948 9276 43004
rect 9276 42948 9280 43004
rect 9216 42944 9280 42948
rect 9296 43004 9360 43008
rect 9296 42948 9300 43004
rect 9300 42948 9356 43004
rect 9356 42948 9360 43004
rect 9296 42944 9360 42948
rect 9376 43004 9440 43008
rect 9376 42948 9380 43004
rect 9380 42948 9436 43004
rect 9436 42948 9440 43004
rect 9376 42944 9440 42948
rect 9456 43004 9520 43008
rect 9456 42948 9460 43004
rect 9460 42948 9516 43004
rect 9516 42948 9520 43004
rect 9456 42944 9520 42948
rect 19216 43004 19280 43008
rect 19216 42948 19220 43004
rect 19220 42948 19276 43004
rect 19276 42948 19280 43004
rect 19216 42944 19280 42948
rect 19296 43004 19360 43008
rect 19296 42948 19300 43004
rect 19300 42948 19356 43004
rect 19356 42948 19360 43004
rect 19296 42944 19360 42948
rect 19376 43004 19440 43008
rect 19376 42948 19380 43004
rect 19380 42948 19436 43004
rect 19436 42948 19440 43004
rect 19376 42944 19440 42948
rect 19456 43004 19520 43008
rect 19456 42948 19460 43004
rect 19460 42948 19516 43004
rect 19516 42948 19520 43004
rect 19456 42944 19520 42948
rect 29216 43004 29280 43008
rect 29216 42948 29220 43004
rect 29220 42948 29276 43004
rect 29276 42948 29280 43004
rect 29216 42944 29280 42948
rect 29296 43004 29360 43008
rect 29296 42948 29300 43004
rect 29300 42948 29356 43004
rect 29356 42948 29360 43004
rect 29296 42944 29360 42948
rect 29376 43004 29440 43008
rect 29376 42948 29380 43004
rect 29380 42948 29436 43004
rect 29436 42948 29440 43004
rect 29376 42944 29440 42948
rect 29456 43004 29520 43008
rect 29456 42948 29460 43004
rect 29460 42948 29516 43004
rect 29516 42948 29520 43004
rect 29456 42944 29520 42948
rect 39216 43004 39280 43008
rect 39216 42948 39220 43004
rect 39220 42948 39276 43004
rect 39276 42948 39280 43004
rect 39216 42944 39280 42948
rect 39296 43004 39360 43008
rect 39296 42948 39300 43004
rect 39300 42948 39356 43004
rect 39356 42948 39360 43004
rect 39296 42944 39360 42948
rect 39376 43004 39440 43008
rect 39376 42948 39380 43004
rect 39380 42948 39436 43004
rect 39436 42948 39440 43004
rect 39376 42944 39440 42948
rect 39456 43004 39520 43008
rect 39456 42948 39460 43004
rect 39460 42948 39516 43004
rect 39516 42948 39520 43004
rect 39456 42944 39520 42948
rect 49216 43004 49280 43008
rect 49216 42948 49220 43004
rect 49220 42948 49276 43004
rect 49276 42948 49280 43004
rect 49216 42944 49280 42948
rect 49296 43004 49360 43008
rect 49296 42948 49300 43004
rect 49300 42948 49356 43004
rect 49356 42948 49360 43004
rect 49296 42944 49360 42948
rect 49376 43004 49440 43008
rect 49376 42948 49380 43004
rect 49380 42948 49436 43004
rect 49436 42948 49440 43004
rect 49376 42944 49440 42948
rect 49456 43004 49520 43008
rect 49456 42948 49460 43004
rect 49460 42948 49516 43004
rect 49516 42948 49520 43004
rect 49456 42944 49520 42948
rect 59216 43004 59280 43008
rect 59216 42948 59220 43004
rect 59220 42948 59276 43004
rect 59276 42948 59280 43004
rect 59216 42944 59280 42948
rect 59296 43004 59360 43008
rect 59296 42948 59300 43004
rect 59300 42948 59356 43004
rect 59356 42948 59360 43004
rect 59296 42944 59360 42948
rect 59376 43004 59440 43008
rect 59376 42948 59380 43004
rect 59380 42948 59436 43004
rect 59436 42948 59440 43004
rect 59376 42944 59440 42948
rect 59456 43004 59520 43008
rect 59456 42948 59460 43004
rect 59460 42948 59516 43004
rect 59516 42948 59520 43004
rect 59456 42944 59520 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 14216 42460 14280 42464
rect 14216 42404 14220 42460
rect 14220 42404 14276 42460
rect 14276 42404 14280 42460
rect 14216 42400 14280 42404
rect 14296 42460 14360 42464
rect 14296 42404 14300 42460
rect 14300 42404 14356 42460
rect 14356 42404 14360 42460
rect 14296 42400 14360 42404
rect 14376 42460 14440 42464
rect 14376 42404 14380 42460
rect 14380 42404 14436 42460
rect 14436 42404 14440 42460
rect 14376 42400 14440 42404
rect 14456 42460 14520 42464
rect 14456 42404 14460 42460
rect 14460 42404 14516 42460
rect 14516 42404 14520 42460
rect 14456 42400 14520 42404
rect 24216 42460 24280 42464
rect 24216 42404 24220 42460
rect 24220 42404 24276 42460
rect 24276 42404 24280 42460
rect 24216 42400 24280 42404
rect 24296 42460 24360 42464
rect 24296 42404 24300 42460
rect 24300 42404 24356 42460
rect 24356 42404 24360 42460
rect 24296 42400 24360 42404
rect 24376 42460 24440 42464
rect 24376 42404 24380 42460
rect 24380 42404 24436 42460
rect 24436 42404 24440 42460
rect 24376 42400 24440 42404
rect 24456 42460 24520 42464
rect 24456 42404 24460 42460
rect 24460 42404 24516 42460
rect 24516 42404 24520 42460
rect 24456 42400 24520 42404
rect 34216 42460 34280 42464
rect 34216 42404 34220 42460
rect 34220 42404 34276 42460
rect 34276 42404 34280 42460
rect 34216 42400 34280 42404
rect 34296 42460 34360 42464
rect 34296 42404 34300 42460
rect 34300 42404 34356 42460
rect 34356 42404 34360 42460
rect 34296 42400 34360 42404
rect 34376 42460 34440 42464
rect 34376 42404 34380 42460
rect 34380 42404 34436 42460
rect 34436 42404 34440 42460
rect 34376 42400 34440 42404
rect 34456 42460 34520 42464
rect 34456 42404 34460 42460
rect 34460 42404 34516 42460
rect 34516 42404 34520 42460
rect 34456 42400 34520 42404
rect 44216 42460 44280 42464
rect 44216 42404 44220 42460
rect 44220 42404 44276 42460
rect 44276 42404 44280 42460
rect 44216 42400 44280 42404
rect 44296 42460 44360 42464
rect 44296 42404 44300 42460
rect 44300 42404 44356 42460
rect 44356 42404 44360 42460
rect 44296 42400 44360 42404
rect 44376 42460 44440 42464
rect 44376 42404 44380 42460
rect 44380 42404 44436 42460
rect 44436 42404 44440 42460
rect 44376 42400 44440 42404
rect 44456 42460 44520 42464
rect 44456 42404 44460 42460
rect 44460 42404 44516 42460
rect 44516 42404 44520 42460
rect 44456 42400 44520 42404
rect 54216 42460 54280 42464
rect 54216 42404 54220 42460
rect 54220 42404 54276 42460
rect 54276 42404 54280 42460
rect 54216 42400 54280 42404
rect 54296 42460 54360 42464
rect 54296 42404 54300 42460
rect 54300 42404 54356 42460
rect 54356 42404 54360 42460
rect 54296 42400 54360 42404
rect 54376 42460 54440 42464
rect 54376 42404 54380 42460
rect 54380 42404 54436 42460
rect 54436 42404 54440 42460
rect 54376 42400 54440 42404
rect 54456 42460 54520 42464
rect 54456 42404 54460 42460
rect 54460 42404 54516 42460
rect 54516 42404 54520 42460
rect 54456 42400 54520 42404
rect 64216 42460 64280 42464
rect 64216 42404 64220 42460
rect 64220 42404 64276 42460
rect 64276 42404 64280 42460
rect 64216 42400 64280 42404
rect 64296 42460 64360 42464
rect 64296 42404 64300 42460
rect 64300 42404 64356 42460
rect 64356 42404 64360 42460
rect 64296 42400 64360 42404
rect 64376 42460 64440 42464
rect 64376 42404 64380 42460
rect 64380 42404 64436 42460
rect 64436 42404 64440 42460
rect 64376 42400 64440 42404
rect 64456 42460 64520 42464
rect 64456 42404 64460 42460
rect 64460 42404 64516 42460
rect 64516 42404 64520 42460
rect 64456 42400 64520 42404
rect 9216 41916 9280 41920
rect 9216 41860 9220 41916
rect 9220 41860 9276 41916
rect 9276 41860 9280 41916
rect 9216 41856 9280 41860
rect 9296 41916 9360 41920
rect 9296 41860 9300 41916
rect 9300 41860 9356 41916
rect 9356 41860 9360 41916
rect 9296 41856 9360 41860
rect 9376 41916 9440 41920
rect 9376 41860 9380 41916
rect 9380 41860 9436 41916
rect 9436 41860 9440 41916
rect 9376 41856 9440 41860
rect 9456 41916 9520 41920
rect 9456 41860 9460 41916
rect 9460 41860 9516 41916
rect 9516 41860 9520 41916
rect 9456 41856 9520 41860
rect 19216 41916 19280 41920
rect 19216 41860 19220 41916
rect 19220 41860 19276 41916
rect 19276 41860 19280 41916
rect 19216 41856 19280 41860
rect 19296 41916 19360 41920
rect 19296 41860 19300 41916
rect 19300 41860 19356 41916
rect 19356 41860 19360 41916
rect 19296 41856 19360 41860
rect 19376 41916 19440 41920
rect 19376 41860 19380 41916
rect 19380 41860 19436 41916
rect 19436 41860 19440 41916
rect 19376 41856 19440 41860
rect 19456 41916 19520 41920
rect 19456 41860 19460 41916
rect 19460 41860 19516 41916
rect 19516 41860 19520 41916
rect 19456 41856 19520 41860
rect 29216 41916 29280 41920
rect 29216 41860 29220 41916
rect 29220 41860 29276 41916
rect 29276 41860 29280 41916
rect 29216 41856 29280 41860
rect 29296 41916 29360 41920
rect 29296 41860 29300 41916
rect 29300 41860 29356 41916
rect 29356 41860 29360 41916
rect 29296 41856 29360 41860
rect 29376 41916 29440 41920
rect 29376 41860 29380 41916
rect 29380 41860 29436 41916
rect 29436 41860 29440 41916
rect 29376 41856 29440 41860
rect 29456 41916 29520 41920
rect 29456 41860 29460 41916
rect 29460 41860 29516 41916
rect 29516 41860 29520 41916
rect 29456 41856 29520 41860
rect 39216 41916 39280 41920
rect 39216 41860 39220 41916
rect 39220 41860 39276 41916
rect 39276 41860 39280 41916
rect 39216 41856 39280 41860
rect 39296 41916 39360 41920
rect 39296 41860 39300 41916
rect 39300 41860 39356 41916
rect 39356 41860 39360 41916
rect 39296 41856 39360 41860
rect 39376 41916 39440 41920
rect 39376 41860 39380 41916
rect 39380 41860 39436 41916
rect 39436 41860 39440 41916
rect 39376 41856 39440 41860
rect 39456 41916 39520 41920
rect 39456 41860 39460 41916
rect 39460 41860 39516 41916
rect 39516 41860 39520 41916
rect 39456 41856 39520 41860
rect 49216 41916 49280 41920
rect 49216 41860 49220 41916
rect 49220 41860 49276 41916
rect 49276 41860 49280 41916
rect 49216 41856 49280 41860
rect 49296 41916 49360 41920
rect 49296 41860 49300 41916
rect 49300 41860 49356 41916
rect 49356 41860 49360 41916
rect 49296 41856 49360 41860
rect 49376 41916 49440 41920
rect 49376 41860 49380 41916
rect 49380 41860 49436 41916
rect 49436 41860 49440 41916
rect 49376 41856 49440 41860
rect 49456 41916 49520 41920
rect 49456 41860 49460 41916
rect 49460 41860 49516 41916
rect 49516 41860 49520 41916
rect 49456 41856 49520 41860
rect 59216 41916 59280 41920
rect 59216 41860 59220 41916
rect 59220 41860 59276 41916
rect 59276 41860 59280 41916
rect 59216 41856 59280 41860
rect 59296 41916 59360 41920
rect 59296 41860 59300 41916
rect 59300 41860 59356 41916
rect 59356 41860 59360 41916
rect 59296 41856 59360 41860
rect 59376 41916 59440 41920
rect 59376 41860 59380 41916
rect 59380 41860 59436 41916
rect 59436 41860 59440 41916
rect 59376 41856 59440 41860
rect 59456 41916 59520 41920
rect 59456 41860 59460 41916
rect 59460 41860 59516 41916
rect 59516 41860 59520 41916
rect 59456 41856 59520 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 14216 41372 14280 41376
rect 14216 41316 14220 41372
rect 14220 41316 14276 41372
rect 14276 41316 14280 41372
rect 14216 41312 14280 41316
rect 14296 41372 14360 41376
rect 14296 41316 14300 41372
rect 14300 41316 14356 41372
rect 14356 41316 14360 41372
rect 14296 41312 14360 41316
rect 14376 41372 14440 41376
rect 14376 41316 14380 41372
rect 14380 41316 14436 41372
rect 14436 41316 14440 41372
rect 14376 41312 14440 41316
rect 14456 41372 14520 41376
rect 14456 41316 14460 41372
rect 14460 41316 14516 41372
rect 14516 41316 14520 41372
rect 14456 41312 14520 41316
rect 24216 41372 24280 41376
rect 24216 41316 24220 41372
rect 24220 41316 24276 41372
rect 24276 41316 24280 41372
rect 24216 41312 24280 41316
rect 24296 41372 24360 41376
rect 24296 41316 24300 41372
rect 24300 41316 24356 41372
rect 24356 41316 24360 41372
rect 24296 41312 24360 41316
rect 24376 41372 24440 41376
rect 24376 41316 24380 41372
rect 24380 41316 24436 41372
rect 24436 41316 24440 41372
rect 24376 41312 24440 41316
rect 24456 41372 24520 41376
rect 24456 41316 24460 41372
rect 24460 41316 24516 41372
rect 24516 41316 24520 41372
rect 24456 41312 24520 41316
rect 34216 41372 34280 41376
rect 34216 41316 34220 41372
rect 34220 41316 34276 41372
rect 34276 41316 34280 41372
rect 34216 41312 34280 41316
rect 34296 41372 34360 41376
rect 34296 41316 34300 41372
rect 34300 41316 34356 41372
rect 34356 41316 34360 41372
rect 34296 41312 34360 41316
rect 34376 41372 34440 41376
rect 34376 41316 34380 41372
rect 34380 41316 34436 41372
rect 34436 41316 34440 41372
rect 34376 41312 34440 41316
rect 34456 41372 34520 41376
rect 34456 41316 34460 41372
rect 34460 41316 34516 41372
rect 34516 41316 34520 41372
rect 34456 41312 34520 41316
rect 44216 41372 44280 41376
rect 44216 41316 44220 41372
rect 44220 41316 44276 41372
rect 44276 41316 44280 41372
rect 44216 41312 44280 41316
rect 44296 41372 44360 41376
rect 44296 41316 44300 41372
rect 44300 41316 44356 41372
rect 44356 41316 44360 41372
rect 44296 41312 44360 41316
rect 44376 41372 44440 41376
rect 44376 41316 44380 41372
rect 44380 41316 44436 41372
rect 44436 41316 44440 41372
rect 44376 41312 44440 41316
rect 44456 41372 44520 41376
rect 44456 41316 44460 41372
rect 44460 41316 44516 41372
rect 44516 41316 44520 41372
rect 44456 41312 44520 41316
rect 54216 41372 54280 41376
rect 54216 41316 54220 41372
rect 54220 41316 54276 41372
rect 54276 41316 54280 41372
rect 54216 41312 54280 41316
rect 54296 41372 54360 41376
rect 54296 41316 54300 41372
rect 54300 41316 54356 41372
rect 54356 41316 54360 41372
rect 54296 41312 54360 41316
rect 54376 41372 54440 41376
rect 54376 41316 54380 41372
rect 54380 41316 54436 41372
rect 54436 41316 54440 41372
rect 54376 41312 54440 41316
rect 54456 41372 54520 41376
rect 54456 41316 54460 41372
rect 54460 41316 54516 41372
rect 54516 41316 54520 41372
rect 54456 41312 54520 41316
rect 64216 41372 64280 41376
rect 64216 41316 64220 41372
rect 64220 41316 64276 41372
rect 64276 41316 64280 41372
rect 64216 41312 64280 41316
rect 64296 41372 64360 41376
rect 64296 41316 64300 41372
rect 64300 41316 64356 41372
rect 64356 41316 64360 41372
rect 64296 41312 64360 41316
rect 64376 41372 64440 41376
rect 64376 41316 64380 41372
rect 64380 41316 64436 41372
rect 64436 41316 64440 41372
rect 64376 41312 64440 41316
rect 64456 41372 64520 41376
rect 64456 41316 64460 41372
rect 64460 41316 64516 41372
rect 64516 41316 64520 41372
rect 64456 41312 64520 41316
rect 9216 40828 9280 40832
rect 9216 40772 9220 40828
rect 9220 40772 9276 40828
rect 9276 40772 9280 40828
rect 9216 40768 9280 40772
rect 9296 40828 9360 40832
rect 9296 40772 9300 40828
rect 9300 40772 9356 40828
rect 9356 40772 9360 40828
rect 9296 40768 9360 40772
rect 9376 40828 9440 40832
rect 9376 40772 9380 40828
rect 9380 40772 9436 40828
rect 9436 40772 9440 40828
rect 9376 40768 9440 40772
rect 9456 40828 9520 40832
rect 9456 40772 9460 40828
rect 9460 40772 9516 40828
rect 9516 40772 9520 40828
rect 9456 40768 9520 40772
rect 19216 40828 19280 40832
rect 19216 40772 19220 40828
rect 19220 40772 19276 40828
rect 19276 40772 19280 40828
rect 19216 40768 19280 40772
rect 19296 40828 19360 40832
rect 19296 40772 19300 40828
rect 19300 40772 19356 40828
rect 19356 40772 19360 40828
rect 19296 40768 19360 40772
rect 19376 40828 19440 40832
rect 19376 40772 19380 40828
rect 19380 40772 19436 40828
rect 19436 40772 19440 40828
rect 19376 40768 19440 40772
rect 19456 40828 19520 40832
rect 19456 40772 19460 40828
rect 19460 40772 19516 40828
rect 19516 40772 19520 40828
rect 19456 40768 19520 40772
rect 29216 40828 29280 40832
rect 29216 40772 29220 40828
rect 29220 40772 29276 40828
rect 29276 40772 29280 40828
rect 29216 40768 29280 40772
rect 29296 40828 29360 40832
rect 29296 40772 29300 40828
rect 29300 40772 29356 40828
rect 29356 40772 29360 40828
rect 29296 40768 29360 40772
rect 29376 40828 29440 40832
rect 29376 40772 29380 40828
rect 29380 40772 29436 40828
rect 29436 40772 29440 40828
rect 29376 40768 29440 40772
rect 29456 40828 29520 40832
rect 29456 40772 29460 40828
rect 29460 40772 29516 40828
rect 29516 40772 29520 40828
rect 29456 40768 29520 40772
rect 39216 40828 39280 40832
rect 39216 40772 39220 40828
rect 39220 40772 39276 40828
rect 39276 40772 39280 40828
rect 39216 40768 39280 40772
rect 39296 40828 39360 40832
rect 39296 40772 39300 40828
rect 39300 40772 39356 40828
rect 39356 40772 39360 40828
rect 39296 40768 39360 40772
rect 39376 40828 39440 40832
rect 39376 40772 39380 40828
rect 39380 40772 39436 40828
rect 39436 40772 39440 40828
rect 39376 40768 39440 40772
rect 39456 40828 39520 40832
rect 39456 40772 39460 40828
rect 39460 40772 39516 40828
rect 39516 40772 39520 40828
rect 39456 40768 39520 40772
rect 49216 40828 49280 40832
rect 49216 40772 49220 40828
rect 49220 40772 49276 40828
rect 49276 40772 49280 40828
rect 49216 40768 49280 40772
rect 49296 40828 49360 40832
rect 49296 40772 49300 40828
rect 49300 40772 49356 40828
rect 49356 40772 49360 40828
rect 49296 40768 49360 40772
rect 49376 40828 49440 40832
rect 49376 40772 49380 40828
rect 49380 40772 49436 40828
rect 49436 40772 49440 40828
rect 49376 40768 49440 40772
rect 49456 40828 49520 40832
rect 49456 40772 49460 40828
rect 49460 40772 49516 40828
rect 49516 40772 49520 40828
rect 49456 40768 49520 40772
rect 59216 40828 59280 40832
rect 59216 40772 59220 40828
rect 59220 40772 59276 40828
rect 59276 40772 59280 40828
rect 59216 40768 59280 40772
rect 59296 40828 59360 40832
rect 59296 40772 59300 40828
rect 59300 40772 59356 40828
rect 59356 40772 59360 40828
rect 59296 40768 59360 40772
rect 59376 40828 59440 40832
rect 59376 40772 59380 40828
rect 59380 40772 59436 40828
rect 59436 40772 59440 40828
rect 59376 40768 59440 40772
rect 59456 40828 59520 40832
rect 59456 40772 59460 40828
rect 59460 40772 59516 40828
rect 59516 40772 59520 40828
rect 59456 40768 59520 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 14216 40284 14280 40288
rect 14216 40228 14220 40284
rect 14220 40228 14276 40284
rect 14276 40228 14280 40284
rect 14216 40224 14280 40228
rect 14296 40284 14360 40288
rect 14296 40228 14300 40284
rect 14300 40228 14356 40284
rect 14356 40228 14360 40284
rect 14296 40224 14360 40228
rect 14376 40284 14440 40288
rect 14376 40228 14380 40284
rect 14380 40228 14436 40284
rect 14436 40228 14440 40284
rect 14376 40224 14440 40228
rect 14456 40284 14520 40288
rect 14456 40228 14460 40284
rect 14460 40228 14516 40284
rect 14516 40228 14520 40284
rect 14456 40224 14520 40228
rect 24216 40284 24280 40288
rect 24216 40228 24220 40284
rect 24220 40228 24276 40284
rect 24276 40228 24280 40284
rect 24216 40224 24280 40228
rect 24296 40284 24360 40288
rect 24296 40228 24300 40284
rect 24300 40228 24356 40284
rect 24356 40228 24360 40284
rect 24296 40224 24360 40228
rect 24376 40284 24440 40288
rect 24376 40228 24380 40284
rect 24380 40228 24436 40284
rect 24436 40228 24440 40284
rect 24376 40224 24440 40228
rect 24456 40284 24520 40288
rect 24456 40228 24460 40284
rect 24460 40228 24516 40284
rect 24516 40228 24520 40284
rect 24456 40224 24520 40228
rect 34216 40284 34280 40288
rect 34216 40228 34220 40284
rect 34220 40228 34276 40284
rect 34276 40228 34280 40284
rect 34216 40224 34280 40228
rect 34296 40284 34360 40288
rect 34296 40228 34300 40284
rect 34300 40228 34356 40284
rect 34356 40228 34360 40284
rect 34296 40224 34360 40228
rect 34376 40284 34440 40288
rect 34376 40228 34380 40284
rect 34380 40228 34436 40284
rect 34436 40228 34440 40284
rect 34376 40224 34440 40228
rect 34456 40284 34520 40288
rect 34456 40228 34460 40284
rect 34460 40228 34516 40284
rect 34516 40228 34520 40284
rect 34456 40224 34520 40228
rect 44216 40284 44280 40288
rect 44216 40228 44220 40284
rect 44220 40228 44276 40284
rect 44276 40228 44280 40284
rect 44216 40224 44280 40228
rect 44296 40284 44360 40288
rect 44296 40228 44300 40284
rect 44300 40228 44356 40284
rect 44356 40228 44360 40284
rect 44296 40224 44360 40228
rect 44376 40284 44440 40288
rect 44376 40228 44380 40284
rect 44380 40228 44436 40284
rect 44436 40228 44440 40284
rect 44376 40224 44440 40228
rect 44456 40284 44520 40288
rect 44456 40228 44460 40284
rect 44460 40228 44516 40284
rect 44516 40228 44520 40284
rect 44456 40224 44520 40228
rect 54216 40284 54280 40288
rect 54216 40228 54220 40284
rect 54220 40228 54276 40284
rect 54276 40228 54280 40284
rect 54216 40224 54280 40228
rect 54296 40284 54360 40288
rect 54296 40228 54300 40284
rect 54300 40228 54356 40284
rect 54356 40228 54360 40284
rect 54296 40224 54360 40228
rect 54376 40284 54440 40288
rect 54376 40228 54380 40284
rect 54380 40228 54436 40284
rect 54436 40228 54440 40284
rect 54376 40224 54440 40228
rect 54456 40284 54520 40288
rect 54456 40228 54460 40284
rect 54460 40228 54516 40284
rect 54516 40228 54520 40284
rect 54456 40224 54520 40228
rect 64216 40284 64280 40288
rect 64216 40228 64220 40284
rect 64220 40228 64276 40284
rect 64276 40228 64280 40284
rect 64216 40224 64280 40228
rect 64296 40284 64360 40288
rect 64296 40228 64300 40284
rect 64300 40228 64356 40284
rect 64356 40228 64360 40284
rect 64296 40224 64360 40228
rect 64376 40284 64440 40288
rect 64376 40228 64380 40284
rect 64380 40228 64436 40284
rect 64436 40228 64440 40284
rect 64376 40224 64440 40228
rect 64456 40284 64520 40288
rect 64456 40228 64460 40284
rect 64460 40228 64516 40284
rect 64516 40228 64520 40284
rect 64456 40224 64520 40228
rect 9216 39740 9280 39744
rect 9216 39684 9220 39740
rect 9220 39684 9276 39740
rect 9276 39684 9280 39740
rect 9216 39680 9280 39684
rect 9296 39740 9360 39744
rect 9296 39684 9300 39740
rect 9300 39684 9356 39740
rect 9356 39684 9360 39740
rect 9296 39680 9360 39684
rect 9376 39740 9440 39744
rect 9376 39684 9380 39740
rect 9380 39684 9436 39740
rect 9436 39684 9440 39740
rect 9376 39680 9440 39684
rect 9456 39740 9520 39744
rect 9456 39684 9460 39740
rect 9460 39684 9516 39740
rect 9516 39684 9520 39740
rect 9456 39680 9520 39684
rect 19216 39740 19280 39744
rect 19216 39684 19220 39740
rect 19220 39684 19276 39740
rect 19276 39684 19280 39740
rect 19216 39680 19280 39684
rect 19296 39740 19360 39744
rect 19296 39684 19300 39740
rect 19300 39684 19356 39740
rect 19356 39684 19360 39740
rect 19296 39680 19360 39684
rect 19376 39740 19440 39744
rect 19376 39684 19380 39740
rect 19380 39684 19436 39740
rect 19436 39684 19440 39740
rect 19376 39680 19440 39684
rect 19456 39740 19520 39744
rect 19456 39684 19460 39740
rect 19460 39684 19516 39740
rect 19516 39684 19520 39740
rect 19456 39680 19520 39684
rect 29216 39740 29280 39744
rect 29216 39684 29220 39740
rect 29220 39684 29276 39740
rect 29276 39684 29280 39740
rect 29216 39680 29280 39684
rect 29296 39740 29360 39744
rect 29296 39684 29300 39740
rect 29300 39684 29356 39740
rect 29356 39684 29360 39740
rect 29296 39680 29360 39684
rect 29376 39740 29440 39744
rect 29376 39684 29380 39740
rect 29380 39684 29436 39740
rect 29436 39684 29440 39740
rect 29376 39680 29440 39684
rect 29456 39740 29520 39744
rect 29456 39684 29460 39740
rect 29460 39684 29516 39740
rect 29516 39684 29520 39740
rect 29456 39680 29520 39684
rect 39216 39740 39280 39744
rect 39216 39684 39220 39740
rect 39220 39684 39276 39740
rect 39276 39684 39280 39740
rect 39216 39680 39280 39684
rect 39296 39740 39360 39744
rect 39296 39684 39300 39740
rect 39300 39684 39356 39740
rect 39356 39684 39360 39740
rect 39296 39680 39360 39684
rect 39376 39740 39440 39744
rect 39376 39684 39380 39740
rect 39380 39684 39436 39740
rect 39436 39684 39440 39740
rect 39376 39680 39440 39684
rect 39456 39740 39520 39744
rect 39456 39684 39460 39740
rect 39460 39684 39516 39740
rect 39516 39684 39520 39740
rect 39456 39680 39520 39684
rect 49216 39740 49280 39744
rect 49216 39684 49220 39740
rect 49220 39684 49276 39740
rect 49276 39684 49280 39740
rect 49216 39680 49280 39684
rect 49296 39740 49360 39744
rect 49296 39684 49300 39740
rect 49300 39684 49356 39740
rect 49356 39684 49360 39740
rect 49296 39680 49360 39684
rect 49376 39740 49440 39744
rect 49376 39684 49380 39740
rect 49380 39684 49436 39740
rect 49436 39684 49440 39740
rect 49376 39680 49440 39684
rect 49456 39740 49520 39744
rect 49456 39684 49460 39740
rect 49460 39684 49516 39740
rect 49516 39684 49520 39740
rect 49456 39680 49520 39684
rect 59216 39740 59280 39744
rect 59216 39684 59220 39740
rect 59220 39684 59276 39740
rect 59276 39684 59280 39740
rect 59216 39680 59280 39684
rect 59296 39740 59360 39744
rect 59296 39684 59300 39740
rect 59300 39684 59356 39740
rect 59356 39684 59360 39740
rect 59296 39680 59360 39684
rect 59376 39740 59440 39744
rect 59376 39684 59380 39740
rect 59380 39684 59436 39740
rect 59436 39684 59440 39740
rect 59376 39680 59440 39684
rect 59456 39740 59520 39744
rect 59456 39684 59460 39740
rect 59460 39684 59516 39740
rect 59516 39684 59520 39740
rect 59456 39680 59520 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 14216 39196 14280 39200
rect 14216 39140 14220 39196
rect 14220 39140 14276 39196
rect 14276 39140 14280 39196
rect 14216 39136 14280 39140
rect 14296 39196 14360 39200
rect 14296 39140 14300 39196
rect 14300 39140 14356 39196
rect 14356 39140 14360 39196
rect 14296 39136 14360 39140
rect 14376 39196 14440 39200
rect 14376 39140 14380 39196
rect 14380 39140 14436 39196
rect 14436 39140 14440 39196
rect 14376 39136 14440 39140
rect 14456 39196 14520 39200
rect 14456 39140 14460 39196
rect 14460 39140 14516 39196
rect 14516 39140 14520 39196
rect 14456 39136 14520 39140
rect 24216 39196 24280 39200
rect 24216 39140 24220 39196
rect 24220 39140 24276 39196
rect 24276 39140 24280 39196
rect 24216 39136 24280 39140
rect 24296 39196 24360 39200
rect 24296 39140 24300 39196
rect 24300 39140 24356 39196
rect 24356 39140 24360 39196
rect 24296 39136 24360 39140
rect 24376 39196 24440 39200
rect 24376 39140 24380 39196
rect 24380 39140 24436 39196
rect 24436 39140 24440 39196
rect 24376 39136 24440 39140
rect 24456 39196 24520 39200
rect 24456 39140 24460 39196
rect 24460 39140 24516 39196
rect 24516 39140 24520 39196
rect 24456 39136 24520 39140
rect 34216 39196 34280 39200
rect 34216 39140 34220 39196
rect 34220 39140 34276 39196
rect 34276 39140 34280 39196
rect 34216 39136 34280 39140
rect 34296 39196 34360 39200
rect 34296 39140 34300 39196
rect 34300 39140 34356 39196
rect 34356 39140 34360 39196
rect 34296 39136 34360 39140
rect 34376 39196 34440 39200
rect 34376 39140 34380 39196
rect 34380 39140 34436 39196
rect 34436 39140 34440 39196
rect 34376 39136 34440 39140
rect 34456 39196 34520 39200
rect 34456 39140 34460 39196
rect 34460 39140 34516 39196
rect 34516 39140 34520 39196
rect 34456 39136 34520 39140
rect 44216 39196 44280 39200
rect 44216 39140 44220 39196
rect 44220 39140 44276 39196
rect 44276 39140 44280 39196
rect 44216 39136 44280 39140
rect 44296 39196 44360 39200
rect 44296 39140 44300 39196
rect 44300 39140 44356 39196
rect 44356 39140 44360 39196
rect 44296 39136 44360 39140
rect 44376 39196 44440 39200
rect 44376 39140 44380 39196
rect 44380 39140 44436 39196
rect 44436 39140 44440 39196
rect 44376 39136 44440 39140
rect 44456 39196 44520 39200
rect 44456 39140 44460 39196
rect 44460 39140 44516 39196
rect 44516 39140 44520 39196
rect 44456 39136 44520 39140
rect 54216 39196 54280 39200
rect 54216 39140 54220 39196
rect 54220 39140 54276 39196
rect 54276 39140 54280 39196
rect 54216 39136 54280 39140
rect 54296 39196 54360 39200
rect 54296 39140 54300 39196
rect 54300 39140 54356 39196
rect 54356 39140 54360 39196
rect 54296 39136 54360 39140
rect 54376 39196 54440 39200
rect 54376 39140 54380 39196
rect 54380 39140 54436 39196
rect 54436 39140 54440 39196
rect 54376 39136 54440 39140
rect 54456 39196 54520 39200
rect 54456 39140 54460 39196
rect 54460 39140 54516 39196
rect 54516 39140 54520 39196
rect 54456 39136 54520 39140
rect 64216 39196 64280 39200
rect 64216 39140 64220 39196
rect 64220 39140 64276 39196
rect 64276 39140 64280 39196
rect 64216 39136 64280 39140
rect 64296 39196 64360 39200
rect 64296 39140 64300 39196
rect 64300 39140 64356 39196
rect 64356 39140 64360 39196
rect 64296 39136 64360 39140
rect 64376 39196 64440 39200
rect 64376 39140 64380 39196
rect 64380 39140 64436 39196
rect 64436 39140 64440 39196
rect 64376 39136 64440 39140
rect 64456 39196 64520 39200
rect 64456 39140 64460 39196
rect 64460 39140 64516 39196
rect 64516 39140 64520 39196
rect 64456 39136 64520 39140
rect 9216 38652 9280 38656
rect 9216 38596 9220 38652
rect 9220 38596 9276 38652
rect 9276 38596 9280 38652
rect 9216 38592 9280 38596
rect 9296 38652 9360 38656
rect 9296 38596 9300 38652
rect 9300 38596 9356 38652
rect 9356 38596 9360 38652
rect 9296 38592 9360 38596
rect 9376 38652 9440 38656
rect 9376 38596 9380 38652
rect 9380 38596 9436 38652
rect 9436 38596 9440 38652
rect 9376 38592 9440 38596
rect 9456 38652 9520 38656
rect 9456 38596 9460 38652
rect 9460 38596 9516 38652
rect 9516 38596 9520 38652
rect 9456 38592 9520 38596
rect 19216 38652 19280 38656
rect 19216 38596 19220 38652
rect 19220 38596 19276 38652
rect 19276 38596 19280 38652
rect 19216 38592 19280 38596
rect 19296 38652 19360 38656
rect 19296 38596 19300 38652
rect 19300 38596 19356 38652
rect 19356 38596 19360 38652
rect 19296 38592 19360 38596
rect 19376 38652 19440 38656
rect 19376 38596 19380 38652
rect 19380 38596 19436 38652
rect 19436 38596 19440 38652
rect 19376 38592 19440 38596
rect 19456 38652 19520 38656
rect 19456 38596 19460 38652
rect 19460 38596 19516 38652
rect 19516 38596 19520 38652
rect 19456 38592 19520 38596
rect 29216 38652 29280 38656
rect 29216 38596 29220 38652
rect 29220 38596 29276 38652
rect 29276 38596 29280 38652
rect 29216 38592 29280 38596
rect 29296 38652 29360 38656
rect 29296 38596 29300 38652
rect 29300 38596 29356 38652
rect 29356 38596 29360 38652
rect 29296 38592 29360 38596
rect 29376 38652 29440 38656
rect 29376 38596 29380 38652
rect 29380 38596 29436 38652
rect 29436 38596 29440 38652
rect 29376 38592 29440 38596
rect 29456 38652 29520 38656
rect 29456 38596 29460 38652
rect 29460 38596 29516 38652
rect 29516 38596 29520 38652
rect 29456 38592 29520 38596
rect 39216 38652 39280 38656
rect 39216 38596 39220 38652
rect 39220 38596 39276 38652
rect 39276 38596 39280 38652
rect 39216 38592 39280 38596
rect 39296 38652 39360 38656
rect 39296 38596 39300 38652
rect 39300 38596 39356 38652
rect 39356 38596 39360 38652
rect 39296 38592 39360 38596
rect 39376 38652 39440 38656
rect 39376 38596 39380 38652
rect 39380 38596 39436 38652
rect 39436 38596 39440 38652
rect 39376 38592 39440 38596
rect 39456 38652 39520 38656
rect 39456 38596 39460 38652
rect 39460 38596 39516 38652
rect 39516 38596 39520 38652
rect 39456 38592 39520 38596
rect 49216 38652 49280 38656
rect 49216 38596 49220 38652
rect 49220 38596 49276 38652
rect 49276 38596 49280 38652
rect 49216 38592 49280 38596
rect 49296 38652 49360 38656
rect 49296 38596 49300 38652
rect 49300 38596 49356 38652
rect 49356 38596 49360 38652
rect 49296 38592 49360 38596
rect 49376 38652 49440 38656
rect 49376 38596 49380 38652
rect 49380 38596 49436 38652
rect 49436 38596 49440 38652
rect 49376 38592 49440 38596
rect 49456 38652 49520 38656
rect 49456 38596 49460 38652
rect 49460 38596 49516 38652
rect 49516 38596 49520 38652
rect 49456 38592 49520 38596
rect 59216 38652 59280 38656
rect 59216 38596 59220 38652
rect 59220 38596 59276 38652
rect 59276 38596 59280 38652
rect 59216 38592 59280 38596
rect 59296 38652 59360 38656
rect 59296 38596 59300 38652
rect 59300 38596 59356 38652
rect 59356 38596 59360 38652
rect 59296 38592 59360 38596
rect 59376 38652 59440 38656
rect 59376 38596 59380 38652
rect 59380 38596 59436 38652
rect 59436 38596 59440 38652
rect 59376 38592 59440 38596
rect 59456 38652 59520 38656
rect 59456 38596 59460 38652
rect 59460 38596 59516 38652
rect 59516 38596 59520 38652
rect 59456 38592 59520 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 14216 38108 14280 38112
rect 14216 38052 14220 38108
rect 14220 38052 14276 38108
rect 14276 38052 14280 38108
rect 14216 38048 14280 38052
rect 14296 38108 14360 38112
rect 14296 38052 14300 38108
rect 14300 38052 14356 38108
rect 14356 38052 14360 38108
rect 14296 38048 14360 38052
rect 14376 38108 14440 38112
rect 14376 38052 14380 38108
rect 14380 38052 14436 38108
rect 14436 38052 14440 38108
rect 14376 38048 14440 38052
rect 14456 38108 14520 38112
rect 14456 38052 14460 38108
rect 14460 38052 14516 38108
rect 14516 38052 14520 38108
rect 14456 38048 14520 38052
rect 24216 38108 24280 38112
rect 24216 38052 24220 38108
rect 24220 38052 24276 38108
rect 24276 38052 24280 38108
rect 24216 38048 24280 38052
rect 24296 38108 24360 38112
rect 24296 38052 24300 38108
rect 24300 38052 24356 38108
rect 24356 38052 24360 38108
rect 24296 38048 24360 38052
rect 24376 38108 24440 38112
rect 24376 38052 24380 38108
rect 24380 38052 24436 38108
rect 24436 38052 24440 38108
rect 24376 38048 24440 38052
rect 24456 38108 24520 38112
rect 24456 38052 24460 38108
rect 24460 38052 24516 38108
rect 24516 38052 24520 38108
rect 24456 38048 24520 38052
rect 34216 38108 34280 38112
rect 34216 38052 34220 38108
rect 34220 38052 34276 38108
rect 34276 38052 34280 38108
rect 34216 38048 34280 38052
rect 34296 38108 34360 38112
rect 34296 38052 34300 38108
rect 34300 38052 34356 38108
rect 34356 38052 34360 38108
rect 34296 38048 34360 38052
rect 34376 38108 34440 38112
rect 34376 38052 34380 38108
rect 34380 38052 34436 38108
rect 34436 38052 34440 38108
rect 34376 38048 34440 38052
rect 34456 38108 34520 38112
rect 34456 38052 34460 38108
rect 34460 38052 34516 38108
rect 34516 38052 34520 38108
rect 34456 38048 34520 38052
rect 44216 38108 44280 38112
rect 44216 38052 44220 38108
rect 44220 38052 44276 38108
rect 44276 38052 44280 38108
rect 44216 38048 44280 38052
rect 44296 38108 44360 38112
rect 44296 38052 44300 38108
rect 44300 38052 44356 38108
rect 44356 38052 44360 38108
rect 44296 38048 44360 38052
rect 44376 38108 44440 38112
rect 44376 38052 44380 38108
rect 44380 38052 44436 38108
rect 44436 38052 44440 38108
rect 44376 38048 44440 38052
rect 44456 38108 44520 38112
rect 44456 38052 44460 38108
rect 44460 38052 44516 38108
rect 44516 38052 44520 38108
rect 44456 38048 44520 38052
rect 54216 38108 54280 38112
rect 54216 38052 54220 38108
rect 54220 38052 54276 38108
rect 54276 38052 54280 38108
rect 54216 38048 54280 38052
rect 54296 38108 54360 38112
rect 54296 38052 54300 38108
rect 54300 38052 54356 38108
rect 54356 38052 54360 38108
rect 54296 38048 54360 38052
rect 54376 38108 54440 38112
rect 54376 38052 54380 38108
rect 54380 38052 54436 38108
rect 54436 38052 54440 38108
rect 54376 38048 54440 38052
rect 54456 38108 54520 38112
rect 54456 38052 54460 38108
rect 54460 38052 54516 38108
rect 54516 38052 54520 38108
rect 54456 38048 54520 38052
rect 64216 38108 64280 38112
rect 64216 38052 64220 38108
rect 64220 38052 64276 38108
rect 64276 38052 64280 38108
rect 64216 38048 64280 38052
rect 64296 38108 64360 38112
rect 64296 38052 64300 38108
rect 64300 38052 64356 38108
rect 64356 38052 64360 38108
rect 64296 38048 64360 38052
rect 64376 38108 64440 38112
rect 64376 38052 64380 38108
rect 64380 38052 64436 38108
rect 64436 38052 64440 38108
rect 64376 38048 64440 38052
rect 64456 38108 64520 38112
rect 64456 38052 64460 38108
rect 64460 38052 64516 38108
rect 64516 38052 64520 38108
rect 64456 38048 64520 38052
rect 9216 37564 9280 37568
rect 9216 37508 9220 37564
rect 9220 37508 9276 37564
rect 9276 37508 9280 37564
rect 9216 37504 9280 37508
rect 9296 37564 9360 37568
rect 9296 37508 9300 37564
rect 9300 37508 9356 37564
rect 9356 37508 9360 37564
rect 9296 37504 9360 37508
rect 9376 37564 9440 37568
rect 9376 37508 9380 37564
rect 9380 37508 9436 37564
rect 9436 37508 9440 37564
rect 9376 37504 9440 37508
rect 9456 37564 9520 37568
rect 9456 37508 9460 37564
rect 9460 37508 9516 37564
rect 9516 37508 9520 37564
rect 9456 37504 9520 37508
rect 19216 37564 19280 37568
rect 19216 37508 19220 37564
rect 19220 37508 19276 37564
rect 19276 37508 19280 37564
rect 19216 37504 19280 37508
rect 19296 37564 19360 37568
rect 19296 37508 19300 37564
rect 19300 37508 19356 37564
rect 19356 37508 19360 37564
rect 19296 37504 19360 37508
rect 19376 37564 19440 37568
rect 19376 37508 19380 37564
rect 19380 37508 19436 37564
rect 19436 37508 19440 37564
rect 19376 37504 19440 37508
rect 19456 37564 19520 37568
rect 19456 37508 19460 37564
rect 19460 37508 19516 37564
rect 19516 37508 19520 37564
rect 19456 37504 19520 37508
rect 29216 37564 29280 37568
rect 29216 37508 29220 37564
rect 29220 37508 29276 37564
rect 29276 37508 29280 37564
rect 29216 37504 29280 37508
rect 29296 37564 29360 37568
rect 29296 37508 29300 37564
rect 29300 37508 29356 37564
rect 29356 37508 29360 37564
rect 29296 37504 29360 37508
rect 29376 37564 29440 37568
rect 29376 37508 29380 37564
rect 29380 37508 29436 37564
rect 29436 37508 29440 37564
rect 29376 37504 29440 37508
rect 29456 37564 29520 37568
rect 29456 37508 29460 37564
rect 29460 37508 29516 37564
rect 29516 37508 29520 37564
rect 29456 37504 29520 37508
rect 39216 37564 39280 37568
rect 39216 37508 39220 37564
rect 39220 37508 39276 37564
rect 39276 37508 39280 37564
rect 39216 37504 39280 37508
rect 39296 37564 39360 37568
rect 39296 37508 39300 37564
rect 39300 37508 39356 37564
rect 39356 37508 39360 37564
rect 39296 37504 39360 37508
rect 39376 37564 39440 37568
rect 39376 37508 39380 37564
rect 39380 37508 39436 37564
rect 39436 37508 39440 37564
rect 39376 37504 39440 37508
rect 39456 37564 39520 37568
rect 39456 37508 39460 37564
rect 39460 37508 39516 37564
rect 39516 37508 39520 37564
rect 39456 37504 39520 37508
rect 49216 37564 49280 37568
rect 49216 37508 49220 37564
rect 49220 37508 49276 37564
rect 49276 37508 49280 37564
rect 49216 37504 49280 37508
rect 49296 37564 49360 37568
rect 49296 37508 49300 37564
rect 49300 37508 49356 37564
rect 49356 37508 49360 37564
rect 49296 37504 49360 37508
rect 49376 37564 49440 37568
rect 49376 37508 49380 37564
rect 49380 37508 49436 37564
rect 49436 37508 49440 37564
rect 49376 37504 49440 37508
rect 49456 37564 49520 37568
rect 49456 37508 49460 37564
rect 49460 37508 49516 37564
rect 49516 37508 49520 37564
rect 49456 37504 49520 37508
rect 59216 37564 59280 37568
rect 59216 37508 59220 37564
rect 59220 37508 59276 37564
rect 59276 37508 59280 37564
rect 59216 37504 59280 37508
rect 59296 37564 59360 37568
rect 59296 37508 59300 37564
rect 59300 37508 59356 37564
rect 59356 37508 59360 37564
rect 59296 37504 59360 37508
rect 59376 37564 59440 37568
rect 59376 37508 59380 37564
rect 59380 37508 59436 37564
rect 59436 37508 59440 37564
rect 59376 37504 59440 37508
rect 59456 37564 59520 37568
rect 59456 37508 59460 37564
rect 59460 37508 59516 37564
rect 59516 37508 59520 37564
rect 59456 37504 59520 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 14216 37020 14280 37024
rect 14216 36964 14220 37020
rect 14220 36964 14276 37020
rect 14276 36964 14280 37020
rect 14216 36960 14280 36964
rect 14296 37020 14360 37024
rect 14296 36964 14300 37020
rect 14300 36964 14356 37020
rect 14356 36964 14360 37020
rect 14296 36960 14360 36964
rect 14376 37020 14440 37024
rect 14376 36964 14380 37020
rect 14380 36964 14436 37020
rect 14436 36964 14440 37020
rect 14376 36960 14440 36964
rect 14456 37020 14520 37024
rect 14456 36964 14460 37020
rect 14460 36964 14516 37020
rect 14516 36964 14520 37020
rect 14456 36960 14520 36964
rect 24216 37020 24280 37024
rect 24216 36964 24220 37020
rect 24220 36964 24276 37020
rect 24276 36964 24280 37020
rect 24216 36960 24280 36964
rect 24296 37020 24360 37024
rect 24296 36964 24300 37020
rect 24300 36964 24356 37020
rect 24356 36964 24360 37020
rect 24296 36960 24360 36964
rect 24376 37020 24440 37024
rect 24376 36964 24380 37020
rect 24380 36964 24436 37020
rect 24436 36964 24440 37020
rect 24376 36960 24440 36964
rect 24456 37020 24520 37024
rect 24456 36964 24460 37020
rect 24460 36964 24516 37020
rect 24516 36964 24520 37020
rect 24456 36960 24520 36964
rect 34216 37020 34280 37024
rect 34216 36964 34220 37020
rect 34220 36964 34276 37020
rect 34276 36964 34280 37020
rect 34216 36960 34280 36964
rect 34296 37020 34360 37024
rect 34296 36964 34300 37020
rect 34300 36964 34356 37020
rect 34356 36964 34360 37020
rect 34296 36960 34360 36964
rect 34376 37020 34440 37024
rect 34376 36964 34380 37020
rect 34380 36964 34436 37020
rect 34436 36964 34440 37020
rect 34376 36960 34440 36964
rect 34456 37020 34520 37024
rect 34456 36964 34460 37020
rect 34460 36964 34516 37020
rect 34516 36964 34520 37020
rect 34456 36960 34520 36964
rect 44216 37020 44280 37024
rect 44216 36964 44220 37020
rect 44220 36964 44276 37020
rect 44276 36964 44280 37020
rect 44216 36960 44280 36964
rect 44296 37020 44360 37024
rect 44296 36964 44300 37020
rect 44300 36964 44356 37020
rect 44356 36964 44360 37020
rect 44296 36960 44360 36964
rect 44376 37020 44440 37024
rect 44376 36964 44380 37020
rect 44380 36964 44436 37020
rect 44436 36964 44440 37020
rect 44376 36960 44440 36964
rect 44456 37020 44520 37024
rect 44456 36964 44460 37020
rect 44460 36964 44516 37020
rect 44516 36964 44520 37020
rect 44456 36960 44520 36964
rect 54216 37020 54280 37024
rect 54216 36964 54220 37020
rect 54220 36964 54276 37020
rect 54276 36964 54280 37020
rect 54216 36960 54280 36964
rect 54296 37020 54360 37024
rect 54296 36964 54300 37020
rect 54300 36964 54356 37020
rect 54356 36964 54360 37020
rect 54296 36960 54360 36964
rect 54376 37020 54440 37024
rect 54376 36964 54380 37020
rect 54380 36964 54436 37020
rect 54436 36964 54440 37020
rect 54376 36960 54440 36964
rect 54456 37020 54520 37024
rect 54456 36964 54460 37020
rect 54460 36964 54516 37020
rect 54516 36964 54520 37020
rect 54456 36960 54520 36964
rect 64216 37020 64280 37024
rect 64216 36964 64220 37020
rect 64220 36964 64276 37020
rect 64276 36964 64280 37020
rect 64216 36960 64280 36964
rect 64296 37020 64360 37024
rect 64296 36964 64300 37020
rect 64300 36964 64356 37020
rect 64356 36964 64360 37020
rect 64296 36960 64360 36964
rect 64376 37020 64440 37024
rect 64376 36964 64380 37020
rect 64380 36964 64436 37020
rect 64436 36964 64440 37020
rect 64376 36960 64440 36964
rect 64456 37020 64520 37024
rect 64456 36964 64460 37020
rect 64460 36964 64516 37020
rect 64516 36964 64520 37020
rect 64456 36960 64520 36964
rect 9216 36476 9280 36480
rect 9216 36420 9220 36476
rect 9220 36420 9276 36476
rect 9276 36420 9280 36476
rect 9216 36416 9280 36420
rect 9296 36476 9360 36480
rect 9296 36420 9300 36476
rect 9300 36420 9356 36476
rect 9356 36420 9360 36476
rect 9296 36416 9360 36420
rect 9376 36476 9440 36480
rect 9376 36420 9380 36476
rect 9380 36420 9436 36476
rect 9436 36420 9440 36476
rect 9376 36416 9440 36420
rect 9456 36476 9520 36480
rect 9456 36420 9460 36476
rect 9460 36420 9516 36476
rect 9516 36420 9520 36476
rect 9456 36416 9520 36420
rect 19216 36476 19280 36480
rect 19216 36420 19220 36476
rect 19220 36420 19276 36476
rect 19276 36420 19280 36476
rect 19216 36416 19280 36420
rect 19296 36476 19360 36480
rect 19296 36420 19300 36476
rect 19300 36420 19356 36476
rect 19356 36420 19360 36476
rect 19296 36416 19360 36420
rect 19376 36476 19440 36480
rect 19376 36420 19380 36476
rect 19380 36420 19436 36476
rect 19436 36420 19440 36476
rect 19376 36416 19440 36420
rect 19456 36476 19520 36480
rect 19456 36420 19460 36476
rect 19460 36420 19516 36476
rect 19516 36420 19520 36476
rect 19456 36416 19520 36420
rect 29216 36476 29280 36480
rect 29216 36420 29220 36476
rect 29220 36420 29276 36476
rect 29276 36420 29280 36476
rect 29216 36416 29280 36420
rect 29296 36476 29360 36480
rect 29296 36420 29300 36476
rect 29300 36420 29356 36476
rect 29356 36420 29360 36476
rect 29296 36416 29360 36420
rect 29376 36476 29440 36480
rect 29376 36420 29380 36476
rect 29380 36420 29436 36476
rect 29436 36420 29440 36476
rect 29376 36416 29440 36420
rect 29456 36476 29520 36480
rect 29456 36420 29460 36476
rect 29460 36420 29516 36476
rect 29516 36420 29520 36476
rect 29456 36416 29520 36420
rect 39216 36476 39280 36480
rect 39216 36420 39220 36476
rect 39220 36420 39276 36476
rect 39276 36420 39280 36476
rect 39216 36416 39280 36420
rect 39296 36476 39360 36480
rect 39296 36420 39300 36476
rect 39300 36420 39356 36476
rect 39356 36420 39360 36476
rect 39296 36416 39360 36420
rect 39376 36476 39440 36480
rect 39376 36420 39380 36476
rect 39380 36420 39436 36476
rect 39436 36420 39440 36476
rect 39376 36416 39440 36420
rect 39456 36476 39520 36480
rect 39456 36420 39460 36476
rect 39460 36420 39516 36476
rect 39516 36420 39520 36476
rect 39456 36416 39520 36420
rect 49216 36476 49280 36480
rect 49216 36420 49220 36476
rect 49220 36420 49276 36476
rect 49276 36420 49280 36476
rect 49216 36416 49280 36420
rect 49296 36476 49360 36480
rect 49296 36420 49300 36476
rect 49300 36420 49356 36476
rect 49356 36420 49360 36476
rect 49296 36416 49360 36420
rect 49376 36476 49440 36480
rect 49376 36420 49380 36476
rect 49380 36420 49436 36476
rect 49436 36420 49440 36476
rect 49376 36416 49440 36420
rect 49456 36476 49520 36480
rect 49456 36420 49460 36476
rect 49460 36420 49516 36476
rect 49516 36420 49520 36476
rect 49456 36416 49520 36420
rect 59216 36476 59280 36480
rect 59216 36420 59220 36476
rect 59220 36420 59276 36476
rect 59276 36420 59280 36476
rect 59216 36416 59280 36420
rect 59296 36476 59360 36480
rect 59296 36420 59300 36476
rect 59300 36420 59356 36476
rect 59356 36420 59360 36476
rect 59296 36416 59360 36420
rect 59376 36476 59440 36480
rect 59376 36420 59380 36476
rect 59380 36420 59436 36476
rect 59436 36420 59440 36476
rect 59376 36416 59440 36420
rect 59456 36476 59520 36480
rect 59456 36420 59460 36476
rect 59460 36420 59516 36476
rect 59516 36420 59520 36476
rect 59456 36416 59520 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 14216 35932 14280 35936
rect 14216 35876 14220 35932
rect 14220 35876 14276 35932
rect 14276 35876 14280 35932
rect 14216 35872 14280 35876
rect 14296 35932 14360 35936
rect 14296 35876 14300 35932
rect 14300 35876 14356 35932
rect 14356 35876 14360 35932
rect 14296 35872 14360 35876
rect 14376 35932 14440 35936
rect 14376 35876 14380 35932
rect 14380 35876 14436 35932
rect 14436 35876 14440 35932
rect 14376 35872 14440 35876
rect 14456 35932 14520 35936
rect 14456 35876 14460 35932
rect 14460 35876 14516 35932
rect 14516 35876 14520 35932
rect 14456 35872 14520 35876
rect 24216 35932 24280 35936
rect 24216 35876 24220 35932
rect 24220 35876 24276 35932
rect 24276 35876 24280 35932
rect 24216 35872 24280 35876
rect 24296 35932 24360 35936
rect 24296 35876 24300 35932
rect 24300 35876 24356 35932
rect 24356 35876 24360 35932
rect 24296 35872 24360 35876
rect 24376 35932 24440 35936
rect 24376 35876 24380 35932
rect 24380 35876 24436 35932
rect 24436 35876 24440 35932
rect 24376 35872 24440 35876
rect 24456 35932 24520 35936
rect 24456 35876 24460 35932
rect 24460 35876 24516 35932
rect 24516 35876 24520 35932
rect 24456 35872 24520 35876
rect 34216 35932 34280 35936
rect 34216 35876 34220 35932
rect 34220 35876 34276 35932
rect 34276 35876 34280 35932
rect 34216 35872 34280 35876
rect 34296 35932 34360 35936
rect 34296 35876 34300 35932
rect 34300 35876 34356 35932
rect 34356 35876 34360 35932
rect 34296 35872 34360 35876
rect 34376 35932 34440 35936
rect 34376 35876 34380 35932
rect 34380 35876 34436 35932
rect 34436 35876 34440 35932
rect 34376 35872 34440 35876
rect 34456 35932 34520 35936
rect 34456 35876 34460 35932
rect 34460 35876 34516 35932
rect 34516 35876 34520 35932
rect 34456 35872 34520 35876
rect 44216 35932 44280 35936
rect 44216 35876 44220 35932
rect 44220 35876 44276 35932
rect 44276 35876 44280 35932
rect 44216 35872 44280 35876
rect 44296 35932 44360 35936
rect 44296 35876 44300 35932
rect 44300 35876 44356 35932
rect 44356 35876 44360 35932
rect 44296 35872 44360 35876
rect 44376 35932 44440 35936
rect 44376 35876 44380 35932
rect 44380 35876 44436 35932
rect 44436 35876 44440 35932
rect 44376 35872 44440 35876
rect 44456 35932 44520 35936
rect 44456 35876 44460 35932
rect 44460 35876 44516 35932
rect 44516 35876 44520 35932
rect 44456 35872 44520 35876
rect 54216 35932 54280 35936
rect 54216 35876 54220 35932
rect 54220 35876 54276 35932
rect 54276 35876 54280 35932
rect 54216 35872 54280 35876
rect 54296 35932 54360 35936
rect 54296 35876 54300 35932
rect 54300 35876 54356 35932
rect 54356 35876 54360 35932
rect 54296 35872 54360 35876
rect 54376 35932 54440 35936
rect 54376 35876 54380 35932
rect 54380 35876 54436 35932
rect 54436 35876 54440 35932
rect 54376 35872 54440 35876
rect 54456 35932 54520 35936
rect 54456 35876 54460 35932
rect 54460 35876 54516 35932
rect 54516 35876 54520 35932
rect 54456 35872 54520 35876
rect 64216 35932 64280 35936
rect 64216 35876 64220 35932
rect 64220 35876 64276 35932
rect 64276 35876 64280 35932
rect 64216 35872 64280 35876
rect 64296 35932 64360 35936
rect 64296 35876 64300 35932
rect 64300 35876 64356 35932
rect 64356 35876 64360 35932
rect 64296 35872 64360 35876
rect 64376 35932 64440 35936
rect 64376 35876 64380 35932
rect 64380 35876 64436 35932
rect 64436 35876 64440 35932
rect 64376 35872 64440 35876
rect 64456 35932 64520 35936
rect 64456 35876 64460 35932
rect 64460 35876 64516 35932
rect 64516 35876 64520 35932
rect 64456 35872 64520 35876
rect 9216 35388 9280 35392
rect 9216 35332 9220 35388
rect 9220 35332 9276 35388
rect 9276 35332 9280 35388
rect 9216 35328 9280 35332
rect 9296 35388 9360 35392
rect 9296 35332 9300 35388
rect 9300 35332 9356 35388
rect 9356 35332 9360 35388
rect 9296 35328 9360 35332
rect 9376 35388 9440 35392
rect 9376 35332 9380 35388
rect 9380 35332 9436 35388
rect 9436 35332 9440 35388
rect 9376 35328 9440 35332
rect 9456 35388 9520 35392
rect 9456 35332 9460 35388
rect 9460 35332 9516 35388
rect 9516 35332 9520 35388
rect 9456 35328 9520 35332
rect 19216 35388 19280 35392
rect 19216 35332 19220 35388
rect 19220 35332 19276 35388
rect 19276 35332 19280 35388
rect 19216 35328 19280 35332
rect 19296 35388 19360 35392
rect 19296 35332 19300 35388
rect 19300 35332 19356 35388
rect 19356 35332 19360 35388
rect 19296 35328 19360 35332
rect 19376 35388 19440 35392
rect 19376 35332 19380 35388
rect 19380 35332 19436 35388
rect 19436 35332 19440 35388
rect 19376 35328 19440 35332
rect 19456 35388 19520 35392
rect 19456 35332 19460 35388
rect 19460 35332 19516 35388
rect 19516 35332 19520 35388
rect 19456 35328 19520 35332
rect 29216 35388 29280 35392
rect 29216 35332 29220 35388
rect 29220 35332 29276 35388
rect 29276 35332 29280 35388
rect 29216 35328 29280 35332
rect 29296 35388 29360 35392
rect 29296 35332 29300 35388
rect 29300 35332 29356 35388
rect 29356 35332 29360 35388
rect 29296 35328 29360 35332
rect 29376 35388 29440 35392
rect 29376 35332 29380 35388
rect 29380 35332 29436 35388
rect 29436 35332 29440 35388
rect 29376 35328 29440 35332
rect 29456 35388 29520 35392
rect 29456 35332 29460 35388
rect 29460 35332 29516 35388
rect 29516 35332 29520 35388
rect 29456 35328 29520 35332
rect 39216 35388 39280 35392
rect 39216 35332 39220 35388
rect 39220 35332 39276 35388
rect 39276 35332 39280 35388
rect 39216 35328 39280 35332
rect 39296 35388 39360 35392
rect 39296 35332 39300 35388
rect 39300 35332 39356 35388
rect 39356 35332 39360 35388
rect 39296 35328 39360 35332
rect 39376 35388 39440 35392
rect 39376 35332 39380 35388
rect 39380 35332 39436 35388
rect 39436 35332 39440 35388
rect 39376 35328 39440 35332
rect 39456 35388 39520 35392
rect 39456 35332 39460 35388
rect 39460 35332 39516 35388
rect 39516 35332 39520 35388
rect 39456 35328 39520 35332
rect 49216 35388 49280 35392
rect 49216 35332 49220 35388
rect 49220 35332 49276 35388
rect 49276 35332 49280 35388
rect 49216 35328 49280 35332
rect 49296 35388 49360 35392
rect 49296 35332 49300 35388
rect 49300 35332 49356 35388
rect 49356 35332 49360 35388
rect 49296 35328 49360 35332
rect 49376 35388 49440 35392
rect 49376 35332 49380 35388
rect 49380 35332 49436 35388
rect 49436 35332 49440 35388
rect 49376 35328 49440 35332
rect 49456 35388 49520 35392
rect 49456 35332 49460 35388
rect 49460 35332 49516 35388
rect 49516 35332 49520 35388
rect 49456 35328 49520 35332
rect 59216 35388 59280 35392
rect 59216 35332 59220 35388
rect 59220 35332 59276 35388
rect 59276 35332 59280 35388
rect 59216 35328 59280 35332
rect 59296 35388 59360 35392
rect 59296 35332 59300 35388
rect 59300 35332 59356 35388
rect 59356 35332 59360 35388
rect 59296 35328 59360 35332
rect 59376 35388 59440 35392
rect 59376 35332 59380 35388
rect 59380 35332 59436 35388
rect 59436 35332 59440 35388
rect 59376 35328 59440 35332
rect 59456 35388 59520 35392
rect 59456 35332 59460 35388
rect 59460 35332 59516 35388
rect 59516 35332 59520 35388
rect 59456 35328 59520 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 14216 34844 14280 34848
rect 14216 34788 14220 34844
rect 14220 34788 14276 34844
rect 14276 34788 14280 34844
rect 14216 34784 14280 34788
rect 14296 34844 14360 34848
rect 14296 34788 14300 34844
rect 14300 34788 14356 34844
rect 14356 34788 14360 34844
rect 14296 34784 14360 34788
rect 14376 34844 14440 34848
rect 14376 34788 14380 34844
rect 14380 34788 14436 34844
rect 14436 34788 14440 34844
rect 14376 34784 14440 34788
rect 14456 34844 14520 34848
rect 14456 34788 14460 34844
rect 14460 34788 14516 34844
rect 14516 34788 14520 34844
rect 14456 34784 14520 34788
rect 24216 34844 24280 34848
rect 24216 34788 24220 34844
rect 24220 34788 24276 34844
rect 24276 34788 24280 34844
rect 24216 34784 24280 34788
rect 24296 34844 24360 34848
rect 24296 34788 24300 34844
rect 24300 34788 24356 34844
rect 24356 34788 24360 34844
rect 24296 34784 24360 34788
rect 24376 34844 24440 34848
rect 24376 34788 24380 34844
rect 24380 34788 24436 34844
rect 24436 34788 24440 34844
rect 24376 34784 24440 34788
rect 24456 34844 24520 34848
rect 24456 34788 24460 34844
rect 24460 34788 24516 34844
rect 24516 34788 24520 34844
rect 24456 34784 24520 34788
rect 34216 34844 34280 34848
rect 34216 34788 34220 34844
rect 34220 34788 34276 34844
rect 34276 34788 34280 34844
rect 34216 34784 34280 34788
rect 34296 34844 34360 34848
rect 34296 34788 34300 34844
rect 34300 34788 34356 34844
rect 34356 34788 34360 34844
rect 34296 34784 34360 34788
rect 34376 34844 34440 34848
rect 34376 34788 34380 34844
rect 34380 34788 34436 34844
rect 34436 34788 34440 34844
rect 34376 34784 34440 34788
rect 34456 34844 34520 34848
rect 34456 34788 34460 34844
rect 34460 34788 34516 34844
rect 34516 34788 34520 34844
rect 34456 34784 34520 34788
rect 44216 34844 44280 34848
rect 44216 34788 44220 34844
rect 44220 34788 44276 34844
rect 44276 34788 44280 34844
rect 44216 34784 44280 34788
rect 44296 34844 44360 34848
rect 44296 34788 44300 34844
rect 44300 34788 44356 34844
rect 44356 34788 44360 34844
rect 44296 34784 44360 34788
rect 44376 34844 44440 34848
rect 44376 34788 44380 34844
rect 44380 34788 44436 34844
rect 44436 34788 44440 34844
rect 44376 34784 44440 34788
rect 44456 34844 44520 34848
rect 44456 34788 44460 34844
rect 44460 34788 44516 34844
rect 44516 34788 44520 34844
rect 44456 34784 44520 34788
rect 54216 34844 54280 34848
rect 54216 34788 54220 34844
rect 54220 34788 54276 34844
rect 54276 34788 54280 34844
rect 54216 34784 54280 34788
rect 54296 34844 54360 34848
rect 54296 34788 54300 34844
rect 54300 34788 54356 34844
rect 54356 34788 54360 34844
rect 54296 34784 54360 34788
rect 54376 34844 54440 34848
rect 54376 34788 54380 34844
rect 54380 34788 54436 34844
rect 54436 34788 54440 34844
rect 54376 34784 54440 34788
rect 54456 34844 54520 34848
rect 54456 34788 54460 34844
rect 54460 34788 54516 34844
rect 54516 34788 54520 34844
rect 54456 34784 54520 34788
rect 64216 34844 64280 34848
rect 64216 34788 64220 34844
rect 64220 34788 64276 34844
rect 64276 34788 64280 34844
rect 64216 34784 64280 34788
rect 64296 34844 64360 34848
rect 64296 34788 64300 34844
rect 64300 34788 64356 34844
rect 64356 34788 64360 34844
rect 64296 34784 64360 34788
rect 64376 34844 64440 34848
rect 64376 34788 64380 34844
rect 64380 34788 64436 34844
rect 64436 34788 64440 34844
rect 64376 34784 64440 34788
rect 64456 34844 64520 34848
rect 64456 34788 64460 34844
rect 64460 34788 64516 34844
rect 64516 34788 64520 34844
rect 64456 34784 64520 34788
rect 9216 34300 9280 34304
rect 9216 34244 9220 34300
rect 9220 34244 9276 34300
rect 9276 34244 9280 34300
rect 9216 34240 9280 34244
rect 9296 34300 9360 34304
rect 9296 34244 9300 34300
rect 9300 34244 9356 34300
rect 9356 34244 9360 34300
rect 9296 34240 9360 34244
rect 9376 34300 9440 34304
rect 9376 34244 9380 34300
rect 9380 34244 9436 34300
rect 9436 34244 9440 34300
rect 9376 34240 9440 34244
rect 9456 34300 9520 34304
rect 9456 34244 9460 34300
rect 9460 34244 9516 34300
rect 9516 34244 9520 34300
rect 9456 34240 9520 34244
rect 19216 34300 19280 34304
rect 19216 34244 19220 34300
rect 19220 34244 19276 34300
rect 19276 34244 19280 34300
rect 19216 34240 19280 34244
rect 19296 34300 19360 34304
rect 19296 34244 19300 34300
rect 19300 34244 19356 34300
rect 19356 34244 19360 34300
rect 19296 34240 19360 34244
rect 19376 34300 19440 34304
rect 19376 34244 19380 34300
rect 19380 34244 19436 34300
rect 19436 34244 19440 34300
rect 19376 34240 19440 34244
rect 19456 34300 19520 34304
rect 19456 34244 19460 34300
rect 19460 34244 19516 34300
rect 19516 34244 19520 34300
rect 19456 34240 19520 34244
rect 29216 34300 29280 34304
rect 29216 34244 29220 34300
rect 29220 34244 29276 34300
rect 29276 34244 29280 34300
rect 29216 34240 29280 34244
rect 29296 34300 29360 34304
rect 29296 34244 29300 34300
rect 29300 34244 29356 34300
rect 29356 34244 29360 34300
rect 29296 34240 29360 34244
rect 29376 34300 29440 34304
rect 29376 34244 29380 34300
rect 29380 34244 29436 34300
rect 29436 34244 29440 34300
rect 29376 34240 29440 34244
rect 29456 34300 29520 34304
rect 29456 34244 29460 34300
rect 29460 34244 29516 34300
rect 29516 34244 29520 34300
rect 29456 34240 29520 34244
rect 39216 34300 39280 34304
rect 39216 34244 39220 34300
rect 39220 34244 39276 34300
rect 39276 34244 39280 34300
rect 39216 34240 39280 34244
rect 39296 34300 39360 34304
rect 39296 34244 39300 34300
rect 39300 34244 39356 34300
rect 39356 34244 39360 34300
rect 39296 34240 39360 34244
rect 39376 34300 39440 34304
rect 39376 34244 39380 34300
rect 39380 34244 39436 34300
rect 39436 34244 39440 34300
rect 39376 34240 39440 34244
rect 39456 34300 39520 34304
rect 39456 34244 39460 34300
rect 39460 34244 39516 34300
rect 39516 34244 39520 34300
rect 39456 34240 39520 34244
rect 49216 34300 49280 34304
rect 49216 34244 49220 34300
rect 49220 34244 49276 34300
rect 49276 34244 49280 34300
rect 49216 34240 49280 34244
rect 49296 34300 49360 34304
rect 49296 34244 49300 34300
rect 49300 34244 49356 34300
rect 49356 34244 49360 34300
rect 49296 34240 49360 34244
rect 49376 34300 49440 34304
rect 49376 34244 49380 34300
rect 49380 34244 49436 34300
rect 49436 34244 49440 34300
rect 49376 34240 49440 34244
rect 49456 34300 49520 34304
rect 49456 34244 49460 34300
rect 49460 34244 49516 34300
rect 49516 34244 49520 34300
rect 49456 34240 49520 34244
rect 59216 34300 59280 34304
rect 59216 34244 59220 34300
rect 59220 34244 59276 34300
rect 59276 34244 59280 34300
rect 59216 34240 59280 34244
rect 59296 34300 59360 34304
rect 59296 34244 59300 34300
rect 59300 34244 59356 34300
rect 59356 34244 59360 34300
rect 59296 34240 59360 34244
rect 59376 34300 59440 34304
rect 59376 34244 59380 34300
rect 59380 34244 59436 34300
rect 59436 34244 59440 34300
rect 59376 34240 59440 34244
rect 59456 34300 59520 34304
rect 59456 34244 59460 34300
rect 59460 34244 59516 34300
rect 59516 34244 59520 34300
rect 59456 34240 59520 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 14216 33756 14280 33760
rect 14216 33700 14220 33756
rect 14220 33700 14276 33756
rect 14276 33700 14280 33756
rect 14216 33696 14280 33700
rect 14296 33756 14360 33760
rect 14296 33700 14300 33756
rect 14300 33700 14356 33756
rect 14356 33700 14360 33756
rect 14296 33696 14360 33700
rect 14376 33756 14440 33760
rect 14376 33700 14380 33756
rect 14380 33700 14436 33756
rect 14436 33700 14440 33756
rect 14376 33696 14440 33700
rect 14456 33756 14520 33760
rect 14456 33700 14460 33756
rect 14460 33700 14516 33756
rect 14516 33700 14520 33756
rect 14456 33696 14520 33700
rect 24216 33756 24280 33760
rect 24216 33700 24220 33756
rect 24220 33700 24276 33756
rect 24276 33700 24280 33756
rect 24216 33696 24280 33700
rect 24296 33756 24360 33760
rect 24296 33700 24300 33756
rect 24300 33700 24356 33756
rect 24356 33700 24360 33756
rect 24296 33696 24360 33700
rect 24376 33756 24440 33760
rect 24376 33700 24380 33756
rect 24380 33700 24436 33756
rect 24436 33700 24440 33756
rect 24376 33696 24440 33700
rect 24456 33756 24520 33760
rect 24456 33700 24460 33756
rect 24460 33700 24516 33756
rect 24516 33700 24520 33756
rect 24456 33696 24520 33700
rect 34216 33756 34280 33760
rect 34216 33700 34220 33756
rect 34220 33700 34276 33756
rect 34276 33700 34280 33756
rect 34216 33696 34280 33700
rect 34296 33756 34360 33760
rect 34296 33700 34300 33756
rect 34300 33700 34356 33756
rect 34356 33700 34360 33756
rect 34296 33696 34360 33700
rect 34376 33756 34440 33760
rect 34376 33700 34380 33756
rect 34380 33700 34436 33756
rect 34436 33700 34440 33756
rect 34376 33696 34440 33700
rect 34456 33756 34520 33760
rect 34456 33700 34460 33756
rect 34460 33700 34516 33756
rect 34516 33700 34520 33756
rect 34456 33696 34520 33700
rect 44216 33756 44280 33760
rect 44216 33700 44220 33756
rect 44220 33700 44276 33756
rect 44276 33700 44280 33756
rect 44216 33696 44280 33700
rect 44296 33756 44360 33760
rect 44296 33700 44300 33756
rect 44300 33700 44356 33756
rect 44356 33700 44360 33756
rect 44296 33696 44360 33700
rect 44376 33756 44440 33760
rect 44376 33700 44380 33756
rect 44380 33700 44436 33756
rect 44436 33700 44440 33756
rect 44376 33696 44440 33700
rect 44456 33756 44520 33760
rect 44456 33700 44460 33756
rect 44460 33700 44516 33756
rect 44516 33700 44520 33756
rect 44456 33696 44520 33700
rect 54216 33756 54280 33760
rect 54216 33700 54220 33756
rect 54220 33700 54276 33756
rect 54276 33700 54280 33756
rect 54216 33696 54280 33700
rect 54296 33756 54360 33760
rect 54296 33700 54300 33756
rect 54300 33700 54356 33756
rect 54356 33700 54360 33756
rect 54296 33696 54360 33700
rect 54376 33756 54440 33760
rect 54376 33700 54380 33756
rect 54380 33700 54436 33756
rect 54436 33700 54440 33756
rect 54376 33696 54440 33700
rect 54456 33756 54520 33760
rect 54456 33700 54460 33756
rect 54460 33700 54516 33756
rect 54516 33700 54520 33756
rect 54456 33696 54520 33700
rect 64216 33756 64280 33760
rect 64216 33700 64220 33756
rect 64220 33700 64276 33756
rect 64276 33700 64280 33756
rect 64216 33696 64280 33700
rect 64296 33756 64360 33760
rect 64296 33700 64300 33756
rect 64300 33700 64356 33756
rect 64356 33700 64360 33756
rect 64296 33696 64360 33700
rect 64376 33756 64440 33760
rect 64376 33700 64380 33756
rect 64380 33700 64436 33756
rect 64436 33700 64440 33756
rect 64376 33696 64440 33700
rect 64456 33756 64520 33760
rect 64456 33700 64460 33756
rect 64460 33700 64516 33756
rect 64516 33700 64520 33756
rect 64456 33696 64520 33700
rect 9216 33212 9280 33216
rect 9216 33156 9220 33212
rect 9220 33156 9276 33212
rect 9276 33156 9280 33212
rect 9216 33152 9280 33156
rect 9296 33212 9360 33216
rect 9296 33156 9300 33212
rect 9300 33156 9356 33212
rect 9356 33156 9360 33212
rect 9296 33152 9360 33156
rect 9376 33212 9440 33216
rect 9376 33156 9380 33212
rect 9380 33156 9436 33212
rect 9436 33156 9440 33212
rect 9376 33152 9440 33156
rect 9456 33212 9520 33216
rect 9456 33156 9460 33212
rect 9460 33156 9516 33212
rect 9516 33156 9520 33212
rect 9456 33152 9520 33156
rect 19216 33212 19280 33216
rect 19216 33156 19220 33212
rect 19220 33156 19276 33212
rect 19276 33156 19280 33212
rect 19216 33152 19280 33156
rect 19296 33212 19360 33216
rect 19296 33156 19300 33212
rect 19300 33156 19356 33212
rect 19356 33156 19360 33212
rect 19296 33152 19360 33156
rect 19376 33212 19440 33216
rect 19376 33156 19380 33212
rect 19380 33156 19436 33212
rect 19436 33156 19440 33212
rect 19376 33152 19440 33156
rect 19456 33212 19520 33216
rect 19456 33156 19460 33212
rect 19460 33156 19516 33212
rect 19516 33156 19520 33212
rect 19456 33152 19520 33156
rect 29216 33212 29280 33216
rect 29216 33156 29220 33212
rect 29220 33156 29276 33212
rect 29276 33156 29280 33212
rect 29216 33152 29280 33156
rect 29296 33212 29360 33216
rect 29296 33156 29300 33212
rect 29300 33156 29356 33212
rect 29356 33156 29360 33212
rect 29296 33152 29360 33156
rect 29376 33212 29440 33216
rect 29376 33156 29380 33212
rect 29380 33156 29436 33212
rect 29436 33156 29440 33212
rect 29376 33152 29440 33156
rect 29456 33212 29520 33216
rect 29456 33156 29460 33212
rect 29460 33156 29516 33212
rect 29516 33156 29520 33212
rect 29456 33152 29520 33156
rect 39216 33212 39280 33216
rect 39216 33156 39220 33212
rect 39220 33156 39276 33212
rect 39276 33156 39280 33212
rect 39216 33152 39280 33156
rect 39296 33212 39360 33216
rect 39296 33156 39300 33212
rect 39300 33156 39356 33212
rect 39356 33156 39360 33212
rect 39296 33152 39360 33156
rect 39376 33212 39440 33216
rect 39376 33156 39380 33212
rect 39380 33156 39436 33212
rect 39436 33156 39440 33212
rect 39376 33152 39440 33156
rect 39456 33212 39520 33216
rect 39456 33156 39460 33212
rect 39460 33156 39516 33212
rect 39516 33156 39520 33212
rect 39456 33152 39520 33156
rect 49216 33212 49280 33216
rect 49216 33156 49220 33212
rect 49220 33156 49276 33212
rect 49276 33156 49280 33212
rect 49216 33152 49280 33156
rect 49296 33212 49360 33216
rect 49296 33156 49300 33212
rect 49300 33156 49356 33212
rect 49356 33156 49360 33212
rect 49296 33152 49360 33156
rect 49376 33212 49440 33216
rect 49376 33156 49380 33212
rect 49380 33156 49436 33212
rect 49436 33156 49440 33212
rect 49376 33152 49440 33156
rect 49456 33212 49520 33216
rect 49456 33156 49460 33212
rect 49460 33156 49516 33212
rect 49516 33156 49520 33212
rect 49456 33152 49520 33156
rect 59216 33212 59280 33216
rect 59216 33156 59220 33212
rect 59220 33156 59276 33212
rect 59276 33156 59280 33212
rect 59216 33152 59280 33156
rect 59296 33212 59360 33216
rect 59296 33156 59300 33212
rect 59300 33156 59356 33212
rect 59356 33156 59360 33212
rect 59296 33152 59360 33156
rect 59376 33212 59440 33216
rect 59376 33156 59380 33212
rect 59380 33156 59436 33212
rect 59436 33156 59440 33212
rect 59376 33152 59440 33156
rect 59456 33212 59520 33216
rect 59456 33156 59460 33212
rect 59460 33156 59516 33212
rect 59516 33156 59520 33212
rect 59456 33152 59520 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 14216 32668 14280 32672
rect 14216 32612 14220 32668
rect 14220 32612 14276 32668
rect 14276 32612 14280 32668
rect 14216 32608 14280 32612
rect 14296 32668 14360 32672
rect 14296 32612 14300 32668
rect 14300 32612 14356 32668
rect 14356 32612 14360 32668
rect 14296 32608 14360 32612
rect 14376 32668 14440 32672
rect 14376 32612 14380 32668
rect 14380 32612 14436 32668
rect 14436 32612 14440 32668
rect 14376 32608 14440 32612
rect 14456 32668 14520 32672
rect 14456 32612 14460 32668
rect 14460 32612 14516 32668
rect 14516 32612 14520 32668
rect 14456 32608 14520 32612
rect 24216 32668 24280 32672
rect 24216 32612 24220 32668
rect 24220 32612 24276 32668
rect 24276 32612 24280 32668
rect 24216 32608 24280 32612
rect 24296 32668 24360 32672
rect 24296 32612 24300 32668
rect 24300 32612 24356 32668
rect 24356 32612 24360 32668
rect 24296 32608 24360 32612
rect 24376 32668 24440 32672
rect 24376 32612 24380 32668
rect 24380 32612 24436 32668
rect 24436 32612 24440 32668
rect 24376 32608 24440 32612
rect 24456 32668 24520 32672
rect 24456 32612 24460 32668
rect 24460 32612 24516 32668
rect 24516 32612 24520 32668
rect 24456 32608 24520 32612
rect 34216 32668 34280 32672
rect 34216 32612 34220 32668
rect 34220 32612 34276 32668
rect 34276 32612 34280 32668
rect 34216 32608 34280 32612
rect 34296 32668 34360 32672
rect 34296 32612 34300 32668
rect 34300 32612 34356 32668
rect 34356 32612 34360 32668
rect 34296 32608 34360 32612
rect 34376 32668 34440 32672
rect 34376 32612 34380 32668
rect 34380 32612 34436 32668
rect 34436 32612 34440 32668
rect 34376 32608 34440 32612
rect 34456 32668 34520 32672
rect 34456 32612 34460 32668
rect 34460 32612 34516 32668
rect 34516 32612 34520 32668
rect 34456 32608 34520 32612
rect 44216 32668 44280 32672
rect 44216 32612 44220 32668
rect 44220 32612 44276 32668
rect 44276 32612 44280 32668
rect 44216 32608 44280 32612
rect 44296 32668 44360 32672
rect 44296 32612 44300 32668
rect 44300 32612 44356 32668
rect 44356 32612 44360 32668
rect 44296 32608 44360 32612
rect 44376 32668 44440 32672
rect 44376 32612 44380 32668
rect 44380 32612 44436 32668
rect 44436 32612 44440 32668
rect 44376 32608 44440 32612
rect 44456 32668 44520 32672
rect 44456 32612 44460 32668
rect 44460 32612 44516 32668
rect 44516 32612 44520 32668
rect 44456 32608 44520 32612
rect 54216 32668 54280 32672
rect 54216 32612 54220 32668
rect 54220 32612 54276 32668
rect 54276 32612 54280 32668
rect 54216 32608 54280 32612
rect 54296 32668 54360 32672
rect 54296 32612 54300 32668
rect 54300 32612 54356 32668
rect 54356 32612 54360 32668
rect 54296 32608 54360 32612
rect 54376 32668 54440 32672
rect 54376 32612 54380 32668
rect 54380 32612 54436 32668
rect 54436 32612 54440 32668
rect 54376 32608 54440 32612
rect 54456 32668 54520 32672
rect 54456 32612 54460 32668
rect 54460 32612 54516 32668
rect 54516 32612 54520 32668
rect 54456 32608 54520 32612
rect 64216 32668 64280 32672
rect 64216 32612 64220 32668
rect 64220 32612 64276 32668
rect 64276 32612 64280 32668
rect 64216 32608 64280 32612
rect 64296 32668 64360 32672
rect 64296 32612 64300 32668
rect 64300 32612 64356 32668
rect 64356 32612 64360 32668
rect 64296 32608 64360 32612
rect 64376 32668 64440 32672
rect 64376 32612 64380 32668
rect 64380 32612 64436 32668
rect 64436 32612 64440 32668
rect 64376 32608 64440 32612
rect 64456 32668 64520 32672
rect 64456 32612 64460 32668
rect 64460 32612 64516 32668
rect 64516 32612 64520 32668
rect 64456 32608 64520 32612
rect 38700 32404 38764 32468
rect 9216 32124 9280 32128
rect 9216 32068 9220 32124
rect 9220 32068 9276 32124
rect 9276 32068 9280 32124
rect 9216 32064 9280 32068
rect 9296 32124 9360 32128
rect 9296 32068 9300 32124
rect 9300 32068 9356 32124
rect 9356 32068 9360 32124
rect 9296 32064 9360 32068
rect 9376 32124 9440 32128
rect 9376 32068 9380 32124
rect 9380 32068 9436 32124
rect 9436 32068 9440 32124
rect 9376 32064 9440 32068
rect 9456 32124 9520 32128
rect 9456 32068 9460 32124
rect 9460 32068 9516 32124
rect 9516 32068 9520 32124
rect 9456 32064 9520 32068
rect 19216 32124 19280 32128
rect 19216 32068 19220 32124
rect 19220 32068 19276 32124
rect 19276 32068 19280 32124
rect 19216 32064 19280 32068
rect 19296 32124 19360 32128
rect 19296 32068 19300 32124
rect 19300 32068 19356 32124
rect 19356 32068 19360 32124
rect 19296 32064 19360 32068
rect 19376 32124 19440 32128
rect 19376 32068 19380 32124
rect 19380 32068 19436 32124
rect 19436 32068 19440 32124
rect 19376 32064 19440 32068
rect 19456 32124 19520 32128
rect 19456 32068 19460 32124
rect 19460 32068 19516 32124
rect 19516 32068 19520 32124
rect 19456 32064 19520 32068
rect 29216 32124 29280 32128
rect 29216 32068 29220 32124
rect 29220 32068 29276 32124
rect 29276 32068 29280 32124
rect 29216 32064 29280 32068
rect 29296 32124 29360 32128
rect 29296 32068 29300 32124
rect 29300 32068 29356 32124
rect 29356 32068 29360 32124
rect 29296 32064 29360 32068
rect 29376 32124 29440 32128
rect 29376 32068 29380 32124
rect 29380 32068 29436 32124
rect 29436 32068 29440 32124
rect 29376 32064 29440 32068
rect 29456 32124 29520 32128
rect 29456 32068 29460 32124
rect 29460 32068 29516 32124
rect 29516 32068 29520 32124
rect 29456 32064 29520 32068
rect 39216 32124 39280 32128
rect 39216 32068 39220 32124
rect 39220 32068 39276 32124
rect 39276 32068 39280 32124
rect 39216 32064 39280 32068
rect 39296 32124 39360 32128
rect 39296 32068 39300 32124
rect 39300 32068 39356 32124
rect 39356 32068 39360 32124
rect 39296 32064 39360 32068
rect 39376 32124 39440 32128
rect 39376 32068 39380 32124
rect 39380 32068 39436 32124
rect 39436 32068 39440 32124
rect 39376 32064 39440 32068
rect 39456 32124 39520 32128
rect 39456 32068 39460 32124
rect 39460 32068 39516 32124
rect 39516 32068 39520 32124
rect 39456 32064 39520 32068
rect 49216 32124 49280 32128
rect 49216 32068 49220 32124
rect 49220 32068 49276 32124
rect 49276 32068 49280 32124
rect 49216 32064 49280 32068
rect 49296 32124 49360 32128
rect 49296 32068 49300 32124
rect 49300 32068 49356 32124
rect 49356 32068 49360 32124
rect 49296 32064 49360 32068
rect 49376 32124 49440 32128
rect 49376 32068 49380 32124
rect 49380 32068 49436 32124
rect 49436 32068 49440 32124
rect 49376 32064 49440 32068
rect 49456 32124 49520 32128
rect 49456 32068 49460 32124
rect 49460 32068 49516 32124
rect 49516 32068 49520 32124
rect 49456 32064 49520 32068
rect 59216 32124 59280 32128
rect 59216 32068 59220 32124
rect 59220 32068 59276 32124
rect 59276 32068 59280 32124
rect 59216 32064 59280 32068
rect 59296 32124 59360 32128
rect 59296 32068 59300 32124
rect 59300 32068 59356 32124
rect 59356 32068 59360 32124
rect 59296 32064 59360 32068
rect 59376 32124 59440 32128
rect 59376 32068 59380 32124
rect 59380 32068 59436 32124
rect 59436 32068 59440 32124
rect 59376 32064 59440 32068
rect 59456 32124 59520 32128
rect 59456 32068 59460 32124
rect 59460 32068 59516 32124
rect 59516 32068 59520 32124
rect 59456 32064 59520 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 14216 31580 14280 31584
rect 14216 31524 14220 31580
rect 14220 31524 14276 31580
rect 14276 31524 14280 31580
rect 14216 31520 14280 31524
rect 14296 31580 14360 31584
rect 14296 31524 14300 31580
rect 14300 31524 14356 31580
rect 14356 31524 14360 31580
rect 14296 31520 14360 31524
rect 14376 31580 14440 31584
rect 14376 31524 14380 31580
rect 14380 31524 14436 31580
rect 14436 31524 14440 31580
rect 14376 31520 14440 31524
rect 14456 31580 14520 31584
rect 14456 31524 14460 31580
rect 14460 31524 14516 31580
rect 14516 31524 14520 31580
rect 14456 31520 14520 31524
rect 24216 31580 24280 31584
rect 24216 31524 24220 31580
rect 24220 31524 24276 31580
rect 24276 31524 24280 31580
rect 24216 31520 24280 31524
rect 24296 31580 24360 31584
rect 24296 31524 24300 31580
rect 24300 31524 24356 31580
rect 24356 31524 24360 31580
rect 24296 31520 24360 31524
rect 24376 31580 24440 31584
rect 24376 31524 24380 31580
rect 24380 31524 24436 31580
rect 24436 31524 24440 31580
rect 24376 31520 24440 31524
rect 24456 31580 24520 31584
rect 24456 31524 24460 31580
rect 24460 31524 24516 31580
rect 24516 31524 24520 31580
rect 24456 31520 24520 31524
rect 34216 31580 34280 31584
rect 34216 31524 34220 31580
rect 34220 31524 34276 31580
rect 34276 31524 34280 31580
rect 34216 31520 34280 31524
rect 34296 31580 34360 31584
rect 34296 31524 34300 31580
rect 34300 31524 34356 31580
rect 34356 31524 34360 31580
rect 34296 31520 34360 31524
rect 34376 31580 34440 31584
rect 34376 31524 34380 31580
rect 34380 31524 34436 31580
rect 34436 31524 34440 31580
rect 34376 31520 34440 31524
rect 34456 31580 34520 31584
rect 34456 31524 34460 31580
rect 34460 31524 34516 31580
rect 34516 31524 34520 31580
rect 34456 31520 34520 31524
rect 44216 31580 44280 31584
rect 44216 31524 44220 31580
rect 44220 31524 44276 31580
rect 44276 31524 44280 31580
rect 44216 31520 44280 31524
rect 44296 31580 44360 31584
rect 44296 31524 44300 31580
rect 44300 31524 44356 31580
rect 44356 31524 44360 31580
rect 44296 31520 44360 31524
rect 44376 31580 44440 31584
rect 44376 31524 44380 31580
rect 44380 31524 44436 31580
rect 44436 31524 44440 31580
rect 44376 31520 44440 31524
rect 44456 31580 44520 31584
rect 44456 31524 44460 31580
rect 44460 31524 44516 31580
rect 44516 31524 44520 31580
rect 44456 31520 44520 31524
rect 54216 31580 54280 31584
rect 54216 31524 54220 31580
rect 54220 31524 54276 31580
rect 54276 31524 54280 31580
rect 54216 31520 54280 31524
rect 54296 31580 54360 31584
rect 54296 31524 54300 31580
rect 54300 31524 54356 31580
rect 54356 31524 54360 31580
rect 54296 31520 54360 31524
rect 54376 31580 54440 31584
rect 54376 31524 54380 31580
rect 54380 31524 54436 31580
rect 54436 31524 54440 31580
rect 54376 31520 54440 31524
rect 54456 31580 54520 31584
rect 54456 31524 54460 31580
rect 54460 31524 54516 31580
rect 54516 31524 54520 31580
rect 54456 31520 54520 31524
rect 64216 31580 64280 31584
rect 64216 31524 64220 31580
rect 64220 31524 64276 31580
rect 64276 31524 64280 31580
rect 64216 31520 64280 31524
rect 64296 31580 64360 31584
rect 64296 31524 64300 31580
rect 64300 31524 64356 31580
rect 64356 31524 64360 31580
rect 64296 31520 64360 31524
rect 64376 31580 64440 31584
rect 64376 31524 64380 31580
rect 64380 31524 64436 31580
rect 64436 31524 64440 31580
rect 64376 31520 64440 31524
rect 64456 31580 64520 31584
rect 64456 31524 64460 31580
rect 64460 31524 64516 31580
rect 64516 31524 64520 31580
rect 64456 31520 64520 31524
rect 9216 31036 9280 31040
rect 9216 30980 9220 31036
rect 9220 30980 9276 31036
rect 9276 30980 9280 31036
rect 9216 30976 9280 30980
rect 9296 31036 9360 31040
rect 9296 30980 9300 31036
rect 9300 30980 9356 31036
rect 9356 30980 9360 31036
rect 9296 30976 9360 30980
rect 9376 31036 9440 31040
rect 9376 30980 9380 31036
rect 9380 30980 9436 31036
rect 9436 30980 9440 31036
rect 9376 30976 9440 30980
rect 9456 31036 9520 31040
rect 9456 30980 9460 31036
rect 9460 30980 9516 31036
rect 9516 30980 9520 31036
rect 9456 30976 9520 30980
rect 19216 31036 19280 31040
rect 19216 30980 19220 31036
rect 19220 30980 19276 31036
rect 19276 30980 19280 31036
rect 19216 30976 19280 30980
rect 19296 31036 19360 31040
rect 19296 30980 19300 31036
rect 19300 30980 19356 31036
rect 19356 30980 19360 31036
rect 19296 30976 19360 30980
rect 19376 31036 19440 31040
rect 19376 30980 19380 31036
rect 19380 30980 19436 31036
rect 19436 30980 19440 31036
rect 19376 30976 19440 30980
rect 19456 31036 19520 31040
rect 19456 30980 19460 31036
rect 19460 30980 19516 31036
rect 19516 30980 19520 31036
rect 19456 30976 19520 30980
rect 29216 31036 29280 31040
rect 29216 30980 29220 31036
rect 29220 30980 29276 31036
rect 29276 30980 29280 31036
rect 29216 30976 29280 30980
rect 29296 31036 29360 31040
rect 29296 30980 29300 31036
rect 29300 30980 29356 31036
rect 29356 30980 29360 31036
rect 29296 30976 29360 30980
rect 29376 31036 29440 31040
rect 29376 30980 29380 31036
rect 29380 30980 29436 31036
rect 29436 30980 29440 31036
rect 29376 30976 29440 30980
rect 29456 31036 29520 31040
rect 29456 30980 29460 31036
rect 29460 30980 29516 31036
rect 29516 30980 29520 31036
rect 29456 30976 29520 30980
rect 39216 31036 39280 31040
rect 39216 30980 39220 31036
rect 39220 30980 39276 31036
rect 39276 30980 39280 31036
rect 39216 30976 39280 30980
rect 39296 31036 39360 31040
rect 39296 30980 39300 31036
rect 39300 30980 39356 31036
rect 39356 30980 39360 31036
rect 39296 30976 39360 30980
rect 39376 31036 39440 31040
rect 39376 30980 39380 31036
rect 39380 30980 39436 31036
rect 39436 30980 39440 31036
rect 39376 30976 39440 30980
rect 39456 31036 39520 31040
rect 39456 30980 39460 31036
rect 39460 30980 39516 31036
rect 39516 30980 39520 31036
rect 39456 30976 39520 30980
rect 49216 31036 49280 31040
rect 49216 30980 49220 31036
rect 49220 30980 49276 31036
rect 49276 30980 49280 31036
rect 49216 30976 49280 30980
rect 49296 31036 49360 31040
rect 49296 30980 49300 31036
rect 49300 30980 49356 31036
rect 49356 30980 49360 31036
rect 49296 30976 49360 30980
rect 49376 31036 49440 31040
rect 49376 30980 49380 31036
rect 49380 30980 49436 31036
rect 49436 30980 49440 31036
rect 49376 30976 49440 30980
rect 49456 31036 49520 31040
rect 49456 30980 49460 31036
rect 49460 30980 49516 31036
rect 49516 30980 49520 31036
rect 49456 30976 49520 30980
rect 59216 31036 59280 31040
rect 59216 30980 59220 31036
rect 59220 30980 59276 31036
rect 59276 30980 59280 31036
rect 59216 30976 59280 30980
rect 59296 31036 59360 31040
rect 59296 30980 59300 31036
rect 59300 30980 59356 31036
rect 59356 30980 59360 31036
rect 59296 30976 59360 30980
rect 59376 31036 59440 31040
rect 59376 30980 59380 31036
rect 59380 30980 59436 31036
rect 59436 30980 59440 31036
rect 59376 30976 59440 30980
rect 59456 31036 59520 31040
rect 59456 30980 59460 31036
rect 59460 30980 59516 31036
rect 59516 30980 59520 31036
rect 59456 30976 59520 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 14216 30492 14280 30496
rect 14216 30436 14220 30492
rect 14220 30436 14276 30492
rect 14276 30436 14280 30492
rect 14216 30432 14280 30436
rect 14296 30492 14360 30496
rect 14296 30436 14300 30492
rect 14300 30436 14356 30492
rect 14356 30436 14360 30492
rect 14296 30432 14360 30436
rect 14376 30492 14440 30496
rect 14376 30436 14380 30492
rect 14380 30436 14436 30492
rect 14436 30436 14440 30492
rect 14376 30432 14440 30436
rect 14456 30492 14520 30496
rect 14456 30436 14460 30492
rect 14460 30436 14516 30492
rect 14516 30436 14520 30492
rect 14456 30432 14520 30436
rect 24216 30492 24280 30496
rect 24216 30436 24220 30492
rect 24220 30436 24276 30492
rect 24276 30436 24280 30492
rect 24216 30432 24280 30436
rect 24296 30492 24360 30496
rect 24296 30436 24300 30492
rect 24300 30436 24356 30492
rect 24356 30436 24360 30492
rect 24296 30432 24360 30436
rect 24376 30492 24440 30496
rect 24376 30436 24380 30492
rect 24380 30436 24436 30492
rect 24436 30436 24440 30492
rect 24376 30432 24440 30436
rect 24456 30492 24520 30496
rect 24456 30436 24460 30492
rect 24460 30436 24516 30492
rect 24516 30436 24520 30492
rect 24456 30432 24520 30436
rect 34216 30492 34280 30496
rect 34216 30436 34220 30492
rect 34220 30436 34276 30492
rect 34276 30436 34280 30492
rect 34216 30432 34280 30436
rect 34296 30492 34360 30496
rect 34296 30436 34300 30492
rect 34300 30436 34356 30492
rect 34356 30436 34360 30492
rect 34296 30432 34360 30436
rect 34376 30492 34440 30496
rect 34376 30436 34380 30492
rect 34380 30436 34436 30492
rect 34436 30436 34440 30492
rect 34376 30432 34440 30436
rect 34456 30492 34520 30496
rect 34456 30436 34460 30492
rect 34460 30436 34516 30492
rect 34516 30436 34520 30492
rect 34456 30432 34520 30436
rect 44216 30492 44280 30496
rect 44216 30436 44220 30492
rect 44220 30436 44276 30492
rect 44276 30436 44280 30492
rect 44216 30432 44280 30436
rect 44296 30492 44360 30496
rect 44296 30436 44300 30492
rect 44300 30436 44356 30492
rect 44356 30436 44360 30492
rect 44296 30432 44360 30436
rect 44376 30492 44440 30496
rect 44376 30436 44380 30492
rect 44380 30436 44436 30492
rect 44436 30436 44440 30492
rect 44376 30432 44440 30436
rect 44456 30492 44520 30496
rect 44456 30436 44460 30492
rect 44460 30436 44516 30492
rect 44516 30436 44520 30492
rect 44456 30432 44520 30436
rect 54216 30492 54280 30496
rect 54216 30436 54220 30492
rect 54220 30436 54276 30492
rect 54276 30436 54280 30492
rect 54216 30432 54280 30436
rect 54296 30492 54360 30496
rect 54296 30436 54300 30492
rect 54300 30436 54356 30492
rect 54356 30436 54360 30492
rect 54296 30432 54360 30436
rect 54376 30492 54440 30496
rect 54376 30436 54380 30492
rect 54380 30436 54436 30492
rect 54436 30436 54440 30492
rect 54376 30432 54440 30436
rect 54456 30492 54520 30496
rect 54456 30436 54460 30492
rect 54460 30436 54516 30492
rect 54516 30436 54520 30492
rect 54456 30432 54520 30436
rect 64216 30492 64280 30496
rect 64216 30436 64220 30492
rect 64220 30436 64276 30492
rect 64276 30436 64280 30492
rect 64216 30432 64280 30436
rect 64296 30492 64360 30496
rect 64296 30436 64300 30492
rect 64300 30436 64356 30492
rect 64356 30436 64360 30492
rect 64296 30432 64360 30436
rect 64376 30492 64440 30496
rect 64376 30436 64380 30492
rect 64380 30436 64436 30492
rect 64436 30436 64440 30492
rect 64376 30432 64440 30436
rect 64456 30492 64520 30496
rect 64456 30436 64460 30492
rect 64460 30436 64516 30492
rect 64516 30436 64520 30492
rect 64456 30432 64520 30436
rect 9216 29948 9280 29952
rect 9216 29892 9220 29948
rect 9220 29892 9276 29948
rect 9276 29892 9280 29948
rect 9216 29888 9280 29892
rect 9296 29948 9360 29952
rect 9296 29892 9300 29948
rect 9300 29892 9356 29948
rect 9356 29892 9360 29948
rect 9296 29888 9360 29892
rect 9376 29948 9440 29952
rect 9376 29892 9380 29948
rect 9380 29892 9436 29948
rect 9436 29892 9440 29948
rect 9376 29888 9440 29892
rect 9456 29948 9520 29952
rect 9456 29892 9460 29948
rect 9460 29892 9516 29948
rect 9516 29892 9520 29948
rect 9456 29888 9520 29892
rect 19216 29948 19280 29952
rect 19216 29892 19220 29948
rect 19220 29892 19276 29948
rect 19276 29892 19280 29948
rect 19216 29888 19280 29892
rect 19296 29948 19360 29952
rect 19296 29892 19300 29948
rect 19300 29892 19356 29948
rect 19356 29892 19360 29948
rect 19296 29888 19360 29892
rect 19376 29948 19440 29952
rect 19376 29892 19380 29948
rect 19380 29892 19436 29948
rect 19436 29892 19440 29948
rect 19376 29888 19440 29892
rect 19456 29948 19520 29952
rect 19456 29892 19460 29948
rect 19460 29892 19516 29948
rect 19516 29892 19520 29948
rect 19456 29888 19520 29892
rect 29216 29948 29280 29952
rect 29216 29892 29220 29948
rect 29220 29892 29276 29948
rect 29276 29892 29280 29948
rect 29216 29888 29280 29892
rect 29296 29948 29360 29952
rect 29296 29892 29300 29948
rect 29300 29892 29356 29948
rect 29356 29892 29360 29948
rect 29296 29888 29360 29892
rect 29376 29948 29440 29952
rect 29376 29892 29380 29948
rect 29380 29892 29436 29948
rect 29436 29892 29440 29948
rect 29376 29888 29440 29892
rect 29456 29948 29520 29952
rect 29456 29892 29460 29948
rect 29460 29892 29516 29948
rect 29516 29892 29520 29948
rect 29456 29888 29520 29892
rect 39216 29948 39280 29952
rect 39216 29892 39220 29948
rect 39220 29892 39276 29948
rect 39276 29892 39280 29948
rect 39216 29888 39280 29892
rect 39296 29948 39360 29952
rect 39296 29892 39300 29948
rect 39300 29892 39356 29948
rect 39356 29892 39360 29948
rect 39296 29888 39360 29892
rect 39376 29948 39440 29952
rect 39376 29892 39380 29948
rect 39380 29892 39436 29948
rect 39436 29892 39440 29948
rect 39376 29888 39440 29892
rect 39456 29948 39520 29952
rect 39456 29892 39460 29948
rect 39460 29892 39516 29948
rect 39516 29892 39520 29948
rect 39456 29888 39520 29892
rect 49216 29948 49280 29952
rect 49216 29892 49220 29948
rect 49220 29892 49276 29948
rect 49276 29892 49280 29948
rect 49216 29888 49280 29892
rect 49296 29948 49360 29952
rect 49296 29892 49300 29948
rect 49300 29892 49356 29948
rect 49356 29892 49360 29948
rect 49296 29888 49360 29892
rect 49376 29948 49440 29952
rect 49376 29892 49380 29948
rect 49380 29892 49436 29948
rect 49436 29892 49440 29948
rect 49376 29888 49440 29892
rect 49456 29948 49520 29952
rect 49456 29892 49460 29948
rect 49460 29892 49516 29948
rect 49516 29892 49520 29948
rect 49456 29888 49520 29892
rect 59216 29948 59280 29952
rect 59216 29892 59220 29948
rect 59220 29892 59276 29948
rect 59276 29892 59280 29948
rect 59216 29888 59280 29892
rect 59296 29948 59360 29952
rect 59296 29892 59300 29948
rect 59300 29892 59356 29948
rect 59356 29892 59360 29948
rect 59296 29888 59360 29892
rect 59376 29948 59440 29952
rect 59376 29892 59380 29948
rect 59380 29892 59436 29948
rect 59436 29892 59440 29948
rect 59376 29888 59440 29892
rect 59456 29948 59520 29952
rect 59456 29892 59460 29948
rect 59460 29892 59516 29948
rect 59516 29892 59520 29948
rect 59456 29888 59520 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 14216 29404 14280 29408
rect 14216 29348 14220 29404
rect 14220 29348 14276 29404
rect 14276 29348 14280 29404
rect 14216 29344 14280 29348
rect 14296 29404 14360 29408
rect 14296 29348 14300 29404
rect 14300 29348 14356 29404
rect 14356 29348 14360 29404
rect 14296 29344 14360 29348
rect 14376 29404 14440 29408
rect 14376 29348 14380 29404
rect 14380 29348 14436 29404
rect 14436 29348 14440 29404
rect 14376 29344 14440 29348
rect 14456 29404 14520 29408
rect 14456 29348 14460 29404
rect 14460 29348 14516 29404
rect 14516 29348 14520 29404
rect 14456 29344 14520 29348
rect 24216 29404 24280 29408
rect 24216 29348 24220 29404
rect 24220 29348 24276 29404
rect 24276 29348 24280 29404
rect 24216 29344 24280 29348
rect 24296 29404 24360 29408
rect 24296 29348 24300 29404
rect 24300 29348 24356 29404
rect 24356 29348 24360 29404
rect 24296 29344 24360 29348
rect 24376 29404 24440 29408
rect 24376 29348 24380 29404
rect 24380 29348 24436 29404
rect 24436 29348 24440 29404
rect 24376 29344 24440 29348
rect 24456 29404 24520 29408
rect 24456 29348 24460 29404
rect 24460 29348 24516 29404
rect 24516 29348 24520 29404
rect 24456 29344 24520 29348
rect 34216 29404 34280 29408
rect 34216 29348 34220 29404
rect 34220 29348 34276 29404
rect 34276 29348 34280 29404
rect 34216 29344 34280 29348
rect 34296 29404 34360 29408
rect 34296 29348 34300 29404
rect 34300 29348 34356 29404
rect 34356 29348 34360 29404
rect 34296 29344 34360 29348
rect 34376 29404 34440 29408
rect 34376 29348 34380 29404
rect 34380 29348 34436 29404
rect 34436 29348 34440 29404
rect 34376 29344 34440 29348
rect 34456 29404 34520 29408
rect 34456 29348 34460 29404
rect 34460 29348 34516 29404
rect 34516 29348 34520 29404
rect 34456 29344 34520 29348
rect 44216 29404 44280 29408
rect 44216 29348 44220 29404
rect 44220 29348 44276 29404
rect 44276 29348 44280 29404
rect 44216 29344 44280 29348
rect 44296 29404 44360 29408
rect 44296 29348 44300 29404
rect 44300 29348 44356 29404
rect 44356 29348 44360 29404
rect 44296 29344 44360 29348
rect 44376 29404 44440 29408
rect 44376 29348 44380 29404
rect 44380 29348 44436 29404
rect 44436 29348 44440 29404
rect 44376 29344 44440 29348
rect 44456 29404 44520 29408
rect 44456 29348 44460 29404
rect 44460 29348 44516 29404
rect 44516 29348 44520 29404
rect 44456 29344 44520 29348
rect 54216 29404 54280 29408
rect 54216 29348 54220 29404
rect 54220 29348 54276 29404
rect 54276 29348 54280 29404
rect 54216 29344 54280 29348
rect 54296 29404 54360 29408
rect 54296 29348 54300 29404
rect 54300 29348 54356 29404
rect 54356 29348 54360 29404
rect 54296 29344 54360 29348
rect 54376 29404 54440 29408
rect 54376 29348 54380 29404
rect 54380 29348 54436 29404
rect 54436 29348 54440 29404
rect 54376 29344 54440 29348
rect 54456 29404 54520 29408
rect 54456 29348 54460 29404
rect 54460 29348 54516 29404
rect 54516 29348 54520 29404
rect 54456 29344 54520 29348
rect 64216 29404 64280 29408
rect 64216 29348 64220 29404
rect 64220 29348 64276 29404
rect 64276 29348 64280 29404
rect 64216 29344 64280 29348
rect 64296 29404 64360 29408
rect 64296 29348 64300 29404
rect 64300 29348 64356 29404
rect 64356 29348 64360 29404
rect 64296 29344 64360 29348
rect 64376 29404 64440 29408
rect 64376 29348 64380 29404
rect 64380 29348 64436 29404
rect 64436 29348 64440 29404
rect 64376 29344 64440 29348
rect 64456 29404 64520 29408
rect 64456 29348 64460 29404
rect 64460 29348 64516 29404
rect 64516 29348 64520 29404
rect 64456 29344 64520 29348
rect 9216 28860 9280 28864
rect 9216 28804 9220 28860
rect 9220 28804 9276 28860
rect 9276 28804 9280 28860
rect 9216 28800 9280 28804
rect 9296 28860 9360 28864
rect 9296 28804 9300 28860
rect 9300 28804 9356 28860
rect 9356 28804 9360 28860
rect 9296 28800 9360 28804
rect 9376 28860 9440 28864
rect 9376 28804 9380 28860
rect 9380 28804 9436 28860
rect 9436 28804 9440 28860
rect 9376 28800 9440 28804
rect 9456 28860 9520 28864
rect 9456 28804 9460 28860
rect 9460 28804 9516 28860
rect 9516 28804 9520 28860
rect 9456 28800 9520 28804
rect 19216 28860 19280 28864
rect 19216 28804 19220 28860
rect 19220 28804 19276 28860
rect 19276 28804 19280 28860
rect 19216 28800 19280 28804
rect 19296 28860 19360 28864
rect 19296 28804 19300 28860
rect 19300 28804 19356 28860
rect 19356 28804 19360 28860
rect 19296 28800 19360 28804
rect 19376 28860 19440 28864
rect 19376 28804 19380 28860
rect 19380 28804 19436 28860
rect 19436 28804 19440 28860
rect 19376 28800 19440 28804
rect 19456 28860 19520 28864
rect 19456 28804 19460 28860
rect 19460 28804 19516 28860
rect 19516 28804 19520 28860
rect 19456 28800 19520 28804
rect 29216 28860 29280 28864
rect 29216 28804 29220 28860
rect 29220 28804 29276 28860
rect 29276 28804 29280 28860
rect 29216 28800 29280 28804
rect 29296 28860 29360 28864
rect 29296 28804 29300 28860
rect 29300 28804 29356 28860
rect 29356 28804 29360 28860
rect 29296 28800 29360 28804
rect 29376 28860 29440 28864
rect 29376 28804 29380 28860
rect 29380 28804 29436 28860
rect 29436 28804 29440 28860
rect 29376 28800 29440 28804
rect 29456 28860 29520 28864
rect 29456 28804 29460 28860
rect 29460 28804 29516 28860
rect 29516 28804 29520 28860
rect 29456 28800 29520 28804
rect 39216 28860 39280 28864
rect 39216 28804 39220 28860
rect 39220 28804 39276 28860
rect 39276 28804 39280 28860
rect 39216 28800 39280 28804
rect 39296 28860 39360 28864
rect 39296 28804 39300 28860
rect 39300 28804 39356 28860
rect 39356 28804 39360 28860
rect 39296 28800 39360 28804
rect 39376 28860 39440 28864
rect 39376 28804 39380 28860
rect 39380 28804 39436 28860
rect 39436 28804 39440 28860
rect 39376 28800 39440 28804
rect 39456 28860 39520 28864
rect 39456 28804 39460 28860
rect 39460 28804 39516 28860
rect 39516 28804 39520 28860
rect 39456 28800 39520 28804
rect 49216 28860 49280 28864
rect 49216 28804 49220 28860
rect 49220 28804 49276 28860
rect 49276 28804 49280 28860
rect 49216 28800 49280 28804
rect 49296 28860 49360 28864
rect 49296 28804 49300 28860
rect 49300 28804 49356 28860
rect 49356 28804 49360 28860
rect 49296 28800 49360 28804
rect 49376 28860 49440 28864
rect 49376 28804 49380 28860
rect 49380 28804 49436 28860
rect 49436 28804 49440 28860
rect 49376 28800 49440 28804
rect 49456 28860 49520 28864
rect 49456 28804 49460 28860
rect 49460 28804 49516 28860
rect 49516 28804 49520 28860
rect 49456 28800 49520 28804
rect 59216 28860 59280 28864
rect 59216 28804 59220 28860
rect 59220 28804 59276 28860
rect 59276 28804 59280 28860
rect 59216 28800 59280 28804
rect 59296 28860 59360 28864
rect 59296 28804 59300 28860
rect 59300 28804 59356 28860
rect 59356 28804 59360 28860
rect 59296 28800 59360 28804
rect 59376 28860 59440 28864
rect 59376 28804 59380 28860
rect 59380 28804 59436 28860
rect 59436 28804 59440 28860
rect 59376 28800 59440 28804
rect 59456 28860 59520 28864
rect 59456 28804 59460 28860
rect 59460 28804 59516 28860
rect 59516 28804 59520 28860
rect 59456 28800 59520 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 14216 28316 14280 28320
rect 14216 28260 14220 28316
rect 14220 28260 14276 28316
rect 14276 28260 14280 28316
rect 14216 28256 14280 28260
rect 14296 28316 14360 28320
rect 14296 28260 14300 28316
rect 14300 28260 14356 28316
rect 14356 28260 14360 28316
rect 14296 28256 14360 28260
rect 14376 28316 14440 28320
rect 14376 28260 14380 28316
rect 14380 28260 14436 28316
rect 14436 28260 14440 28316
rect 14376 28256 14440 28260
rect 14456 28316 14520 28320
rect 14456 28260 14460 28316
rect 14460 28260 14516 28316
rect 14516 28260 14520 28316
rect 14456 28256 14520 28260
rect 24216 28316 24280 28320
rect 24216 28260 24220 28316
rect 24220 28260 24276 28316
rect 24276 28260 24280 28316
rect 24216 28256 24280 28260
rect 24296 28316 24360 28320
rect 24296 28260 24300 28316
rect 24300 28260 24356 28316
rect 24356 28260 24360 28316
rect 24296 28256 24360 28260
rect 24376 28316 24440 28320
rect 24376 28260 24380 28316
rect 24380 28260 24436 28316
rect 24436 28260 24440 28316
rect 24376 28256 24440 28260
rect 24456 28316 24520 28320
rect 24456 28260 24460 28316
rect 24460 28260 24516 28316
rect 24516 28260 24520 28316
rect 24456 28256 24520 28260
rect 34216 28316 34280 28320
rect 34216 28260 34220 28316
rect 34220 28260 34276 28316
rect 34276 28260 34280 28316
rect 34216 28256 34280 28260
rect 34296 28316 34360 28320
rect 34296 28260 34300 28316
rect 34300 28260 34356 28316
rect 34356 28260 34360 28316
rect 34296 28256 34360 28260
rect 34376 28316 34440 28320
rect 34376 28260 34380 28316
rect 34380 28260 34436 28316
rect 34436 28260 34440 28316
rect 34376 28256 34440 28260
rect 34456 28316 34520 28320
rect 34456 28260 34460 28316
rect 34460 28260 34516 28316
rect 34516 28260 34520 28316
rect 34456 28256 34520 28260
rect 44216 28316 44280 28320
rect 44216 28260 44220 28316
rect 44220 28260 44276 28316
rect 44276 28260 44280 28316
rect 44216 28256 44280 28260
rect 44296 28316 44360 28320
rect 44296 28260 44300 28316
rect 44300 28260 44356 28316
rect 44356 28260 44360 28316
rect 44296 28256 44360 28260
rect 44376 28316 44440 28320
rect 44376 28260 44380 28316
rect 44380 28260 44436 28316
rect 44436 28260 44440 28316
rect 44376 28256 44440 28260
rect 44456 28316 44520 28320
rect 44456 28260 44460 28316
rect 44460 28260 44516 28316
rect 44516 28260 44520 28316
rect 44456 28256 44520 28260
rect 54216 28316 54280 28320
rect 54216 28260 54220 28316
rect 54220 28260 54276 28316
rect 54276 28260 54280 28316
rect 54216 28256 54280 28260
rect 54296 28316 54360 28320
rect 54296 28260 54300 28316
rect 54300 28260 54356 28316
rect 54356 28260 54360 28316
rect 54296 28256 54360 28260
rect 54376 28316 54440 28320
rect 54376 28260 54380 28316
rect 54380 28260 54436 28316
rect 54436 28260 54440 28316
rect 54376 28256 54440 28260
rect 54456 28316 54520 28320
rect 54456 28260 54460 28316
rect 54460 28260 54516 28316
rect 54516 28260 54520 28316
rect 54456 28256 54520 28260
rect 64216 28316 64280 28320
rect 64216 28260 64220 28316
rect 64220 28260 64276 28316
rect 64276 28260 64280 28316
rect 64216 28256 64280 28260
rect 64296 28316 64360 28320
rect 64296 28260 64300 28316
rect 64300 28260 64356 28316
rect 64356 28260 64360 28316
rect 64296 28256 64360 28260
rect 64376 28316 64440 28320
rect 64376 28260 64380 28316
rect 64380 28260 64436 28316
rect 64436 28260 64440 28316
rect 64376 28256 64440 28260
rect 64456 28316 64520 28320
rect 64456 28260 64460 28316
rect 64460 28260 64516 28316
rect 64516 28260 64520 28316
rect 64456 28256 64520 28260
rect 9216 27772 9280 27776
rect 9216 27716 9220 27772
rect 9220 27716 9276 27772
rect 9276 27716 9280 27772
rect 9216 27712 9280 27716
rect 9296 27772 9360 27776
rect 9296 27716 9300 27772
rect 9300 27716 9356 27772
rect 9356 27716 9360 27772
rect 9296 27712 9360 27716
rect 9376 27772 9440 27776
rect 9376 27716 9380 27772
rect 9380 27716 9436 27772
rect 9436 27716 9440 27772
rect 9376 27712 9440 27716
rect 9456 27772 9520 27776
rect 9456 27716 9460 27772
rect 9460 27716 9516 27772
rect 9516 27716 9520 27772
rect 9456 27712 9520 27716
rect 19216 27772 19280 27776
rect 19216 27716 19220 27772
rect 19220 27716 19276 27772
rect 19276 27716 19280 27772
rect 19216 27712 19280 27716
rect 19296 27772 19360 27776
rect 19296 27716 19300 27772
rect 19300 27716 19356 27772
rect 19356 27716 19360 27772
rect 19296 27712 19360 27716
rect 19376 27772 19440 27776
rect 19376 27716 19380 27772
rect 19380 27716 19436 27772
rect 19436 27716 19440 27772
rect 19376 27712 19440 27716
rect 19456 27772 19520 27776
rect 19456 27716 19460 27772
rect 19460 27716 19516 27772
rect 19516 27716 19520 27772
rect 19456 27712 19520 27716
rect 29216 27772 29280 27776
rect 29216 27716 29220 27772
rect 29220 27716 29276 27772
rect 29276 27716 29280 27772
rect 29216 27712 29280 27716
rect 29296 27772 29360 27776
rect 29296 27716 29300 27772
rect 29300 27716 29356 27772
rect 29356 27716 29360 27772
rect 29296 27712 29360 27716
rect 29376 27772 29440 27776
rect 29376 27716 29380 27772
rect 29380 27716 29436 27772
rect 29436 27716 29440 27772
rect 29376 27712 29440 27716
rect 29456 27772 29520 27776
rect 29456 27716 29460 27772
rect 29460 27716 29516 27772
rect 29516 27716 29520 27772
rect 29456 27712 29520 27716
rect 39216 27772 39280 27776
rect 39216 27716 39220 27772
rect 39220 27716 39276 27772
rect 39276 27716 39280 27772
rect 39216 27712 39280 27716
rect 39296 27772 39360 27776
rect 39296 27716 39300 27772
rect 39300 27716 39356 27772
rect 39356 27716 39360 27772
rect 39296 27712 39360 27716
rect 39376 27772 39440 27776
rect 39376 27716 39380 27772
rect 39380 27716 39436 27772
rect 39436 27716 39440 27772
rect 39376 27712 39440 27716
rect 39456 27772 39520 27776
rect 39456 27716 39460 27772
rect 39460 27716 39516 27772
rect 39516 27716 39520 27772
rect 39456 27712 39520 27716
rect 49216 27772 49280 27776
rect 49216 27716 49220 27772
rect 49220 27716 49276 27772
rect 49276 27716 49280 27772
rect 49216 27712 49280 27716
rect 49296 27772 49360 27776
rect 49296 27716 49300 27772
rect 49300 27716 49356 27772
rect 49356 27716 49360 27772
rect 49296 27712 49360 27716
rect 49376 27772 49440 27776
rect 49376 27716 49380 27772
rect 49380 27716 49436 27772
rect 49436 27716 49440 27772
rect 49376 27712 49440 27716
rect 49456 27772 49520 27776
rect 49456 27716 49460 27772
rect 49460 27716 49516 27772
rect 49516 27716 49520 27772
rect 49456 27712 49520 27716
rect 59216 27772 59280 27776
rect 59216 27716 59220 27772
rect 59220 27716 59276 27772
rect 59276 27716 59280 27772
rect 59216 27712 59280 27716
rect 59296 27772 59360 27776
rect 59296 27716 59300 27772
rect 59300 27716 59356 27772
rect 59356 27716 59360 27772
rect 59296 27712 59360 27716
rect 59376 27772 59440 27776
rect 59376 27716 59380 27772
rect 59380 27716 59436 27772
rect 59436 27716 59440 27772
rect 59376 27712 59440 27716
rect 59456 27772 59520 27776
rect 59456 27716 59460 27772
rect 59460 27716 59516 27772
rect 59516 27716 59520 27772
rect 59456 27712 59520 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 14216 27228 14280 27232
rect 14216 27172 14220 27228
rect 14220 27172 14276 27228
rect 14276 27172 14280 27228
rect 14216 27168 14280 27172
rect 14296 27228 14360 27232
rect 14296 27172 14300 27228
rect 14300 27172 14356 27228
rect 14356 27172 14360 27228
rect 14296 27168 14360 27172
rect 14376 27228 14440 27232
rect 14376 27172 14380 27228
rect 14380 27172 14436 27228
rect 14436 27172 14440 27228
rect 14376 27168 14440 27172
rect 14456 27228 14520 27232
rect 14456 27172 14460 27228
rect 14460 27172 14516 27228
rect 14516 27172 14520 27228
rect 14456 27168 14520 27172
rect 24216 27228 24280 27232
rect 24216 27172 24220 27228
rect 24220 27172 24276 27228
rect 24276 27172 24280 27228
rect 24216 27168 24280 27172
rect 24296 27228 24360 27232
rect 24296 27172 24300 27228
rect 24300 27172 24356 27228
rect 24356 27172 24360 27228
rect 24296 27168 24360 27172
rect 24376 27228 24440 27232
rect 24376 27172 24380 27228
rect 24380 27172 24436 27228
rect 24436 27172 24440 27228
rect 24376 27168 24440 27172
rect 24456 27228 24520 27232
rect 24456 27172 24460 27228
rect 24460 27172 24516 27228
rect 24516 27172 24520 27228
rect 24456 27168 24520 27172
rect 34216 27228 34280 27232
rect 34216 27172 34220 27228
rect 34220 27172 34276 27228
rect 34276 27172 34280 27228
rect 34216 27168 34280 27172
rect 34296 27228 34360 27232
rect 34296 27172 34300 27228
rect 34300 27172 34356 27228
rect 34356 27172 34360 27228
rect 34296 27168 34360 27172
rect 34376 27228 34440 27232
rect 34376 27172 34380 27228
rect 34380 27172 34436 27228
rect 34436 27172 34440 27228
rect 34376 27168 34440 27172
rect 34456 27228 34520 27232
rect 34456 27172 34460 27228
rect 34460 27172 34516 27228
rect 34516 27172 34520 27228
rect 34456 27168 34520 27172
rect 44216 27228 44280 27232
rect 44216 27172 44220 27228
rect 44220 27172 44276 27228
rect 44276 27172 44280 27228
rect 44216 27168 44280 27172
rect 44296 27228 44360 27232
rect 44296 27172 44300 27228
rect 44300 27172 44356 27228
rect 44356 27172 44360 27228
rect 44296 27168 44360 27172
rect 44376 27228 44440 27232
rect 44376 27172 44380 27228
rect 44380 27172 44436 27228
rect 44436 27172 44440 27228
rect 44376 27168 44440 27172
rect 44456 27228 44520 27232
rect 44456 27172 44460 27228
rect 44460 27172 44516 27228
rect 44516 27172 44520 27228
rect 44456 27168 44520 27172
rect 54216 27228 54280 27232
rect 54216 27172 54220 27228
rect 54220 27172 54276 27228
rect 54276 27172 54280 27228
rect 54216 27168 54280 27172
rect 54296 27228 54360 27232
rect 54296 27172 54300 27228
rect 54300 27172 54356 27228
rect 54356 27172 54360 27228
rect 54296 27168 54360 27172
rect 54376 27228 54440 27232
rect 54376 27172 54380 27228
rect 54380 27172 54436 27228
rect 54436 27172 54440 27228
rect 54376 27168 54440 27172
rect 54456 27228 54520 27232
rect 54456 27172 54460 27228
rect 54460 27172 54516 27228
rect 54516 27172 54520 27228
rect 54456 27168 54520 27172
rect 64216 27228 64280 27232
rect 64216 27172 64220 27228
rect 64220 27172 64276 27228
rect 64276 27172 64280 27228
rect 64216 27168 64280 27172
rect 64296 27228 64360 27232
rect 64296 27172 64300 27228
rect 64300 27172 64356 27228
rect 64356 27172 64360 27228
rect 64296 27168 64360 27172
rect 64376 27228 64440 27232
rect 64376 27172 64380 27228
rect 64380 27172 64436 27228
rect 64436 27172 64440 27228
rect 64376 27168 64440 27172
rect 64456 27228 64520 27232
rect 64456 27172 64460 27228
rect 64460 27172 64516 27228
rect 64516 27172 64520 27228
rect 64456 27168 64520 27172
rect 9216 26684 9280 26688
rect 9216 26628 9220 26684
rect 9220 26628 9276 26684
rect 9276 26628 9280 26684
rect 9216 26624 9280 26628
rect 9296 26684 9360 26688
rect 9296 26628 9300 26684
rect 9300 26628 9356 26684
rect 9356 26628 9360 26684
rect 9296 26624 9360 26628
rect 9376 26684 9440 26688
rect 9376 26628 9380 26684
rect 9380 26628 9436 26684
rect 9436 26628 9440 26684
rect 9376 26624 9440 26628
rect 9456 26684 9520 26688
rect 9456 26628 9460 26684
rect 9460 26628 9516 26684
rect 9516 26628 9520 26684
rect 9456 26624 9520 26628
rect 19216 26684 19280 26688
rect 19216 26628 19220 26684
rect 19220 26628 19276 26684
rect 19276 26628 19280 26684
rect 19216 26624 19280 26628
rect 19296 26684 19360 26688
rect 19296 26628 19300 26684
rect 19300 26628 19356 26684
rect 19356 26628 19360 26684
rect 19296 26624 19360 26628
rect 19376 26684 19440 26688
rect 19376 26628 19380 26684
rect 19380 26628 19436 26684
rect 19436 26628 19440 26684
rect 19376 26624 19440 26628
rect 19456 26684 19520 26688
rect 19456 26628 19460 26684
rect 19460 26628 19516 26684
rect 19516 26628 19520 26684
rect 19456 26624 19520 26628
rect 29216 26684 29280 26688
rect 29216 26628 29220 26684
rect 29220 26628 29276 26684
rect 29276 26628 29280 26684
rect 29216 26624 29280 26628
rect 29296 26684 29360 26688
rect 29296 26628 29300 26684
rect 29300 26628 29356 26684
rect 29356 26628 29360 26684
rect 29296 26624 29360 26628
rect 29376 26684 29440 26688
rect 29376 26628 29380 26684
rect 29380 26628 29436 26684
rect 29436 26628 29440 26684
rect 29376 26624 29440 26628
rect 29456 26684 29520 26688
rect 29456 26628 29460 26684
rect 29460 26628 29516 26684
rect 29516 26628 29520 26684
rect 29456 26624 29520 26628
rect 39216 26684 39280 26688
rect 39216 26628 39220 26684
rect 39220 26628 39276 26684
rect 39276 26628 39280 26684
rect 39216 26624 39280 26628
rect 39296 26684 39360 26688
rect 39296 26628 39300 26684
rect 39300 26628 39356 26684
rect 39356 26628 39360 26684
rect 39296 26624 39360 26628
rect 39376 26684 39440 26688
rect 39376 26628 39380 26684
rect 39380 26628 39436 26684
rect 39436 26628 39440 26684
rect 39376 26624 39440 26628
rect 39456 26684 39520 26688
rect 39456 26628 39460 26684
rect 39460 26628 39516 26684
rect 39516 26628 39520 26684
rect 39456 26624 39520 26628
rect 49216 26684 49280 26688
rect 49216 26628 49220 26684
rect 49220 26628 49276 26684
rect 49276 26628 49280 26684
rect 49216 26624 49280 26628
rect 49296 26684 49360 26688
rect 49296 26628 49300 26684
rect 49300 26628 49356 26684
rect 49356 26628 49360 26684
rect 49296 26624 49360 26628
rect 49376 26684 49440 26688
rect 49376 26628 49380 26684
rect 49380 26628 49436 26684
rect 49436 26628 49440 26684
rect 49376 26624 49440 26628
rect 49456 26684 49520 26688
rect 49456 26628 49460 26684
rect 49460 26628 49516 26684
rect 49516 26628 49520 26684
rect 49456 26624 49520 26628
rect 59216 26684 59280 26688
rect 59216 26628 59220 26684
rect 59220 26628 59276 26684
rect 59276 26628 59280 26684
rect 59216 26624 59280 26628
rect 59296 26684 59360 26688
rect 59296 26628 59300 26684
rect 59300 26628 59356 26684
rect 59356 26628 59360 26684
rect 59296 26624 59360 26628
rect 59376 26684 59440 26688
rect 59376 26628 59380 26684
rect 59380 26628 59436 26684
rect 59436 26628 59440 26684
rect 59376 26624 59440 26628
rect 59456 26684 59520 26688
rect 59456 26628 59460 26684
rect 59460 26628 59516 26684
rect 59516 26628 59520 26684
rect 59456 26624 59520 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 14216 26140 14280 26144
rect 14216 26084 14220 26140
rect 14220 26084 14276 26140
rect 14276 26084 14280 26140
rect 14216 26080 14280 26084
rect 14296 26140 14360 26144
rect 14296 26084 14300 26140
rect 14300 26084 14356 26140
rect 14356 26084 14360 26140
rect 14296 26080 14360 26084
rect 14376 26140 14440 26144
rect 14376 26084 14380 26140
rect 14380 26084 14436 26140
rect 14436 26084 14440 26140
rect 14376 26080 14440 26084
rect 14456 26140 14520 26144
rect 14456 26084 14460 26140
rect 14460 26084 14516 26140
rect 14516 26084 14520 26140
rect 14456 26080 14520 26084
rect 24216 26140 24280 26144
rect 24216 26084 24220 26140
rect 24220 26084 24276 26140
rect 24276 26084 24280 26140
rect 24216 26080 24280 26084
rect 24296 26140 24360 26144
rect 24296 26084 24300 26140
rect 24300 26084 24356 26140
rect 24356 26084 24360 26140
rect 24296 26080 24360 26084
rect 24376 26140 24440 26144
rect 24376 26084 24380 26140
rect 24380 26084 24436 26140
rect 24436 26084 24440 26140
rect 24376 26080 24440 26084
rect 24456 26140 24520 26144
rect 24456 26084 24460 26140
rect 24460 26084 24516 26140
rect 24516 26084 24520 26140
rect 24456 26080 24520 26084
rect 34216 26140 34280 26144
rect 34216 26084 34220 26140
rect 34220 26084 34276 26140
rect 34276 26084 34280 26140
rect 34216 26080 34280 26084
rect 34296 26140 34360 26144
rect 34296 26084 34300 26140
rect 34300 26084 34356 26140
rect 34356 26084 34360 26140
rect 34296 26080 34360 26084
rect 34376 26140 34440 26144
rect 34376 26084 34380 26140
rect 34380 26084 34436 26140
rect 34436 26084 34440 26140
rect 34376 26080 34440 26084
rect 34456 26140 34520 26144
rect 34456 26084 34460 26140
rect 34460 26084 34516 26140
rect 34516 26084 34520 26140
rect 34456 26080 34520 26084
rect 44216 26140 44280 26144
rect 44216 26084 44220 26140
rect 44220 26084 44276 26140
rect 44276 26084 44280 26140
rect 44216 26080 44280 26084
rect 44296 26140 44360 26144
rect 44296 26084 44300 26140
rect 44300 26084 44356 26140
rect 44356 26084 44360 26140
rect 44296 26080 44360 26084
rect 44376 26140 44440 26144
rect 44376 26084 44380 26140
rect 44380 26084 44436 26140
rect 44436 26084 44440 26140
rect 44376 26080 44440 26084
rect 44456 26140 44520 26144
rect 44456 26084 44460 26140
rect 44460 26084 44516 26140
rect 44516 26084 44520 26140
rect 44456 26080 44520 26084
rect 54216 26140 54280 26144
rect 54216 26084 54220 26140
rect 54220 26084 54276 26140
rect 54276 26084 54280 26140
rect 54216 26080 54280 26084
rect 54296 26140 54360 26144
rect 54296 26084 54300 26140
rect 54300 26084 54356 26140
rect 54356 26084 54360 26140
rect 54296 26080 54360 26084
rect 54376 26140 54440 26144
rect 54376 26084 54380 26140
rect 54380 26084 54436 26140
rect 54436 26084 54440 26140
rect 54376 26080 54440 26084
rect 54456 26140 54520 26144
rect 54456 26084 54460 26140
rect 54460 26084 54516 26140
rect 54516 26084 54520 26140
rect 54456 26080 54520 26084
rect 64216 26140 64280 26144
rect 64216 26084 64220 26140
rect 64220 26084 64276 26140
rect 64276 26084 64280 26140
rect 64216 26080 64280 26084
rect 64296 26140 64360 26144
rect 64296 26084 64300 26140
rect 64300 26084 64356 26140
rect 64356 26084 64360 26140
rect 64296 26080 64360 26084
rect 64376 26140 64440 26144
rect 64376 26084 64380 26140
rect 64380 26084 64436 26140
rect 64436 26084 64440 26140
rect 64376 26080 64440 26084
rect 64456 26140 64520 26144
rect 64456 26084 64460 26140
rect 64460 26084 64516 26140
rect 64516 26084 64520 26140
rect 64456 26080 64520 26084
rect 9216 25596 9280 25600
rect 9216 25540 9220 25596
rect 9220 25540 9276 25596
rect 9276 25540 9280 25596
rect 9216 25536 9280 25540
rect 9296 25596 9360 25600
rect 9296 25540 9300 25596
rect 9300 25540 9356 25596
rect 9356 25540 9360 25596
rect 9296 25536 9360 25540
rect 9376 25596 9440 25600
rect 9376 25540 9380 25596
rect 9380 25540 9436 25596
rect 9436 25540 9440 25596
rect 9376 25536 9440 25540
rect 9456 25596 9520 25600
rect 9456 25540 9460 25596
rect 9460 25540 9516 25596
rect 9516 25540 9520 25596
rect 9456 25536 9520 25540
rect 19216 25596 19280 25600
rect 19216 25540 19220 25596
rect 19220 25540 19276 25596
rect 19276 25540 19280 25596
rect 19216 25536 19280 25540
rect 19296 25596 19360 25600
rect 19296 25540 19300 25596
rect 19300 25540 19356 25596
rect 19356 25540 19360 25596
rect 19296 25536 19360 25540
rect 19376 25596 19440 25600
rect 19376 25540 19380 25596
rect 19380 25540 19436 25596
rect 19436 25540 19440 25596
rect 19376 25536 19440 25540
rect 19456 25596 19520 25600
rect 19456 25540 19460 25596
rect 19460 25540 19516 25596
rect 19516 25540 19520 25596
rect 19456 25536 19520 25540
rect 29216 25596 29280 25600
rect 29216 25540 29220 25596
rect 29220 25540 29276 25596
rect 29276 25540 29280 25596
rect 29216 25536 29280 25540
rect 29296 25596 29360 25600
rect 29296 25540 29300 25596
rect 29300 25540 29356 25596
rect 29356 25540 29360 25596
rect 29296 25536 29360 25540
rect 29376 25596 29440 25600
rect 29376 25540 29380 25596
rect 29380 25540 29436 25596
rect 29436 25540 29440 25596
rect 29376 25536 29440 25540
rect 29456 25596 29520 25600
rect 29456 25540 29460 25596
rect 29460 25540 29516 25596
rect 29516 25540 29520 25596
rect 29456 25536 29520 25540
rect 39216 25596 39280 25600
rect 39216 25540 39220 25596
rect 39220 25540 39276 25596
rect 39276 25540 39280 25596
rect 39216 25536 39280 25540
rect 39296 25596 39360 25600
rect 39296 25540 39300 25596
rect 39300 25540 39356 25596
rect 39356 25540 39360 25596
rect 39296 25536 39360 25540
rect 39376 25596 39440 25600
rect 39376 25540 39380 25596
rect 39380 25540 39436 25596
rect 39436 25540 39440 25596
rect 39376 25536 39440 25540
rect 39456 25596 39520 25600
rect 39456 25540 39460 25596
rect 39460 25540 39516 25596
rect 39516 25540 39520 25596
rect 39456 25536 39520 25540
rect 49216 25596 49280 25600
rect 49216 25540 49220 25596
rect 49220 25540 49276 25596
rect 49276 25540 49280 25596
rect 49216 25536 49280 25540
rect 49296 25596 49360 25600
rect 49296 25540 49300 25596
rect 49300 25540 49356 25596
rect 49356 25540 49360 25596
rect 49296 25536 49360 25540
rect 49376 25596 49440 25600
rect 49376 25540 49380 25596
rect 49380 25540 49436 25596
rect 49436 25540 49440 25596
rect 49376 25536 49440 25540
rect 49456 25596 49520 25600
rect 49456 25540 49460 25596
rect 49460 25540 49516 25596
rect 49516 25540 49520 25596
rect 49456 25536 49520 25540
rect 59216 25596 59280 25600
rect 59216 25540 59220 25596
rect 59220 25540 59276 25596
rect 59276 25540 59280 25596
rect 59216 25536 59280 25540
rect 59296 25596 59360 25600
rect 59296 25540 59300 25596
rect 59300 25540 59356 25596
rect 59356 25540 59360 25596
rect 59296 25536 59360 25540
rect 59376 25596 59440 25600
rect 59376 25540 59380 25596
rect 59380 25540 59436 25596
rect 59436 25540 59440 25596
rect 59376 25536 59440 25540
rect 59456 25596 59520 25600
rect 59456 25540 59460 25596
rect 59460 25540 59516 25596
rect 59516 25540 59520 25596
rect 59456 25536 59520 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 14216 25052 14280 25056
rect 14216 24996 14220 25052
rect 14220 24996 14276 25052
rect 14276 24996 14280 25052
rect 14216 24992 14280 24996
rect 14296 25052 14360 25056
rect 14296 24996 14300 25052
rect 14300 24996 14356 25052
rect 14356 24996 14360 25052
rect 14296 24992 14360 24996
rect 14376 25052 14440 25056
rect 14376 24996 14380 25052
rect 14380 24996 14436 25052
rect 14436 24996 14440 25052
rect 14376 24992 14440 24996
rect 14456 25052 14520 25056
rect 14456 24996 14460 25052
rect 14460 24996 14516 25052
rect 14516 24996 14520 25052
rect 14456 24992 14520 24996
rect 24216 25052 24280 25056
rect 24216 24996 24220 25052
rect 24220 24996 24276 25052
rect 24276 24996 24280 25052
rect 24216 24992 24280 24996
rect 24296 25052 24360 25056
rect 24296 24996 24300 25052
rect 24300 24996 24356 25052
rect 24356 24996 24360 25052
rect 24296 24992 24360 24996
rect 24376 25052 24440 25056
rect 24376 24996 24380 25052
rect 24380 24996 24436 25052
rect 24436 24996 24440 25052
rect 24376 24992 24440 24996
rect 24456 25052 24520 25056
rect 24456 24996 24460 25052
rect 24460 24996 24516 25052
rect 24516 24996 24520 25052
rect 24456 24992 24520 24996
rect 34216 25052 34280 25056
rect 34216 24996 34220 25052
rect 34220 24996 34276 25052
rect 34276 24996 34280 25052
rect 34216 24992 34280 24996
rect 34296 25052 34360 25056
rect 34296 24996 34300 25052
rect 34300 24996 34356 25052
rect 34356 24996 34360 25052
rect 34296 24992 34360 24996
rect 34376 25052 34440 25056
rect 34376 24996 34380 25052
rect 34380 24996 34436 25052
rect 34436 24996 34440 25052
rect 34376 24992 34440 24996
rect 34456 25052 34520 25056
rect 34456 24996 34460 25052
rect 34460 24996 34516 25052
rect 34516 24996 34520 25052
rect 34456 24992 34520 24996
rect 44216 25052 44280 25056
rect 44216 24996 44220 25052
rect 44220 24996 44276 25052
rect 44276 24996 44280 25052
rect 44216 24992 44280 24996
rect 44296 25052 44360 25056
rect 44296 24996 44300 25052
rect 44300 24996 44356 25052
rect 44356 24996 44360 25052
rect 44296 24992 44360 24996
rect 44376 25052 44440 25056
rect 44376 24996 44380 25052
rect 44380 24996 44436 25052
rect 44436 24996 44440 25052
rect 44376 24992 44440 24996
rect 44456 25052 44520 25056
rect 44456 24996 44460 25052
rect 44460 24996 44516 25052
rect 44516 24996 44520 25052
rect 44456 24992 44520 24996
rect 54216 25052 54280 25056
rect 54216 24996 54220 25052
rect 54220 24996 54276 25052
rect 54276 24996 54280 25052
rect 54216 24992 54280 24996
rect 54296 25052 54360 25056
rect 54296 24996 54300 25052
rect 54300 24996 54356 25052
rect 54356 24996 54360 25052
rect 54296 24992 54360 24996
rect 54376 25052 54440 25056
rect 54376 24996 54380 25052
rect 54380 24996 54436 25052
rect 54436 24996 54440 25052
rect 54376 24992 54440 24996
rect 54456 25052 54520 25056
rect 54456 24996 54460 25052
rect 54460 24996 54516 25052
rect 54516 24996 54520 25052
rect 54456 24992 54520 24996
rect 64216 25052 64280 25056
rect 64216 24996 64220 25052
rect 64220 24996 64276 25052
rect 64276 24996 64280 25052
rect 64216 24992 64280 24996
rect 64296 25052 64360 25056
rect 64296 24996 64300 25052
rect 64300 24996 64356 25052
rect 64356 24996 64360 25052
rect 64296 24992 64360 24996
rect 64376 25052 64440 25056
rect 64376 24996 64380 25052
rect 64380 24996 64436 25052
rect 64436 24996 64440 25052
rect 64376 24992 64440 24996
rect 64456 25052 64520 25056
rect 64456 24996 64460 25052
rect 64460 24996 64516 25052
rect 64516 24996 64520 25052
rect 64456 24992 64520 24996
rect 9216 24508 9280 24512
rect 9216 24452 9220 24508
rect 9220 24452 9276 24508
rect 9276 24452 9280 24508
rect 9216 24448 9280 24452
rect 9296 24508 9360 24512
rect 9296 24452 9300 24508
rect 9300 24452 9356 24508
rect 9356 24452 9360 24508
rect 9296 24448 9360 24452
rect 9376 24508 9440 24512
rect 9376 24452 9380 24508
rect 9380 24452 9436 24508
rect 9436 24452 9440 24508
rect 9376 24448 9440 24452
rect 9456 24508 9520 24512
rect 9456 24452 9460 24508
rect 9460 24452 9516 24508
rect 9516 24452 9520 24508
rect 9456 24448 9520 24452
rect 19216 24508 19280 24512
rect 19216 24452 19220 24508
rect 19220 24452 19276 24508
rect 19276 24452 19280 24508
rect 19216 24448 19280 24452
rect 19296 24508 19360 24512
rect 19296 24452 19300 24508
rect 19300 24452 19356 24508
rect 19356 24452 19360 24508
rect 19296 24448 19360 24452
rect 19376 24508 19440 24512
rect 19376 24452 19380 24508
rect 19380 24452 19436 24508
rect 19436 24452 19440 24508
rect 19376 24448 19440 24452
rect 19456 24508 19520 24512
rect 19456 24452 19460 24508
rect 19460 24452 19516 24508
rect 19516 24452 19520 24508
rect 19456 24448 19520 24452
rect 29216 24508 29280 24512
rect 29216 24452 29220 24508
rect 29220 24452 29276 24508
rect 29276 24452 29280 24508
rect 29216 24448 29280 24452
rect 29296 24508 29360 24512
rect 29296 24452 29300 24508
rect 29300 24452 29356 24508
rect 29356 24452 29360 24508
rect 29296 24448 29360 24452
rect 29376 24508 29440 24512
rect 29376 24452 29380 24508
rect 29380 24452 29436 24508
rect 29436 24452 29440 24508
rect 29376 24448 29440 24452
rect 29456 24508 29520 24512
rect 29456 24452 29460 24508
rect 29460 24452 29516 24508
rect 29516 24452 29520 24508
rect 29456 24448 29520 24452
rect 39216 24508 39280 24512
rect 39216 24452 39220 24508
rect 39220 24452 39276 24508
rect 39276 24452 39280 24508
rect 39216 24448 39280 24452
rect 39296 24508 39360 24512
rect 39296 24452 39300 24508
rect 39300 24452 39356 24508
rect 39356 24452 39360 24508
rect 39296 24448 39360 24452
rect 39376 24508 39440 24512
rect 39376 24452 39380 24508
rect 39380 24452 39436 24508
rect 39436 24452 39440 24508
rect 39376 24448 39440 24452
rect 39456 24508 39520 24512
rect 39456 24452 39460 24508
rect 39460 24452 39516 24508
rect 39516 24452 39520 24508
rect 39456 24448 39520 24452
rect 49216 24508 49280 24512
rect 49216 24452 49220 24508
rect 49220 24452 49276 24508
rect 49276 24452 49280 24508
rect 49216 24448 49280 24452
rect 49296 24508 49360 24512
rect 49296 24452 49300 24508
rect 49300 24452 49356 24508
rect 49356 24452 49360 24508
rect 49296 24448 49360 24452
rect 49376 24508 49440 24512
rect 49376 24452 49380 24508
rect 49380 24452 49436 24508
rect 49436 24452 49440 24508
rect 49376 24448 49440 24452
rect 49456 24508 49520 24512
rect 49456 24452 49460 24508
rect 49460 24452 49516 24508
rect 49516 24452 49520 24508
rect 49456 24448 49520 24452
rect 59216 24508 59280 24512
rect 59216 24452 59220 24508
rect 59220 24452 59276 24508
rect 59276 24452 59280 24508
rect 59216 24448 59280 24452
rect 59296 24508 59360 24512
rect 59296 24452 59300 24508
rect 59300 24452 59356 24508
rect 59356 24452 59360 24508
rect 59296 24448 59360 24452
rect 59376 24508 59440 24512
rect 59376 24452 59380 24508
rect 59380 24452 59436 24508
rect 59436 24452 59440 24508
rect 59376 24448 59440 24452
rect 59456 24508 59520 24512
rect 59456 24452 59460 24508
rect 59460 24452 59516 24508
rect 59516 24452 59520 24508
rect 59456 24448 59520 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 14216 23964 14280 23968
rect 14216 23908 14220 23964
rect 14220 23908 14276 23964
rect 14276 23908 14280 23964
rect 14216 23904 14280 23908
rect 14296 23964 14360 23968
rect 14296 23908 14300 23964
rect 14300 23908 14356 23964
rect 14356 23908 14360 23964
rect 14296 23904 14360 23908
rect 14376 23964 14440 23968
rect 14376 23908 14380 23964
rect 14380 23908 14436 23964
rect 14436 23908 14440 23964
rect 14376 23904 14440 23908
rect 14456 23964 14520 23968
rect 14456 23908 14460 23964
rect 14460 23908 14516 23964
rect 14516 23908 14520 23964
rect 14456 23904 14520 23908
rect 24216 23964 24280 23968
rect 24216 23908 24220 23964
rect 24220 23908 24276 23964
rect 24276 23908 24280 23964
rect 24216 23904 24280 23908
rect 24296 23964 24360 23968
rect 24296 23908 24300 23964
rect 24300 23908 24356 23964
rect 24356 23908 24360 23964
rect 24296 23904 24360 23908
rect 24376 23964 24440 23968
rect 24376 23908 24380 23964
rect 24380 23908 24436 23964
rect 24436 23908 24440 23964
rect 24376 23904 24440 23908
rect 24456 23964 24520 23968
rect 24456 23908 24460 23964
rect 24460 23908 24516 23964
rect 24516 23908 24520 23964
rect 24456 23904 24520 23908
rect 34216 23964 34280 23968
rect 34216 23908 34220 23964
rect 34220 23908 34276 23964
rect 34276 23908 34280 23964
rect 34216 23904 34280 23908
rect 34296 23964 34360 23968
rect 34296 23908 34300 23964
rect 34300 23908 34356 23964
rect 34356 23908 34360 23964
rect 34296 23904 34360 23908
rect 34376 23964 34440 23968
rect 34376 23908 34380 23964
rect 34380 23908 34436 23964
rect 34436 23908 34440 23964
rect 34376 23904 34440 23908
rect 34456 23964 34520 23968
rect 34456 23908 34460 23964
rect 34460 23908 34516 23964
rect 34516 23908 34520 23964
rect 34456 23904 34520 23908
rect 44216 23964 44280 23968
rect 44216 23908 44220 23964
rect 44220 23908 44276 23964
rect 44276 23908 44280 23964
rect 44216 23904 44280 23908
rect 44296 23964 44360 23968
rect 44296 23908 44300 23964
rect 44300 23908 44356 23964
rect 44356 23908 44360 23964
rect 44296 23904 44360 23908
rect 44376 23964 44440 23968
rect 44376 23908 44380 23964
rect 44380 23908 44436 23964
rect 44436 23908 44440 23964
rect 44376 23904 44440 23908
rect 44456 23964 44520 23968
rect 44456 23908 44460 23964
rect 44460 23908 44516 23964
rect 44516 23908 44520 23964
rect 44456 23904 44520 23908
rect 54216 23964 54280 23968
rect 54216 23908 54220 23964
rect 54220 23908 54276 23964
rect 54276 23908 54280 23964
rect 54216 23904 54280 23908
rect 54296 23964 54360 23968
rect 54296 23908 54300 23964
rect 54300 23908 54356 23964
rect 54356 23908 54360 23964
rect 54296 23904 54360 23908
rect 54376 23964 54440 23968
rect 54376 23908 54380 23964
rect 54380 23908 54436 23964
rect 54436 23908 54440 23964
rect 54376 23904 54440 23908
rect 54456 23964 54520 23968
rect 54456 23908 54460 23964
rect 54460 23908 54516 23964
rect 54516 23908 54520 23964
rect 54456 23904 54520 23908
rect 64216 23964 64280 23968
rect 64216 23908 64220 23964
rect 64220 23908 64276 23964
rect 64276 23908 64280 23964
rect 64216 23904 64280 23908
rect 64296 23964 64360 23968
rect 64296 23908 64300 23964
rect 64300 23908 64356 23964
rect 64356 23908 64360 23964
rect 64296 23904 64360 23908
rect 64376 23964 64440 23968
rect 64376 23908 64380 23964
rect 64380 23908 64436 23964
rect 64436 23908 64440 23964
rect 64376 23904 64440 23908
rect 64456 23964 64520 23968
rect 64456 23908 64460 23964
rect 64460 23908 64516 23964
rect 64516 23908 64520 23964
rect 64456 23904 64520 23908
rect 9216 23420 9280 23424
rect 9216 23364 9220 23420
rect 9220 23364 9276 23420
rect 9276 23364 9280 23420
rect 9216 23360 9280 23364
rect 9296 23420 9360 23424
rect 9296 23364 9300 23420
rect 9300 23364 9356 23420
rect 9356 23364 9360 23420
rect 9296 23360 9360 23364
rect 9376 23420 9440 23424
rect 9376 23364 9380 23420
rect 9380 23364 9436 23420
rect 9436 23364 9440 23420
rect 9376 23360 9440 23364
rect 9456 23420 9520 23424
rect 9456 23364 9460 23420
rect 9460 23364 9516 23420
rect 9516 23364 9520 23420
rect 9456 23360 9520 23364
rect 19216 23420 19280 23424
rect 19216 23364 19220 23420
rect 19220 23364 19276 23420
rect 19276 23364 19280 23420
rect 19216 23360 19280 23364
rect 19296 23420 19360 23424
rect 19296 23364 19300 23420
rect 19300 23364 19356 23420
rect 19356 23364 19360 23420
rect 19296 23360 19360 23364
rect 19376 23420 19440 23424
rect 19376 23364 19380 23420
rect 19380 23364 19436 23420
rect 19436 23364 19440 23420
rect 19376 23360 19440 23364
rect 19456 23420 19520 23424
rect 19456 23364 19460 23420
rect 19460 23364 19516 23420
rect 19516 23364 19520 23420
rect 19456 23360 19520 23364
rect 29216 23420 29280 23424
rect 29216 23364 29220 23420
rect 29220 23364 29276 23420
rect 29276 23364 29280 23420
rect 29216 23360 29280 23364
rect 29296 23420 29360 23424
rect 29296 23364 29300 23420
rect 29300 23364 29356 23420
rect 29356 23364 29360 23420
rect 29296 23360 29360 23364
rect 29376 23420 29440 23424
rect 29376 23364 29380 23420
rect 29380 23364 29436 23420
rect 29436 23364 29440 23420
rect 29376 23360 29440 23364
rect 29456 23420 29520 23424
rect 29456 23364 29460 23420
rect 29460 23364 29516 23420
rect 29516 23364 29520 23420
rect 29456 23360 29520 23364
rect 39216 23420 39280 23424
rect 39216 23364 39220 23420
rect 39220 23364 39276 23420
rect 39276 23364 39280 23420
rect 39216 23360 39280 23364
rect 39296 23420 39360 23424
rect 39296 23364 39300 23420
rect 39300 23364 39356 23420
rect 39356 23364 39360 23420
rect 39296 23360 39360 23364
rect 39376 23420 39440 23424
rect 39376 23364 39380 23420
rect 39380 23364 39436 23420
rect 39436 23364 39440 23420
rect 39376 23360 39440 23364
rect 39456 23420 39520 23424
rect 39456 23364 39460 23420
rect 39460 23364 39516 23420
rect 39516 23364 39520 23420
rect 39456 23360 39520 23364
rect 49216 23420 49280 23424
rect 49216 23364 49220 23420
rect 49220 23364 49276 23420
rect 49276 23364 49280 23420
rect 49216 23360 49280 23364
rect 49296 23420 49360 23424
rect 49296 23364 49300 23420
rect 49300 23364 49356 23420
rect 49356 23364 49360 23420
rect 49296 23360 49360 23364
rect 49376 23420 49440 23424
rect 49376 23364 49380 23420
rect 49380 23364 49436 23420
rect 49436 23364 49440 23420
rect 49376 23360 49440 23364
rect 49456 23420 49520 23424
rect 49456 23364 49460 23420
rect 49460 23364 49516 23420
rect 49516 23364 49520 23420
rect 49456 23360 49520 23364
rect 59216 23420 59280 23424
rect 59216 23364 59220 23420
rect 59220 23364 59276 23420
rect 59276 23364 59280 23420
rect 59216 23360 59280 23364
rect 59296 23420 59360 23424
rect 59296 23364 59300 23420
rect 59300 23364 59356 23420
rect 59356 23364 59360 23420
rect 59296 23360 59360 23364
rect 59376 23420 59440 23424
rect 59376 23364 59380 23420
rect 59380 23364 59436 23420
rect 59436 23364 59440 23420
rect 59376 23360 59440 23364
rect 59456 23420 59520 23424
rect 59456 23364 59460 23420
rect 59460 23364 59516 23420
rect 59516 23364 59520 23420
rect 59456 23360 59520 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 14216 22876 14280 22880
rect 14216 22820 14220 22876
rect 14220 22820 14276 22876
rect 14276 22820 14280 22876
rect 14216 22816 14280 22820
rect 14296 22876 14360 22880
rect 14296 22820 14300 22876
rect 14300 22820 14356 22876
rect 14356 22820 14360 22876
rect 14296 22816 14360 22820
rect 14376 22876 14440 22880
rect 14376 22820 14380 22876
rect 14380 22820 14436 22876
rect 14436 22820 14440 22876
rect 14376 22816 14440 22820
rect 14456 22876 14520 22880
rect 14456 22820 14460 22876
rect 14460 22820 14516 22876
rect 14516 22820 14520 22876
rect 14456 22816 14520 22820
rect 24216 22876 24280 22880
rect 24216 22820 24220 22876
rect 24220 22820 24276 22876
rect 24276 22820 24280 22876
rect 24216 22816 24280 22820
rect 24296 22876 24360 22880
rect 24296 22820 24300 22876
rect 24300 22820 24356 22876
rect 24356 22820 24360 22876
rect 24296 22816 24360 22820
rect 24376 22876 24440 22880
rect 24376 22820 24380 22876
rect 24380 22820 24436 22876
rect 24436 22820 24440 22876
rect 24376 22816 24440 22820
rect 24456 22876 24520 22880
rect 24456 22820 24460 22876
rect 24460 22820 24516 22876
rect 24516 22820 24520 22876
rect 24456 22816 24520 22820
rect 34216 22876 34280 22880
rect 34216 22820 34220 22876
rect 34220 22820 34276 22876
rect 34276 22820 34280 22876
rect 34216 22816 34280 22820
rect 34296 22876 34360 22880
rect 34296 22820 34300 22876
rect 34300 22820 34356 22876
rect 34356 22820 34360 22876
rect 34296 22816 34360 22820
rect 34376 22876 34440 22880
rect 34376 22820 34380 22876
rect 34380 22820 34436 22876
rect 34436 22820 34440 22876
rect 34376 22816 34440 22820
rect 34456 22876 34520 22880
rect 34456 22820 34460 22876
rect 34460 22820 34516 22876
rect 34516 22820 34520 22876
rect 34456 22816 34520 22820
rect 44216 22876 44280 22880
rect 44216 22820 44220 22876
rect 44220 22820 44276 22876
rect 44276 22820 44280 22876
rect 44216 22816 44280 22820
rect 44296 22876 44360 22880
rect 44296 22820 44300 22876
rect 44300 22820 44356 22876
rect 44356 22820 44360 22876
rect 44296 22816 44360 22820
rect 44376 22876 44440 22880
rect 44376 22820 44380 22876
rect 44380 22820 44436 22876
rect 44436 22820 44440 22876
rect 44376 22816 44440 22820
rect 44456 22876 44520 22880
rect 44456 22820 44460 22876
rect 44460 22820 44516 22876
rect 44516 22820 44520 22876
rect 44456 22816 44520 22820
rect 54216 22876 54280 22880
rect 54216 22820 54220 22876
rect 54220 22820 54276 22876
rect 54276 22820 54280 22876
rect 54216 22816 54280 22820
rect 54296 22876 54360 22880
rect 54296 22820 54300 22876
rect 54300 22820 54356 22876
rect 54356 22820 54360 22876
rect 54296 22816 54360 22820
rect 54376 22876 54440 22880
rect 54376 22820 54380 22876
rect 54380 22820 54436 22876
rect 54436 22820 54440 22876
rect 54376 22816 54440 22820
rect 54456 22876 54520 22880
rect 54456 22820 54460 22876
rect 54460 22820 54516 22876
rect 54516 22820 54520 22876
rect 54456 22816 54520 22820
rect 64216 22876 64280 22880
rect 64216 22820 64220 22876
rect 64220 22820 64276 22876
rect 64276 22820 64280 22876
rect 64216 22816 64280 22820
rect 64296 22876 64360 22880
rect 64296 22820 64300 22876
rect 64300 22820 64356 22876
rect 64356 22820 64360 22876
rect 64296 22816 64360 22820
rect 64376 22876 64440 22880
rect 64376 22820 64380 22876
rect 64380 22820 64436 22876
rect 64436 22820 64440 22876
rect 64376 22816 64440 22820
rect 64456 22876 64520 22880
rect 64456 22820 64460 22876
rect 64460 22820 64516 22876
rect 64516 22820 64520 22876
rect 64456 22816 64520 22820
rect 9216 22332 9280 22336
rect 9216 22276 9220 22332
rect 9220 22276 9276 22332
rect 9276 22276 9280 22332
rect 9216 22272 9280 22276
rect 9296 22332 9360 22336
rect 9296 22276 9300 22332
rect 9300 22276 9356 22332
rect 9356 22276 9360 22332
rect 9296 22272 9360 22276
rect 9376 22332 9440 22336
rect 9376 22276 9380 22332
rect 9380 22276 9436 22332
rect 9436 22276 9440 22332
rect 9376 22272 9440 22276
rect 9456 22332 9520 22336
rect 9456 22276 9460 22332
rect 9460 22276 9516 22332
rect 9516 22276 9520 22332
rect 9456 22272 9520 22276
rect 19216 22332 19280 22336
rect 19216 22276 19220 22332
rect 19220 22276 19276 22332
rect 19276 22276 19280 22332
rect 19216 22272 19280 22276
rect 19296 22332 19360 22336
rect 19296 22276 19300 22332
rect 19300 22276 19356 22332
rect 19356 22276 19360 22332
rect 19296 22272 19360 22276
rect 19376 22332 19440 22336
rect 19376 22276 19380 22332
rect 19380 22276 19436 22332
rect 19436 22276 19440 22332
rect 19376 22272 19440 22276
rect 19456 22332 19520 22336
rect 19456 22276 19460 22332
rect 19460 22276 19516 22332
rect 19516 22276 19520 22332
rect 19456 22272 19520 22276
rect 29216 22332 29280 22336
rect 29216 22276 29220 22332
rect 29220 22276 29276 22332
rect 29276 22276 29280 22332
rect 29216 22272 29280 22276
rect 29296 22332 29360 22336
rect 29296 22276 29300 22332
rect 29300 22276 29356 22332
rect 29356 22276 29360 22332
rect 29296 22272 29360 22276
rect 29376 22332 29440 22336
rect 29376 22276 29380 22332
rect 29380 22276 29436 22332
rect 29436 22276 29440 22332
rect 29376 22272 29440 22276
rect 29456 22332 29520 22336
rect 29456 22276 29460 22332
rect 29460 22276 29516 22332
rect 29516 22276 29520 22332
rect 29456 22272 29520 22276
rect 39216 22332 39280 22336
rect 39216 22276 39220 22332
rect 39220 22276 39276 22332
rect 39276 22276 39280 22332
rect 39216 22272 39280 22276
rect 39296 22332 39360 22336
rect 39296 22276 39300 22332
rect 39300 22276 39356 22332
rect 39356 22276 39360 22332
rect 39296 22272 39360 22276
rect 39376 22332 39440 22336
rect 39376 22276 39380 22332
rect 39380 22276 39436 22332
rect 39436 22276 39440 22332
rect 39376 22272 39440 22276
rect 39456 22332 39520 22336
rect 39456 22276 39460 22332
rect 39460 22276 39516 22332
rect 39516 22276 39520 22332
rect 39456 22272 39520 22276
rect 49216 22332 49280 22336
rect 49216 22276 49220 22332
rect 49220 22276 49276 22332
rect 49276 22276 49280 22332
rect 49216 22272 49280 22276
rect 49296 22332 49360 22336
rect 49296 22276 49300 22332
rect 49300 22276 49356 22332
rect 49356 22276 49360 22332
rect 49296 22272 49360 22276
rect 49376 22332 49440 22336
rect 49376 22276 49380 22332
rect 49380 22276 49436 22332
rect 49436 22276 49440 22332
rect 49376 22272 49440 22276
rect 49456 22332 49520 22336
rect 49456 22276 49460 22332
rect 49460 22276 49516 22332
rect 49516 22276 49520 22332
rect 49456 22272 49520 22276
rect 59216 22332 59280 22336
rect 59216 22276 59220 22332
rect 59220 22276 59276 22332
rect 59276 22276 59280 22332
rect 59216 22272 59280 22276
rect 59296 22332 59360 22336
rect 59296 22276 59300 22332
rect 59300 22276 59356 22332
rect 59356 22276 59360 22332
rect 59296 22272 59360 22276
rect 59376 22332 59440 22336
rect 59376 22276 59380 22332
rect 59380 22276 59436 22332
rect 59436 22276 59440 22332
rect 59376 22272 59440 22276
rect 59456 22332 59520 22336
rect 59456 22276 59460 22332
rect 59460 22276 59516 22332
rect 59516 22276 59520 22332
rect 59456 22272 59520 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 14216 21788 14280 21792
rect 14216 21732 14220 21788
rect 14220 21732 14276 21788
rect 14276 21732 14280 21788
rect 14216 21728 14280 21732
rect 14296 21788 14360 21792
rect 14296 21732 14300 21788
rect 14300 21732 14356 21788
rect 14356 21732 14360 21788
rect 14296 21728 14360 21732
rect 14376 21788 14440 21792
rect 14376 21732 14380 21788
rect 14380 21732 14436 21788
rect 14436 21732 14440 21788
rect 14376 21728 14440 21732
rect 14456 21788 14520 21792
rect 14456 21732 14460 21788
rect 14460 21732 14516 21788
rect 14516 21732 14520 21788
rect 14456 21728 14520 21732
rect 24216 21788 24280 21792
rect 24216 21732 24220 21788
rect 24220 21732 24276 21788
rect 24276 21732 24280 21788
rect 24216 21728 24280 21732
rect 24296 21788 24360 21792
rect 24296 21732 24300 21788
rect 24300 21732 24356 21788
rect 24356 21732 24360 21788
rect 24296 21728 24360 21732
rect 24376 21788 24440 21792
rect 24376 21732 24380 21788
rect 24380 21732 24436 21788
rect 24436 21732 24440 21788
rect 24376 21728 24440 21732
rect 24456 21788 24520 21792
rect 24456 21732 24460 21788
rect 24460 21732 24516 21788
rect 24516 21732 24520 21788
rect 24456 21728 24520 21732
rect 34216 21788 34280 21792
rect 34216 21732 34220 21788
rect 34220 21732 34276 21788
rect 34276 21732 34280 21788
rect 34216 21728 34280 21732
rect 34296 21788 34360 21792
rect 34296 21732 34300 21788
rect 34300 21732 34356 21788
rect 34356 21732 34360 21788
rect 34296 21728 34360 21732
rect 34376 21788 34440 21792
rect 34376 21732 34380 21788
rect 34380 21732 34436 21788
rect 34436 21732 34440 21788
rect 34376 21728 34440 21732
rect 34456 21788 34520 21792
rect 34456 21732 34460 21788
rect 34460 21732 34516 21788
rect 34516 21732 34520 21788
rect 34456 21728 34520 21732
rect 44216 21788 44280 21792
rect 44216 21732 44220 21788
rect 44220 21732 44276 21788
rect 44276 21732 44280 21788
rect 44216 21728 44280 21732
rect 44296 21788 44360 21792
rect 44296 21732 44300 21788
rect 44300 21732 44356 21788
rect 44356 21732 44360 21788
rect 44296 21728 44360 21732
rect 44376 21788 44440 21792
rect 44376 21732 44380 21788
rect 44380 21732 44436 21788
rect 44436 21732 44440 21788
rect 44376 21728 44440 21732
rect 44456 21788 44520 21792
rect 44456 21732 44460 21788
rect 44460 21732 44516 21788
rect 44516 21732 44520 21788
rect 44456 21728 44520 21732
rect 54216 21788 54280 21792
rect 54216 21732 54220 21788
rect 54220 21732 54276 21788
rect 54276 21732 54280 21788
rect 54216 21728 54280 21732
rect 54296 21788 54360 21792
rect 54296 21732 54300 21788
rect 54300 21732 54356 21788
rect 54356 21732 54360 21788
rect 54296 21728 54360 21732
rect 54376 21788 54440 21792
rect 54376 21732 54380 21788
rect 54380 21732 54436 21788
rect 54436 21732 54440 21788
rect 54376 21728 54440 21732
rect 54456 21788 54520 21792
rect 54456 21732 54460 21788
rect 54460 21732 54516 21788
rect 54516 21732 54520 21788
rect 54456 21728 54520 21732
rect 64216 21788 64280 21792
rect 64216 21732 64220 21788
rect 64220 21732 64276 21788
rect 64276 21732 64280 21788
rect 64216 21728 64280 21732
rect 64296 21788 64360 21792
rect 64296 21732 64300 21788
rect 64300 21732 64356 21788
rect 64356 21732 64360 21788
rect 64296 21728 64360 21732
rect 64376 21788 64440 21792
rect 64376 21732 64380 21788
rect 64380 21732 64436 21788
rect 64436 21732 64440 21788
rect 64376 21728 64440 21732
rect 64456 21788 64520 21792
rect 64456 21732 64460 21788
rect 64460 21732 64516 21788
rect 64516 21732 64520 21788
rect 64456 21728 64520 21732
rect 39068 21388 39132 21452
rect 9216 21244 9280 21248
rect 9216 21188 9220 21244
rect 9220 21188 9276 21244
rect 9276 21188 9280 21244
rect 9216 21184 9280 21188
rect 9296 21244 9360 21248
rect 9296 21188 9300 21244
rect 9300 21188 9356 21244
rect 9356 21188 9360 21244
rect 9296 21184 9360 21188
rect 9376 21244 9440 21248
rect 9376 21188 9380 21244
rect 9380 21188 9436 21244
rect 9436 21188 9440 21244
rect 9376 21184 9440 21188
rect 9456 21244 9520 21248
rect 9456 21188 9460 21244
rect 9460 21188 9516 21244
rect 9516 21188 9520 21244
rect 9456 21184 9520 21188
rect 19216 21244 19280 21248
rect 19216 21188 19220 21244
rect 19220 21188 19276 21244
rect 19276 21188 19280 21244
rect 19216 21184 19280 21188
rect 19296 21244 19360 21248
rect 19296 21188 19300 21244
rect 19300 21188 19356 21244
rect 19356 21188 19360 21244
rect 19296 21184 19360 21188
rect 19376 21244 19440 21248
rect 19376 21188 19380 21244
rect 19380 21188 19436 21244
rect 19436 21188 19440 21244
rect 19376 21184 19440 21188
rect 19456 21244 19520 21248
rect 19456 21188 19460 21244
rect 19460 21188 19516 21244
rect 19516 21188 19520 21244
rect 19456 21184 19520 21188
rect 29216 21244 29280 21248
rect 29216 21188 29220 21244
rect 29220 21188 29276 21244
rect 29276 21188 29280 21244
rect 29216 21184 29280 21188
rect 29296 21244 29360 21248
rect 29296 21188 29300 21244
rect 29300 21188 29356 21244
rect 29356 21188 29360 21244
rect 29296 21184 29360 21188
rect 29376 21244 29440 21248
rect 29376 21188 29380 21244
rect 29380 21188 29436 21244
rect 29436 21188 29440 21244
rect 29376 21184 29440 21188
rect 29456 21244 29520 21248
rect 29456 21188 29460 21244
rect 29460 21188 29516 21244
rect 29516 21188 29520 21244
rect 29456 21184 29520 21188
rect 39216 21244 39280 21248
rect 39216 21188 39220 21244
rect 39220 21188 39276 21244
rect 39276 21188 39280 21244
rect 39216 21184 39280 21188
rect 39296 21244 39360 21248
rect 39296 21188 39300 21244
rect 39300 21188 39356 21244
rect 39356 21188 39360 21244
rect 39296 21184 39360 21188
rect 39376 21244 39440 21248
rect 39376 21188 39380 21244
rect 39380 21188 39436 21244
rect 39436 21188 39440 21244
rect 39376 21184 39440 21188
rect 39456 21244 39520 21248
rect 39456 21188 39460 21244
rect 39460 21188 39516 21244
rect 39516 21188 39520 21244
rect 39456 21184 39520 21188
rect 49216 21244 49280 21248
rect 49216 21188 49220 21244
rect 49220 21188 49276 21244
rect 49276 21188 49280 21244
rect 49216 21184 49280 21188
rect 49296 21244 49360 21248
rect 49296 21188 49300 21244
rect 49300 21188 49356 21244
rect 49356 21188 49360 21244
rect 49296 21184 49360 21188
rect 49376 21244 49440 21248
rect 49376 21188 49380 21244
rect 49380 21188 49436 21244
rect 49436 21188 49440 21244
rect 49376 21184 49440 21188
rect 49456 21244 49520 21248
rect 49456 21188 49460 21244
rect 49460 21188 49516 21244
rect 49516 21188 49520 21244
rect 49456 21184 49520 21188
rect 59216 21244 59280 21248
rect 59216 21188 59220 21244
rect 59220 21188 59276 21244
rect 59276 21188 59280 21244
rect 59216 21184 59280 21188
rect 59296 21244 59360 21248
rect 59296 21188 59300 21244
rect 59300 21188 59356 21244
rect 59356 21188 59360 21244
rect 59296 21184 59360 21188
rect 59376 21244 59440 21248
rect 59376 21188 59380 21244
rect 59380 21188 59436 21244
rect 59436 21188 59440 21244
rect 59376 21184 59440 21188
rect 59456 21244 59520 21248
rect 59456 21188 59460 21244
rect 59460 21188 59516 21244
rect 59516 21188 59520 21244
rect 59456 21184 59520 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 14216 20700 14280 20704
rect 14216 20644 14220 20700
rect 14220 20644 14276 20700
rect 14276 20644 14280 20700
rect 14216 20640 14280 20644
rect 14296 20700 14360 20704
rect 14296 20644 14300 20700
rect 14300 20644 14356 20700
rect 14356 20644 14360 20700
rect 14296 20640 14360 20644
rect 14376 20700 14440 20704
rect 14376 20644 14380 20700
rect 14380 20644 14436 20700
rect 14436 20644 14440 20700
rect 14376 20640 14440 20644
rect 14456 20700 14520 20704
rect 14456 20644 14460 20700
rect 14460 20644 14516 20700
rect 14516 20644 14520 20700
rect 14456 20640 14520 20644
rect 24216 20700 24280 20704
rect 24216 20644 24220 20700
rect 24220 20644 24276 20700
rect 24276 20644 24280 20700
rect 24216 20640 24280 20644
rect 24296 20700 24360 20704
rect 24296 20644 24300 20700
rect 24300 20644 24356 20700
rect 24356 20644 24360 20700
rect 24296 20640 24360 20644
rect 24376 20700 24440 20704
rect 24376 20644 24380 20700
rect 24380 20644 24436 20700
rect 24436 20644 24440 20700
rect 24376 20640 24440 20644
rect 24456 20700 24520 20704
rect 24456 20644 24460 20700
rect 24460 20644 24516 20700
rect 24516 20644 24520 20700
rect 24456 20640 24520 20644
rect 34216 20700 34280 20704
rect 34216 20644 34220 20700
rect 34220 20644 34276 20700
rect 34276 20644 34280 20700
rect 34216 20640 34280 20644
rect 34296 20700 34360 20704
rect 34296 20644 34300 20700
rect 34300 20644 34356 20700
rect 34356 20644 34360 20700
rect 34296 20640 34360 20644
rect 34376 20700 34440 20704
rect 34376 20644 34380 20700
rect 34380 20644 34436 20700
rect 34436 20644 34440 20700
rect 34376 20640 34440 20644
rect 34456 20700 34520 20704
rect 34456 20644 34460 20700
rect 34460 20644 34516 20700
rect 34516 20644 34520 20700
rect 34456 20640 34520 20644
rect 44216 20700 44280 20704
rect 44216 20644 44220 20700
rect 44220 20644 44276 20700
rect 44276 20644 44280 20700
rect 44216 20640 44280 20644
rect 44296 20700 44360 20704
rect 44296 20644 44300 20700
rect 44300 20644 44356 20700
rect 44356 20644 44360 20700
rect 44296 20640 44360 20644
rect 44376 20700 44440 20704
rect 44376 20644 44380 20700
rect 44380 20644 44436 20700
rect 44436 20644 44440 20700
rect 44376 20640 44440 20644
rect 44456 20700 44520 20704
rect 44456 20644 44460 20700
rect 44460 20644 44516 20700
rect 44516 20644 44520 20700
rect 44456 20640 44520 20644
rect 54216 20700 54280 20704
rect 54216 20644 54220 20700
rect 54220 20644 54276 20700
rect 54276 20644 54280 20700
rect 54216 20640 54280 20644
rect 54296 20700 54360 20704
rect 54296 20644 54300 20700
rect 54300 20644 54356 20700
rect 54356 20644 54360 20700
rect 54296 20640 54360 20644
rect 54376 20700 54440 20704
rect 54376 20644 54380 20700
rect 54380 20644 54436 20700
rect 54436 20644 54440 20700
rect 54376 20640 54440 20644
rect 54456 20700 54520 20704
rect 54456 20644 54460 20700
rect 54460 20644 54516 20700
rect 54516 20644 54520 20700
rect 54456 20640 54520 20644
rect 64216 20700 64280 20704
rect 64216 20644 64220 20700
rect 64220 20644 64276 20700
rect 64276 20644 64280 20700
rect 64216 20640 64280 20644
rect 64296 20700 64360 20704
rect 64296 20644 64300 20700
rect 64300 20644 64356 20700
rect 64356 20644 64360 20700
rect 64296 20640 64360 20644
rect 64376 20700 64440 20704
rect 64376 20644 64380 20700
rect 64380 20644 64436 20700
rect 64436 20644 64440 20700
rect 64376 20640 64440 20644
rect 64456 20700 64520 20704
rect 64456 20644 64460 20700
rect 64460 20644 64516 20700
rect 64516 20644 64520 20700
rect 64456 20640 64520 20644
rect 9216 20156 9280 20160
rect 9216 20100 9220 20156
rect 9220 20100 9276 20156
rect 9276 20100 9280 20156
rect 9216 20096 9280 20100
rect 9296 20156 9360 20160
rect 9296 20100 9300 20156
rect 9300 20100 9356 20156
rect 9356 20100 9360 20156
rect 9296 20096 9360 20100
rect 9376 20156 9440 20160
rect 9376 20100 9380 20156
rect 9380 20100 9436 20156
rect 9436 20100 9440 20156
rect 9376 20096 9440 20100
rect 9456 20156 9520 20160
rect 9456 20100 9460 20156
rect 9460 20100 9516 20156
rect 9516 20100 9520 20156
rect 9456 20096 9520 20100
rect 19216 20156 19280 20160
rect 19216 20100 19220 20156
rect 19220 20100 19276 20156
rect 19276 20100 19280 20156
rect 19216 20096 19280 20100
rect 19296 20156 19360 20160
rect 19296 20100 19300 20156
rect 19300 20100 19356 20156
rect 19356 20100 19360 20156
rect 19296 20096 19360 20100
rect 19376 20156 19440 20160
rect 19376 20100 19380 20156
rect 19380 20100 19436 20156
rect 19436 20100 19440 20156
rect 19376 20096 19440 20100
rect 19456 20156 19520 20160
rect 19456 20100 19460 20156
rect 19460 20100 19516 20156
rect 19516 20100 19520 20156
rect 19456 20096 19520 20100
rect 29216 20156 29280 20160
rect 29216 20100 29220 20156
rect 29220 20100 29276 20156
rect 29276 20100 29280 20156
rect 29216 20096 29280 20100
rect 29296 20156 29360 20160
rect 29296 20100 29300 20156
rect 29300 20100 29356 20156
rect 29356 20100 29360 20156
rect 29296 20096 29360 20100
rect 29376 20156 29440 20160
rect 29376 20100 29380 20156
rect 29380 20100 29436 20156
rect 29436 20100 29440 20156
rect 29376 20096 29440 20100
rect 29456 20156 29520 20160
rect 29456 20100 29460 20156
rect 29460 20100 29516 20156
rect 29516 20100 29520 20156
rect 29456 20096 29520 20100
rect 39216 20156 39280 20160
rect 39216 20100 39220 20156
rect 39220 20100 39276 20156
rect 39276 20100 39280 20156
rect 39216 20096 39280 20100
rect 39296 20156 39360 20160
rect 39296 20100 39300 20156
rect 39300 20100 39356 20156
rect 39356 20100 39360 20156
rect 39296 20096 39360 20100
rect 39376 20156 39440 20160
rect 39376 20100 39380 20156
rect 39380 20100 39436 20156
rect 39436 20100 39440 20156
rect 39376 20096 39440 20100
rect 39456 20156 39520 20160
rect 39456 20100 39460 20156
rect 39460 20100 39516 20156
rect 39516 20100 39520 20156
rect 39456 20096 39520 20100
rect 49216 20156 49280 20160
rect 49216 20100 49220 20156
rect 49220 20100 49276 20156
rect 49276 20100 49280 20156
rect 49216 20096 49280 20100
rect 49296 20156 49360 20160
rect 49296 20100 49300 20156
rect 49300 20100 49356 20156
rect 49356 20100 49360 20156
rect 49296 20096 49360 20100
rect 49376 20156 49440 20160
rect 49376 20100 49380 20156
rect 49380 20100 49436 20156
rect 49436 20100 49440 20156
rect 49376 20096 49440 20100
rect 49456 20156 49520 20160
rect 49456 20100 49460 20156
rect 49460 20100 49516 20156
rect 49516 20100 49520 20156
rect 49456 20096 49520 20100
rect 59216 20156 59280 20160
rect 59216 20100 59220 20156
rect 59220 20100 59276 20156
rect 59276 20100 59280 20156
rect 59216 20096 59280 20100
rect 59296 20156 59360 20160
rect 59296 20100 59300 20156
rect 59300 20100 59356 20156
rect 59356 20100 59360 20156
rect 59296 20096 59360 20100
rect 59376 20156 59440 20160
rect 59376 20100 59380 20156
rect 59380 20100 59436 20156
rect 59436 20100 59440 20156
rect 59376 20096 59440 20100
rect 59456 20156 59520 20160
rect 59456 20100 59460 20156
rect 59460 20100 59516 20156
rect 59516 20100 59520 20156
rect 59456 20096 59520 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 14216 19612 14280 19616
rect 14216 19556 14220 19612
rect 14220 19556 14276 19612
rect 14276 19556 14280 19612
rect 14216 19552 14280 19556
rect 14296 19612 14360 19616
rect 14296 19556 14300 19612
rect 14300 19556 14356 19612
rect 14356 19556 14360 19612
rect 14296 19552 14360 19556
rect 14376 19612 14440 19616
rect 14376 19556 14380 19612
rect 14380 19556 14436 19612
rect 14436 19556 14440 19612
rect 14376 19552 14440 19556
rect 14456 19612 14520 19616
rect 14456 19556 14460 19612
rect 14460 19556 14516 19612
rect 14516 19556 14520 19612
rect 14456 19552 14520 19556
rect 24216 19612 24280 19616
rect 24216 19556 24220 19612
rect 24220 19556 24276 19612
rect 24276 19556 24280 19612
rect 24216 19552 24280 19556
rect 24296 19612 24360 19616
rect 24296 19556 24300 19612
rect 24300 19556 24356 19612
rect 24356 19556 24360 19612
rect 24296 19552 24360 19556
rect 24376 19612 24440 19616
rect 24376 19556 24380 19612
rect 24380 19556 24436 19612
rect 24436 19556 24440 19612
rect 24376 19552 24440 19556
rect 24456 19612 24520 19616
rect 24456 19556 24460 19612
rect 24460 19556 24516 19612
rect 24516 19556 24520 19612
rect 24456 19552 24520 19556
rect 34216 19612 34280 19616
rect 34216 19556 34220 19612
rect 34220 19556 34276 19612
rect 34276 19556 34280 19612
rect 34216 19552 34280 19556
rect 34296 19612 34360 19616
rect 34296 19556 34300 19612
rect 34300 19556 34356 19612
rect 34356 19556 34360 19612
rect 34296 19552 34360 19556
rect 34376 19612 34440 19616
rect 34376 19556 34380 19612
rect 34380 19556 34436 19612
rect 34436 19556 34440 19612
rect 34376 19552 34440 19556
rect 34456 19612 34520 19616
rect 34456 19556 34460 19612
rect 34460 19556 34516 19612
rect 34516 19556 34520 19612
rect 34456 19552 34520 19556
rect 44216 19612 44280 19616
rect 44216 19556 44220 19612
rect 44220 19556 44276 19612
rect 44276 19556 44280 19612
rect 44216 19552 44280 19556
rect 44296 19612 44360 19616
rect 44296 19556 44300 19612
rect 44300 19556 44356 19612
rect 44356 19556 44360 19612
rect 44296 19552 44360 19556
rect 44376 19612 44440 19616
rect 44376 19556 44380 19612
rect 44380 19556 44436 19612
rect 44436 19556 44440 19612
rect 44376 19552 44440 19556
rect 44456 19612 44520 19616
rect 44456 19556 44460 19612
rect 44460 19556 44516 19612
rect 44516 19556 44520 19612
rect 44456 19552 44520 19556
rect 54216 19612 54280 19616
rect 54216 19556 54220 19612
rect 54220 19556 54276 19612
rect 54276 19556 54280 19612
rect 54216 19552 54280 19556
rect 54296 19612 54360 19616
rect 54296 19556 54300 19612
rect 54300 19556 54356 19612
rect 54356 19556 54360 19612
rect 54296 19552 54360 19556
rect 54376 19612 54440 19616
rect 54376 19556 54380 19612
rect 54380 19556 54436 19612
rect 54436 19556 54440 19612
rect 54376 19552 54440 19556
rect 54456 19612 54520 19616
rect 54456 19556 54460 19612
rect 54460 19556 54516 19612
rect 54516 19556 54520 19612
rect 54456 19552 54520 19556
rect 64216 19612 64280 19616
rect 64216 19556 64220 19612
rect 64220 19556 64276 19612
rect 64276 19556 64280 19612
rect 64216 19552 64280 19556
rect 64296 19612 64360 19616
rect 64296 19556 64300 19612
rect 64300 19556 64356 19612
rect 64356 19556 64360 19612
rect 64296 19552 64360 19556
rect 64376 19612 64440 19616
rect 64376 19556 64380 19612
rect 64380 19556 64436 19612
rect 64436 19556 64440 19612
rect 64376 19552 64440 19556
rect 64456 19612 64520 19616
rect 64456 19556 64460 19612
rect 64460 19556 64516 19612
rect 64516 19556 64520 19612
rect 64456 19552 64520 19556
rect 9216 19068 9280 19072
rect 9216 19012 9220 19068
rect 9220 19012 9276 19068
rect 9276 19012 9280 19068
rect 9216 19008 9280 19012
rect 9296 19068 9360 19072
rect 9296 19012 9300 19068
rect 9300 19012 9356 19068
rect 9356 19012 9360 19068
rect 9296 19008 9360 19012
rect 9376 19068 9440 19072
rect 9376 19012 9380 19068
rect 9380 19012 9436 19068
rect 9436 19012 9440 19068
rect 9376 19008 9440 19012
rect 9456 19068 9520 19072
rect 9456 19012 9460 19068
rect 9460 19012 9516 19068
rect 9516 19012 9520 19068
rect 9456 19008 9520 19012
rect 39216 19068 39280 19072
rect 39216 19012 39220 19068
rect 39220 19012 39276 19068
rect 39276 19012 39280 19068
rect 39216 19008 39280 19012
rect 39296 19068 39360 19072
rect 39296 19012 39300 19068
rect 39300 19012 39356 19068
rect 39356 19012 39360 19068
rect 39296 19008 39360 19012
rect 39376 19068 39440 19072
rect 39376 19012 39380 19068
rect 39380 19012 39436 19068
rect 39436 19012 39440 19068
rect 39376 19008 39440 19012
rect 39456 19068 39520 19072
rect 39456 19012 39460 19068
rect 39460 19012 39516 19068
rect 39516 19012 39520 19068
rect 39456 19008 39520 19012
rect 49216 19068 49280 19072
rect 49216 19012 49220 19068
rect 49220 19012 49276 19068
rect 49276 19012 49280 19068
rect 49216 19008 49280 19012
rect 49296 19068 49360 19072
rect 49296 19012 49300 19068
rect 49300 19012 49356 19068
rect 49356 19012 49360 19068
rect 49296 19008 49360 19012
rect 49376 19068 49440 19072
rect 49376 19012 49380 19068
rect 49380 19012 49436 19068
rect 49436 19012 49440 19068
rect 49376 19008 49440 19012
rect 49456 19068 49520 19072
rect 49456 19012 49460 19068
rect 49460 19012 49516 19068
rect 49516 19012 49520 19068
rect 49456 19008 49520 19012
rect 59216 19068 59280 19072
rect 59216 19012 59220 19068
rect 59220 19012 59276 19068
rect 59276 19012 59280 19068
rect 59216 19008 59280 19012
rect 59296 19068 59360 19072
rect 59296 19012 59300 19068
rect 59300 19012 59356 19068
rect 59356 19012 59360 19068
rect 59296 19008 59360 19012
rect 59376 19068 59440 19072
rect 59376 19012 59380 19068
rect 59380 19012 59436 19068
rect 59436 19012 59440 19068
rect 59376 19008 59440 19012
rect 59456 19068 59520 19072
rect 59456 19012 59460 19068
rect 59460 19012 59516 19068
rect 59516 19012 59520 19068
rect 59456 19008 59520 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 14216 18524 14280 18528
rect 14216 18468 14220 18524
rect 14220 18468 14276 18524
rect 14276 18468 14280 18524
rect 14216 18464 14280 18468
rect 14296 18524 14360 18528
rect 14296 18468 14300 18524
rect 14300 18468 14356 18524
rect 14356 18468 14360 18524
rect 14296 18464 14360 18468
rect 14376 18524 14440 18528
rect 14376 18468 14380 18524
rect 14380 18468 14436 18524
rect 14436 18468 14440 18524
rect 14376 18464 14440 18468
rect 14456 18524 14520 18528
rect 14456 18468 14460 18524
rect 14460 18468 14516 18524
rect 14516 18468 14520 18524
rect 14456 18464 14520 18468
rect 44216 18524 44280 18528
rect 44216 18468 44220 18524
rect 44220 18468 44276 18524
rect 44276 18468 44280 18524
rect 44216 18464 44280 18468
rect 44296 18524 44360 18528
rect 44296 18468 44300 18524
rect 44300 18468 44356 18524
rect 44356 18468 44360 18524
rect 44296 18464 44360 18468
rect 44376 18524 44440 18528
rect 44376 18468 44380 18524
rect 44380 18468 44436 18524
rect 44436 18468 44440 18524
rect 44376 18464 44440 18468
rect 44456 18524 44520 18528
rect 44456 18468 44460 18524
rect 44460 18468 44516 18524
rect 44516 18468 44520 18524
rect 44456 18464 44520 18468
rect 54216 18524 54280 18528
rect 54216 18468 54220 18524
rect 54220 18468 54276 18524
rect 54276 18468 54280 18524
rect 54216 18464 54280 18468
rect 54296 18524 54360 18528
rect 54296 18468 54300 18524
rect 54300 18468 54356 18524
rect 54356 18468 54360 18524
rect 54296 18464 54360 18468
rect 54376 18524 54440 18528
rect 54376 18468 54380 18524
rect 54380 18468 54436 18524
rect 54436 18468 54440 18524
rect 54376 18464 54440 18468
rect 54456 18524 54520 18528
rect 54456 18468 54460 18524
rect 54460 18468 54516 18524
rect 54516 18468 54520 18524
rect 54456 18464 54520 18468
rect 64216 18524 64280 18528
rect 64216 18468 64220 18524
rect 64220 18468 64276 18524
rect 64276 18468 64280 18524
rect 64216 18464 64280 18468
rect 64296 18524 64360 18528
rect 64296 18468 64300 18524
rect 64300 18468 64356 18524
rect 64356 18468 64360 18524
rect 64296 18464 64360 18468
rect 64376 18524 64440 18528
rect 64376 18468 64380 18524
rect 64380 18468 64436 18524
rect 64436 18468 64440 18524
rect 64376 18464 64440 18468
rect 64456 18524 64520 18528
rect 64456 18468 64460 18524
rect 64460 18468 64516 18524
rect 64516 18468 64520 18524
rect 64456 18464 64520 18468
rect 9216 17980 9280 17984
rect 9216 17924 9220 17980
rect 9220 17924 9276 17980
rect 9276 17924 9280 17980
rect 9216 17920 9280 17924
rect 9296 17980 9360 17984
rect 9296 17924 9300 17980
rect 9300 17924 9356 17980
rect 9356 17924 9360 17980
rect 9296 17920 9360 17924
rect 9376 17980 9440 17984
rect 9376 17924 9380 17980
rect 9380 17924 9436 17980
rect 9436 17924 9440 17980
rect 9376 17920 9440 17924
rect 9456 17980 9520 17984
rect 9456 17924 9460 17980
rect 9460 17924 9516 17980
rect 9516 17924 9520 17980
rect 9456 17920 9520 17924
rect 39216 17980 39280 17984
rect 39216 17924 39220 17980
rect 39220 17924 39276 17980
rect 39276 17924 39280 17980
rect 39216 17920 39280 17924
rect 39296 17980 39360 17984
rect 39296 17924 39300 17980
rect 39300 17924 39356 17980
rect 39356 17924 39360 17980
rect 39296 17920 39360 17924
rect 39376 17980 39440 17984
rect 39376 17924 39380 17980
rect 39380 17924 39436 17980
rect 39436 17924 39440 17980
rect 39376 17920 39440 17924
rect 39456 17980 39520 17984
rect 39456 17924 39460 17980
rect 39460 17924 39516 17980
rect 39516 17924 39520 17980
rect 39456 17920 39520 17924
rect 49216 17980 49280 17984
rect 49216 17924 49220 17980
rect 49220 17924 49276 17980
rect 49276 17924 49280 17980
rect 49216 17920 49280 17924
rect 49296 17980 49360 17984
rect 49296 17924 49300 17980
rect 49300 17924 49356 17980
rect 49356 17924 49360 17980
rect 49296 17920 49360 17924
rect 49376 17980 49440 17984
rect 49376 17924 49380 17980
rect 49380 17924 49436 17980
rect 49436 17924 49440 17980
rect 49376 17920 49440 17924
rect 49456 17980 49520 17984
rect 49456 17924 49460 17980
rect 49460 17924 49516 17980
rect 49516 17924 49520 17980
rect 49456 17920 49520 17924
rect 59216 17980 59280 17984
rect 59216 17924 59220 17980
rect 59220 17924 59276 17980
rect 59276 17924 59280 17980
rect 59216 17920 59280 17924
rect 59296 17980 59360 17984
rect 59296 17924 59300 17980
rect 59300 17924 59356 17980
rect 59356 17924 59360 17980
rect 59296 17920 59360 17924
rect 59376 17980 59440 17984
rect 59376 17924 59380 17980
rect 59380 17924 59436 17980
rect 59436 17924 59440 17980
rect 59376 17920 59440 17924
rect 59456 17980 59520 17984
rect 59456 17924 59460 17980
rect 59460 17924 59516 17980
rect 59516 17924 59520 17980
rect 59456 17920 59520 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 14216 17436 14280 17440
rect 14216 17380 14220 17436
rect 14220 17380 14276 17436
rect 14276 17380 14280 17436
rect 14216 17376 14280 17380
rect 14296 17436 14360 17440
rect 14296 17380 14300 17436
rect 14300 17380 14356 17436
rect 14356 17380 14360 17436
rect 14296 17376 14360 17380
rect 14376 17436 14440 17440
rect 14376 17380 14380 17436
rect 14380 17380 14436 17436
rect 14436 17380 14440 17436
rect 14376 17376 14440 17380
rect 14456 17436 14520 17440
rect 14456 17380 14460 17436
rect 14460 17380 14516 17436
rect 14516 17380 14520 17436
rect 14456 17376 14520 17380
rect 44216 17436 44280 17440
rect 44216 17380 44220 17436
rect 44220 17380 44276 17436
rect 44276 17380 44280 17436
rect 44216 17376 44280 17380
rect 44296 17436 44360 17440
rect 44296 17380 44300 17436
rect 44300 17380 44356 17436
rect 44356 17380 44360 17436
rect 44296 17376 44360 17380
rect 44376 17436 44440 17440
rect 44376 17380 44380 17436
rect 44380 17380 44436 17436
rect 44436 17380 44440 17436
rect 44376 17376 44440 17380
rect 44456 17436 44520 17440
rect 44456 17380 44460 17436
rect 44460 17380 44516 17436
rect 44516 17380 44520 17436
rect 44456 17376 44520 17380
rect 54216 17436 54280 17440
rect 54216 17380 54220 17436
rect 54220 17380 54276 17436
rect 54276 17380 54280 17436
rect 54216 17376 54280 17380
rect 54296 17436 54360 17440
rect 54296 17380 54300 17436
rect 54300 17380 54356 17436
rect 54356 17380 54360 17436
rect 54296 17376 54360 17380
rect 54376 17436 54440 17440
rect 54376 17380 54380 17436
rect 54380 17380 54436 17436
rect 54436 17380 54440 17436
rect 54376 17376 54440 17380
rect 54456 17436 54520 17440
rect 54456 17380 54460 17436
rect 54460 17380 54516 17436
rect 54516 17380 54520 17436
rect 54456 17376 54520 17380
rect 64216 17436 64280 17440
rect 64216 17380 64220 17436
rect 64220 17380 64276 17436
rect 64276 17380 64280 17436
rect 64216 17376 64280 17380
rect 64296 17436 64360 17440
rect 64296 17380 64300 17436
rect 64300 17380 64356 17436
rect 64356 17380 64360 17436
rect 64296 17376 64360 17380
rect 64376 17436 64440 17440
rect 64376 17380 64380 17436
rect 64380 17380 64436 17436
rect 64436 17380 64440 17436
rect 64376 17376 64440 17380
rect 64456 17436 64520 17440
rect 64456 17380 64460 17436
rect 64460 17380 64516 17436
rect 64516 17380 64520 17436
rect 64456 17376 64520 17380
rect 39804 17172 39868 17236
rect 9216 16892 9280 16896
rect 9216 16836 9220 16892
rect 9220 16836 9276 16892
rect 9276 16836 9280 16892
rect 9216 16832 9280 16836
rect 9296 16892 9360 16896
rect 9296 16836 9300 16892
rect 9300 16836 9356 16892
rect 9356 16836 9360 16892
rect 9296 16832 9360 16836
rect 9376 16892 9440 16896
rect 9376 16836 9380 16892
rect 9380 16836 9436 16892
rect 9436 16836 9440 16892
rect 9376 16832 9440 16836
rect 9456 16892 9520 16896
rect 9456 16836 9460 16892
rect 9460 16836 9516 16892
rect 9516 16836 9520 16892
rect 9456 16832 9520 16836
rect 39216 16892 39280 16896
rect 39216 16836 39220 16892
rect 39220 16836 39276 16892
rect 39276 16836 39280 16892
rect 39216 16832 39280 16836
rect 39296 16892 39360 16896
rect 39296 16836 39300 16892
rect 39300 16836 39356 16892
rect 39356 16836 39360 16892
rect 39296 16832 39360 16836
rect 39376 16892 39440 16896
rect 39376 16836 39380 16892
rect 39380 16836 39436 16892
rect 39436 16836 39440 16892
rect 39376 16832 39440 16836
rect 39456 16892 39520 16896
rect 39456 16836 39460 16892
rect 39460 16836 39516 16892
rect 39516 16836 39520 16892
rect 39456 16832 39520 16836
rect 49216 16892 49280 16896
rect 49216 16836 49220 16892
rect 49220 16836 49276 16892
rect 49276 16836 49280 16892
rect 49216 16832 49280 16836
rect 49296 16892 49360 16896
rect 49296 16836 49300 16892
rect 49300 16836 49356 16892
rect 49356 16836 49360 16892
rect 49296 16832 49360 16836
rect 49376 16892 49440 16896
rect 49376 16836 49380 16892
rect 49380 16836 49436 16892
rect 49436 16836 49440 16892
rect 49376 16832 49440 16836
rect 49456 16892 49520 16896
rect 49456 16836 49460 16892
rect 49460 16836 49516 16892
rect 49516 16836 49520 16892
rect 49456 16832 49520 16836
rect 59216 16892 59280 16896
rect 59216 16836 59220 16892
rect 59220 16836 59276 16892
rect 59276 16836 59280 16892
rect 59216 16832 59280 16836
rect 59296 16892 59360 16896
rect 59296 16836 59300 16892
rect 59300 16836 59356 16892
rect 59356 16836 59360 16892
rect 59296 16832 59360 16836
rect 59376 16892 59440 16896
rect 59376 16836 59380 16892
rect 59380 16836 59436 16892
rect 59436 16836 59440 16892
rect 59376 16832 59440 16836
rect 59456 16892 59520 16896
rect 59456 16836 59460 16892
rect 59460 16836 59516 16892
rect 59516 16836 59520 16892
rect 59456 16832 59520 16836
rect 29216 16374 29280 16438
rect 29296 16374 29360 16438
rect 29376 16374 29440 16438
rect 29456 16374 29520 16438
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 14216 16348 14280 16352
rect 14216 16292 14220 16348
rect 14220 16292 14276 16348
rect 14276 16292 14280 16348
rect 14216 16288 14280 16292
rect 14296 16348 14360 16352
rect 14296 16292 14300 16348
rect 14300 16292 14356 16348
rect 14356 16292 14360 16348
rect 14296 16288 14360 16292
rect 14376 16348 14440 16352
rect 14376 16292 14380 16348
rect 14380 16292 14436 16348
rect 14436 16292 14440 16348
rect 14376 16288 14440 16292
rect 14456 16348 14520 16352
rect 14456 16292 14460 16348
rect 14460 16292 14516 16348
rect 14516 16292 14520 16348
rect 14456 16288 14520 16292
rect 29216 16294 29280 16358
rect 29296 16294 29360 16358
rect 29376 16294 29440 16358
rect 29456 16294 29520 16358
rect 44216 16348 44280 16352
rect 44216 16292 44220 16348
rect 44220 16292 44276 16348
rect 44276 16292 44280 16348
rect 44216 16288 44280 16292
rect 44296 16348 44360 16352
rect 44296 16292 44300 16348
rect 44300 16292 44356 16348
rect 44356 16292 44360 16348
rect 44296 16288 44360 16292
rect 44376 16348 44440 16352
rect 44376 16292 44380 16348
rect 44380 16292 44436 16348
rect 44436 16292 44440 16348
rect 44376 16288 44440 16292
rect 44456 16348 44520 16352
rect 44456 16292 44460 16348
rect 44460 16292 44516 16348
rect 44516 16292 44520 16348
rect 44456 16288 44520 16292
rect 54216 16348 54280 16352
rect 54216 16292 54220 16348
rect 54220 16292 54276 16348
rect 54276 16292 54280 16348
rect 54216 16288 54280 16292
rect 54296 16348 54360 16352
rect 54296 16292 54300 16348
rect 54300 16292 54356 16348
rect 54356 16292 54360 16348
rect 54296 16288 54360 16292
rect 54376 16348 54440 16352
rect 54376 16292 54380 16348
rect 54380 16292 54436 16348
rect 54436 16292 54440 16348
rect 54376 16288 54440 16292
rect 54456 16348 54520 16352
rect 54456 16292 54460 16348
rect 54460 16292 54516 16348
rect 54516 16292 54520 16348
rect 54456 16288 54520 16292
rect 64216 16348 64280 16352
rect 64216 16292 64220 16348
rect 64220 16292 64276 16348
rect 64276 16292 64280 16348
rect 64216 16288 64280 16292
rect 64296 16348 64360 16352
rect 64296 16292 64300 16348
rect 64300 16292 64356 16348
rect 64356 16292 64360 16348
rect 64296 16288 64360 16292
rect 64376 16348 64440 16352
rect 64376 16292 64380 16348
rect 64380 16292 64436 16348
rect 64436 16292 64440 16348
rect 64376 16288 64440 16292
rect 64456 16348 64520 16352
rect 64456 16292 64460 16348
rect 64460 16292 64516 16348
rect 64516 16292 64520 16348
rect 64456 16288 64520 16292
rect 29216 16214 29280 16278
rect 29296 16214 29360 16278
rect 29376 16214 29440 16278
rect 29456 16214 29520 16278
rect 29216 16134 29280 16198
rect 29296 16134 29360 16198
rect 29376 16134 29440 16198
rect 29456 16134 29520 16198
rect 29216 16054 29280 16118
rect 29296 16054 29360 16118
rect 29376 16054 29440 16118
rect 29456 16054 29520 16118
rect 9216 15804 9280 15808
rect 9216 15748 9220 15804
rect 9220 15748 9276 15804
rect 9276 15748 9280 15804
rect 9216 15744 9280 15748
rect 9296 15804 9360 15808
rect 9296 15748 9300 15804
rect 9300 15748 9356 15804
rect 9356 15748 9360 15804
rect 9296 15744 9360 15748
rect 9376 15804 9440 15808
rect 9376 15748 9380 15804
rect 9380 15748 9436 15804
rect 9436 15748 9440 15804
rect 9376 15744 9440 15748
rect 9456 15804 9520 15808
rect 9456 15748 9460 15804
rect 9460 15748 9516 15804
rect 9516 15748 9520 15804
rect 9456 15744 9520 15748
rect 39216 15804 39280 15808
rect 39216 15748 39220 15804
rect 39220 15748 39276 15804
rect 39276 15748 39280 15804
rect 39216 15744 39280 15748
rect 39296 15804 39360 15808
rect 39296 15748 39300 15804
rect 39300 15748 39356 15804
rect 39356 15748 39360 15804
rect 39296 15744 39360 15748
rect 39376 15804 39440 15808
rect 39376 15748 39380 15804
rect 39380 15748 39436 15804
rect 39436 15748 39440 15804
rect 39376 15744 39440 15748
rect 39456 15804 39520 15808
rect 39456 15748 39460 15804
rect 39460 15748 39516 15804
rect 39516 15748 39520 15804
rect 39456 15744 39520 15748
rect 49216 15804 49280 15808
rect 49216 15748 49220 15804
rect 49220 15748 49276 15804
rect 49276 15748 49280 15804
rect 49216 15744 49280 15748
rect 49296 15804 49360 15808
rect 49296 15748 49300 15804
rect 49300 15748 49356 15804
rect 49356 15748 49360 15804
rect 49296 15744 49360 15748
rect 49376 15804 49440 15808
rect 49376 15748 49380 15804
rect 49380 15748 49436 15804
rect 49436 15748 49440 15804
rect 49376 15744 49440 15748
rect 49456 15804 49520 15808
rect 49456 15748 49460 15804
rect 49460 15748 49516 15804
rect 49516 15748 49520 15804
rect 49456 15744 49520 15748
rect 59216 15804 59280 15808
rect 59216 15748 59220 15804
rect 59220 15748 59276 15804
rect 59276 15748 59280 15804
rect 59216 15744 59280 15748
rect 59296 15804 59360 15808
rect 59296 15748 59300 15804
rect 59300 15748 59356 15804
rect 59356 15748 59360 15804
rect 59296 15744 59360 15748
rect 59376 15804 59440 15808
rect 59376 15748 59380 15804
rect 59380 15748 59436 15804
rect 59436 15748 59440 15804
rect 59376 15744 59440 15748
rect 59456 15804 59520 15808
rect 59456 15748 59460 15804
rect 59460 15748 59516 15804
rect 59516 15748 59520 15804
rect 59456 15744 59520 15748
rect 24216 15574 24280 15638
rect 24296 15574 24360 15638
rect 24376 15574 24440 15638
rect 24456 15574 24520 15638
rect 24216 15494 24280 15558
rect 24296 15494 24360 15558
rect 24376 15494 24440 15558
rect 24456 15494 24520 15558
rect 24216 15414 24280 15478
rect 24296 15414 24360 15478
rect 24376 15414 24440 15478
rect 24456 15414 24520 15478
rect 24216 15334 24280 15398
rect 24296 15334 24360 15398
rect 24376 15334 24440 15398
rect 24456 15334 24520 15398
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 14216 15260 14280 15264
rect 14216 15204 14220 15260
rect 14220 15204 14276 15260
rect 14276 15204 14280 15260
rect 14216 15200 14280 15204
rect 14296 15260 14360 15264
rect 14296 15204 14300 15260
rect 14300 15204 14356 15260
rect 14356 15204 14360 15260
rect 14296 15200 14360 15204
rect 14376 15260 14440 15264
rect 14376 15204 14380 15260
rect 14380 15204 14436 15260
rect 14436 15204 14440 15260
rect 14376 15200 14440 15204
rect 14456 15260 14520 15264
rect 14456 15204 14460 15260
rect 14460 15204 14516 15260
rect 14516 15204 14520 15260
rect 14456 15200 14520 15204
rect 24216 15254 24280 15318
rect 24296 15254 24360 15318
rect 24376 15254 24440 15318
rect 24456 15254 24520 15318
rect 44216 15260 44280 15264
rect 44216 15204 44220 15260
rect 44220 15204 44276 15260
rect 44276 15204 44280 15260
rect 44216 15200 44280 15204
rect 44296 15260 44360 15264
rect 44296 15204 44300 15260
rect 44300 15204 44356 15260
rect 44356 15204 44360 15260
rect 44296 15200 44360 15204
rect 44376 15260 44440 15264
rect 44376 15204 44380 15260
rect 44380 15204 44436 15260
rect 44436 15204 44440 15260
rect 44376 15200 44440 15204
rect 44456 15260 44520 15264
rect 44456 15204 44460 15260
rect 44460 15204 44516 15260
rect 44516 15204 44520 15260
rect 44456 15200 44520 15204
rect 54216 15260 54280 15264
rect 54216 15204 54220 15260
rect 54220 15204 54276 15260
rect 54276 15204 54280 15260
rect 54216 15200 54280 15204
rect 54296 15260 54360 15264
rect 54296 15204 54300 15260
rect 54300 15204 54356 15260
rect 54356 15204 54360 15260
rect 54296 15200 54360 15204
rect 54376 15260 54440 15264
rect 54376 15204 54380 15260
rect 54380 15204 54436 15260
rect 54436 15204 54440 15260
rect 54376 15200 54440 15204
rect 54456 15260 54520 15264
rect 54456 15204 54460 15260
rect 54460 15204 54516 15260
rect 54516 15204 54520 15260
rect 54456 15200 54520 15204
rect 64216 15260 64280 15264
rect 64216 15204 64220 15260
rect 64220 15204 64276 15260
rect 64276 15204 64280 15260
rect 64216 15200 64280 15204
rect 64296 15260 64360 15264
rect 64296 15204 64300 15260
rect 64300 15204 64356 15260
rect 64356 15204 64360 15260
rect 64296 15200 64360 15204
rect 64376 15260 64440 15264
rect 64376 15204 64380 15260
rect 64380 15204 64436 15260
rect 64436 15204 64440 15260
rect 64376 15200 64440 15204
rect 64456 15260 64520 15264
rect 64456 15204 64460 15260
rect 64460 15204 64516 15260
rect 64516 15204 64520 15260
rect 64456 15200 64520 15204
rect 9216 14716 9280 14720
rect 9216 14660 9220 14716
rect 9220 14660 9276 14716
rect 9276 14660 9280 14716
rect 9216 14656 9280 14660
rect 9296 14716 9360 14720
rect 9296 14660 9300 14716
rect 9300 14660 9356 14716
rect 9356 14660 9360 14716
rect 9296 14656 9360 14660
rect 9376 14716 9440 14720
rect 9376 14660 9380 14716
rect 9380 14660 9436 14716
rect 9436 14660 9440 14716
rect 9376 14656 9440 14660
rect 9456 14716 9520 14720
rect 9456 14660 9460 14716
rect 9460 14660 9516 14716
rect 9516 14660 9520 14716
rect 9456 14656 9520 14660
rect 39216 14716 39280 14720
rect 39216 14660 39220 14716
rect 39220 14660 39276 14716
rect 39276 14660 39280 14716
rect 39216 14656 39280 14660
rect 39296 14716 39360 14720
rect 39296 14660 39300 14716
rect 39300 14660 39356 14716
rect 39356 14660 39360 14716
rect 39296 14656 39360 14660
rect 39376 14716 39440 14720
rect 39376 14660 39380 14716
rect 39380 14660 39436 14716
rect 39436 14660 39440 14716
rect 39376 14656 39440 14660
rect 39456 14716 39520 14720
rect 39456 14660 39460 14716
rect 39460 14660 39516 14716
rect 39516 14660 39520 14716
rect 39456 14656 39520 14660
rect 49216 14716 49280 14720
rect 49216 14660 49220 14716
rect 49220 14660 49276 14716
rect 49276 14660 49280 14716
rect 49216 14656 49280 14660
rect 49296 14716 49360 14720
rect 49296 14660 49300 14716
rect 49300 14660 49356 14716
rect 49356 14660 49360 14716
rect 49296 14656 49360 14660
rect 49376 14716 49440 14720
rect 49376 14660 49380 14716
rect 49380 14660 49436 14716
rect 49436 14660 49440 14716
rect 49376 14656 49440 14660
rect 49456 14716 49520 14720
rect 49456 14660 49460 14716
rect 49460 14660 49516 14716
rect 49516 14660 49520 14716
rect 49456 14656 49520 14660
rect 59216 14716 59280 14720
rect 59216 14660 59220 14716
rect 59220 14660 59276 14716
rect 59276 14660 59280 14716
rect 59216 14656 59280 14660
rect 59296 14716 59360 14720
rect 59296 14660 59300 14716
rect 59300 14660 59356 14716
rect 59356 14660 59360 14716
rect 59296 14656 59360 14660
rect 59376 14716 59440 14720
rect 59376 14660 59380 14716
rect 59380 14660 59436 14716
rect 59436 14660 59440 14716
rect 59376 14656 59440 14660
rect 59456 14716 59520 14720
rect 59456 14660 59460 14716
rect 59460 14660 59516 14716
rect 59516 14660 59520 14716
rect 59456 14656 59520 14660
rect 40172 14452 40236 14516
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 14216 14172 14280 14176
rect 14216 14116 14220 14172
rect 14220 14116 14276 14172
rect 14276 14116 14280 14172
rect 14216 14112 14280 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 44216 14172 44280 14176
rect 44216 14116 44220 14172
rect 44220 14116 44276 14172
rect 44276 14116 44280 14172
rect 44216 14112 44280 14116
rect 44296 14172 44360 14176
rect 44296 14116 44300 14172
rect 44300 14116 44356 14172
rect 44356 14116 44360 14172
rect 44296 14112 44360 14116
rect 44376 14172 44440 14176
rect 44376 14116 44380 14172
rect 44380 14116 44436 14172
rect 44436 14116 44440 14172
rect 44376 14112 44440 14116
rect 44456 14172 44520 14176
rect 44456 14116 44460 14172
rect 44460 14116 44516 14172
rect 44516 14116 44520 14172
rect 44456 14112 44520 14116
rect 54216 14172 54280 14176
rect 54216 14116 54220 14172
rect 54220 14116 54276 14172
rect 54276 14116 54280 14172
rect 54216 14112 54280 14116
rect 54296 14172 54360 14176
rect 54296 14116 54300 14172
rect 54300 14116 54356 14172
rect 54356 14116 54360 14172
rect 54296 14112 54360 14116
rect 54376 14172 54440 14176
rect 54376 14116 54380 14172
rect 54380 14116 54436 14172
rect 54436 14116 54440 14172
rect 54376 14112 54440 14116
rect 54456 14172 54520 14176
rect 54456 14116 54460 14172
rect 54460 14116 54516 14172
rect 54516 14116 54520 14172
rect 54456 14112 54520 14116
rect 64216 14172 64280 14176
rect 64216 14116 64220 14172
rect 64220 14116 64276 14172
rect 64276 14116 64280 14172
rect 64216 14112 64280 14116
rect 64296 14172 64360 14176
rect 64296 14116 64300 14172
rect 64300 14116 64356 14172
rect 64356 14116 64360 14172
rect 64296 14112 64360 14116
rect 64376 14172 64440 14176
rect 64376 14116 64380 14172
rect 64380 14116 64436 14172
rect 64436 14116 64440 14172
rect 64376 14112 64440 14116
rect 64456 14172 64520 14176
rect 64456 14116 64460 14172
rect 64460 14116 64516 14172
rect 64516 14116 64520 14172
rect 64456 14112 64520 14116
rect 15700 13772 15764 13836
rect 16252 13832 16316 13836
rect 16252 13776 16302 13832
rect 16302 13776 16316 13832
rect 16252 13772 16316 13776
rect 9216 13628 9280 13632
rect 9216 13572 9220 13628
rect 9220 13572 9276 13628
rect 9276 13572 9280 13628
rect 9216 13568 9280 13572
rect 9296 13628 9360 13632
rect 9296 13572 9300 13628
rect 9300 13572 9356 13628
rect 9356 13572 9360 13628
rect 9296 13568 9360 13572
rect 9376 13628 9440 13632
rect 9376 13572 9380 13628
rect 9380 13572 9436 13628
rect 9436 13572 9440 13628
rect 9376 13568 9440 13572
rect 9456 13628 9520 13632
rect 9456 13572 9460 13628
rect 9460 13572 9516 13628
rect 9516 13572 9520 13628
rect 9456 13568 9520 13572
rect 39216 13628 39280 13632
rect 39216 13572 39220 13628
rect 39220 13572 39276 13628
rect 39276 13572 39280 13628
rect 39216 13568 39280 13572
rect 39296 13628 39360 13632
rect 39296 13572 39300 13628
rect 39300 13572 39356 13628
rect 39356 13572 39360 13628
rect 39296 13568 39360 13572
rect 39376 13628 39440 13632
rect 39376 13572 39380 13628
rect 39380 13572 39436 13628
rect 39436 13572 39440 13628
rect 39376 13568 39440 13572
rect 39456 13628 39520 13632
rect 39456 13572 39460 13628
rect 39460 13572 39516 13628
rect 39516 13572 39520 13628
rect 39456 13568 39520 13572
rect 49216 13628 49280 13632
rect 49216 13572 49220 13628
rect 49220 13572 49276 13628
rect 49276 13572 49280 13628
rect 49216 13568 49280 13572
rect 49296 13628 49360 13632
rect 49296 13572 49300 13628
rect 49300 13572 49356 13628
rect 49356 13572 49360 13628
rect 49296 13568 49360 13572
rect 49376 13628 49440 13632
rect 49376 13572 49380 13628
rect 49380 13572 49436 13628
rect 49436 13572 49440 13628
rect 49376 13568 49440 13572
rect 49456 13628 49520 13632
rect 49456 13572 49460 13628
rect 49460 13572 49516 13628
rect 49516 13572 49520 13628
rect 49456 13568 49520 13572
rect 59216 13628 59280 13632
rect 59216 13572 59220 13628
rect 59220 13572 59276 13628
rect 59276 13572 59280 13628
rect 59216 13568 59280 13572
rect 59296 13628 59360 13632
rect 59296 13572 59300 13628
rect 59300 13572 59356 13628
rect 59356 13572 59360 13628
rect 59296 13568 59360 13572
rect 59376 13628 59440 13632
rect 59376 13572 59380 13628
rect 59380 13572 59436 13628
rect 59436 13572 59440 13628
rect 59376 13568 59440 13572
rect 59456 13628 59520 13632
rect 59456 13572 59460 13628
rect 59460 13572 59516 13628
rect 59516 13572 59520 13628
rect 59456 13568 59520 13572
rect 13492 13152 13556 13156
rect 13492 13096 13542 13152
rect 13542 13096 13556 13152
rect 13492 13092 13556 13096
rect 39068 13092 39132 13156
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 14216 13084 14280 13088
rect 14216 13028 14220 13084
rect 14220 13028 14276 13084
rect 14276 13028 14280 13084
rect 14216 13024 14280 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 44216 13084 44280 13088
rect 44216 13028 44220 13084
rect 44220 13028 44276 13084
rect 44276 13028 44280 13084
rect 44216 13024 44280 13028
rect 44296 13084 44360 13088
rect 44296 13028 44300 13084
rect 44300 13028 44356 13084
rect 44356 13028 44360 13084
rect 44296 13024 44360 13028
rect 44376 13084 44440 13088
rect 44376 13028 44380 13084
rect 44380 13028 44436 13084
rect 44436 13028 44440 13084
rect 44376 13024 44440 13028
rect 44456 13084 44520 13088
rect 44456 13028 44460 13084
rect 44460 13028 44516 13084
rect 44516 13028 44520 13084
rect 44456 13024 44520 13028
rect 54216 13084 54280 13088
rect 54216 13028 54220 13084
rect 54220 13028 54276 13084
rect 54276 13028 54280 13084
rect 54216 13024 54280 13028
rect 54296 13084 54360 13088
rect 54296 13028 54300 13084
rect 54300 13028 54356 13084
rect 54356 13028 54360 13084
rect 54296 13024 54360 13028
rect 54376 13084 54440 13088
rect 54376 13028 54380 13084
rect 54380 13028 54436 13084
rect 54436 13028 54440 13084
rect 54376 13024 54440 13028
rect 54456 13084 54520 13088
rect 54456 13028 54460 13084
rect 54460 13028 54516 13084
rect 54516 13028 54520 13084
rect 54456 13024 54520 13028
rect 64216 13084 64280 13088
rect 64216 13028 64220 13084
rect 64220 13028 64276 13084
rect 64276 13028 64280 13084
rect 64216 13024 64280 13028
rect 64296 13084 64360 13088
rect 64296 13028 64300 13084
rect 64300 13028 64356 13084
rect 64356 13028 64360 13084
rect 64296 13024 64360 13028
rect 64376 13084 64440 13088
rect 64376 13028 64380 13084
rect 64380 13028 64436 13084
rect 64436 13028 64440 13084
rect 64376 13024 64440 13028
rect 64456 13084 64520 13088
rect 64456 13028 64460 13084
rect 64460 13028 64516 13084
rect 64516 13028 64520 13084
rect 64456 13024 64520 13028
rect 39804 12956 39868 13020
rect 13124 12548 13188 12612
rect 40724 12548 40788 12612
rect 9216 12540 9280 12544
rect 9216 12484 9220 12540
rect 9220 12484 9276 12540
rect 9276 12484 9280 12540
rect 9216 12480 9280 12484
rect 9296 12540 9360 12544
rect 9296 12484 9300 12540
rect 9300 12484 9356 12540
rect 9356 12484 9360 12540
rect 9296 12480 9360 12484
rect 9376 12540 9440 12544
rect 9376 12484 9380 12540
rect 9380 12484 9436 12540
rect 9436 12484 9440 12540
rect 9376 12480 9440 12484
rect 9456 12540 9520 12544
rect 9456 12484 9460 12540
rect 9460 12484 9516 12540
rect 9516 12484 9520 12540
rect 9456 12480 9520 12484
rect 39216 12540 39280 12544
rect 39216 12484 39220 12540
rect 39220 12484 39276 12540
rect 39276 12484 39280 12540
rect 39216 12480 39280 12484
rect 39296 12540 39360 12544
rect 39296 12484 39300 12540
rect 39300 12484 39356 12540
rect 39356 12484 39360 12540
rect 39296 12480 39360 12484
rect 39376 12540 39440 12544
rect 39376 12484 39380 12540
rect 39380 12484 39436 12540
rect 39436 12484 39440 12540
rect 39376 12480 39440 12484
rect 39456 12540 39520 12544
rect 39456 12484 39460 12540
rect 39460 12484 39516 12540
rect 39516 12484 39520 12540
rect 39456 12480 39520 12484
rect 49216 12540 49280 12544
rect 49216 12484 49220 12540
rect 49220 12484 49276 12540
rect 49276 12484 49280 12540
rect 49216 12480 49280 12484
rect 49296 12540 49360 12544
rect 49296 12484 49300 12540
rect 49300 12484 49356 12540
rect 49356 12484 49360 12540
rect 49296 12480 49360 12484
rect 49376 12540 49440 12544
rect 49376 12484 49380 12540
rect 49380 12484 49436 12540
rect 49436 12484 49440 12540
rect 49376 12480 49440 12484
rect 49456 12540 49520 12544
rect 49456 12484 49460 12540
rect 49460 12484 49516 12540
rect 49516 12484 49520 12540
rect 49456 12480 49520 12484
rect 59216 12540 59280 12544
rect 59216 12484 59220 12540
rect 59220 12484 59276 12540
rect 59276 12484 59280 12540
rect 59216 12480 59280 12484
rect 59296 12540 59360 12544
rect 59296 12484 59300 12540
rect 59300 12484 59356 12540
rect 59356 12484 59360 12540
rect 59296 12480 59360 12484
rect 59376 12540 59440 12544
rect 59376 12484 59380 12540
rect 59380 12484 59436 12540
rect 59436 12484 59440 12540
rect 59376 12480 59440 12484
rect 59456 12540 59520 12544
rect 59456 12484 59460 12540
rect 59460 12484 59516 12540
rect 59516 12484 59520 12540
rect 59456 12480 59520 12484
rect 39620 12412 39684 12476
rect 38700 12140 38764 12204
rect 39804 12200 39868 12204
rect 39804 12144 39818 12200
rect 39818 12144 39868 12200
rect 39804 12140 39868 12144
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 14216 11996 14280 12000
rect 14216 11940 14220 11996
rect 14220 11940 14276 11996
rect 14276 11940 14280 11996
rect 14216 11936 14280 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 44216 11996 44280 12000
rect 44216 11940 44220 11996
rect 44220 11940 44276 11996
rect 44276 11940 44280 11996
rect 44216 11936 44280 11940
rect 44296 11996 44360 12000
rect 44296 11940 44300 11996
rect 44300 11940 44356 11996
rect 44356 11940 44360 11996
rect 44296 11936 44360 11940
rect 44376 11996 44440 12000
rect 44376 11940 44380 11996
rect 44380 11940 44436 11996
rect 44436 11940 44440 11996
rect 44376 11936 44440 11940
rect 44456 11996 44520 12000
rect 44456 11940 44460 11996
rect 44460 11940 44516 11996
rect 44516 11940 44520 11996
rect 44456 11936 44520 11940
rect 54216 11996 54280 12000
rect 54216 11940 54220 11996
rect 54220 11940 54276 11996
rect 54276 11940 54280 11996
rect 54216 11936 54280 11940
rect 54296 11996 54360 12000
rect 54296 11940 54300 11996
rect 54300 11940 54356 11996
rect 54356 11940 54360 11996
rect 54296 11936 54360 11940
rect 54376 11996 54440 12000
rect 54376 11940 54380 11996
rect 54380 11940 54436 11996
rect 54436 11940 54440 11996
rect 54376 11936 54440 11940
rect 54456 11996 54520 12000
rect 54456 11940 54460 11996
rect 54460 11940 54516 11996
rect 54516 11940 54520 11996
rect 54456 11936 54520 11940
rect 64216 11996 64280 12000
rect 64216 11940 64220 11996
rect 64220 11940 64276 11996
rect 64276 11940 64280 11996
rect 64216 11936 64280 11940
rect 64296 11996 64360 12000
rect 64296 11940 64300 11996
rect 64300 11940 64356 11996
rect 64356 11940 64360 11996
rect 64296 11936 64360 11940
rect 64376 11996 64440 12000
rect 64376 11940 64380 11996
rect 64380 11940 64436 11996
rect 64436 11940 64440 11996
rect 64376 11936 64440 11940
rect 64456 11996 64520 12000
rect 64456 11940 64460 11996
rect 64460 11940 64516 11996
rect 64516 11940 64520 11996
rect 64456 11936 64520 11940
rect 24216 11843 24280 11907
rect 24296 11843 24360 11907
rect 24376 11843 24440 11907
rect 24456 11843 24520 11907
rect 24216 11763 24280 11827
rect 24296 11763 24360 11827
rect 24376 11763 24440 11827
rect 24456 11763 24520 11827
rect 24216 11683 24280 11747
rect 24296 11683 24360 11747
rect 24376 11683 24440 11747
rect 24456 11683 24520 11747
rect 14780 11656 14844 11660
rect 14780 11600 14830 11656
rect 14830 11600 14844 11656
rect 14780 11596 14844 11600
rect 24216 11603 24280 11667
rect 24296 11603 24360 11667
rect 24376 11603 24440 11667
rect 24456 11603 24520 11667
rect 34216 11843 34280 11907
rect 34296 11843 34360 11907
rect 34376 11843 34440 11907
rect 34456 11843 34520 11907
rect 34216 11763 34280 11827
rect 34296 11763 34360 11827
rect 34376 11763 34440 11827
rect 34456 11763 34520 11827
rect 34216 11683 34280 11747
rect 34296 11683 34360 11747
rect 34376 11683 34440 11747
rect 34456 11683 34520 11747
rect 34216 11603 34280 11667
rect 34296 11603 34360 11667
rect 34376 11603 34440 11667
rect 34456 11603 34520 11667
rect 9216 11452 9280 11456
rect 9216 11396 9220 11452
rect 9220 11396 9276 11452
rect 9276 11396 9280 11452
rect 9216 11392 9280 11396
rect 9296 11452 9360 11456
rect 9296 11396 9300 11452
rect 9300 11396 9356 11452
rect 9356 11396 9360 11452
rect 9296 11392 9360 11396
rect 9376 11452 9440 11456
rect 9376 11396 9380 11452
rect 9380 11396 9436 11452
rect 9436 11396 9440 11452
rect 9376 11392 9440 11396
rect 9456 11452 9520 11456
rect 9456 11396 9460 11452
rect 9460 11396 9516 11452
rect 9516 11396 9520 11452
rect 9456 11392 9520 11396
rect 39216 11452 39280 11456
rect 39216 11396 39220 11452
rect 39220 11396 39276 11452
rect 39276 11396 39280 11452
rect 39216 11392 39280 11396
rect 39296 11452 39360 11456
rect 39296 11396 39300 11452
rect 39300 11396 39356 11452
rect 39356 11396 39360 11452
rect 39296 11392 39360 11396
rect 39376 11452 39440 11456
rect 39376 11396 39380 11452
rect 39380 11396 39436 11452
rect 39436 11396 39440 11452
rect 39376 11392 39440 11396
rect 39456 11452 39520 11456
rect 39456 11396 39460 11452
rect 39460 11396 39516 11452
rect 39516 11396 39520 11452
rect 39456 11392 39520 11396
rect 49216 11452 49280 11456
rect 49216 11396 49220 11452
rect 49220 11396 49276 11452
rect 49276 11396 49280 11452
rect 49216 11392 49280 11396
rect 49296 11452 49360 11456
rect 49296 11396 49300 11452
rect 49300 11396 49356 11452
rect 49356 11396 49360 11452
rect 49296 11392 49360 11396
rect 49376 11452 49440 11456
rect 49376 11396 49380 11452
rect 49380 11396 49436 11452
rect 49436 11396 49440 11452
rect 49376 11392 49440 11396
rect 49456 11452 49520 11456
rect 49456 11396 49460 11452
rect 49460 11396 49516 11452
rect 49516 11396 49520 11452
rect 49456 11392 49520 11396
rect 59216 11452 59280 11456
rect 59216 11396 59220 11452
rect 59220 11396 59276 11452
rect 59276 11396 59280 11452
rect 59216 11392 59280 11396
rect 59296 11452 59360 11456
rect 59296 11396 59300 11452
rect 59300 11396 59356 11452
rect 59356 11396 59360 11452
rect 59296 11392 59360 11396
rect 59376 11452 59440 11456
rect 59376 11396 59380 11452
rect 59380 11396 59436 11452
rect 59436 11396 59440 11452
rect 59376 11392 59440 11396
rect 59456 11452 59520 11456
rect 59456 11396 59460 11452
rect 59460 11396 59516 11452
rect 59516 11396 59520 11452
rect 59456 11392 59520 11396
rect 13860 11384 13924 11388
rect 13860 11328 13874 11384
rect 13874 11328 13924 11384
rect 13860 11324 13924 11328
rect 9628 11248 9692 11252
rect 9628 11192 9678 11248
rect 9678 11192 9692 11248
rect 9628 11188 9692 11192
rect 42564 11052 42628 11116
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 14216 10908 14280 10912
rect 14216 10852 14220 10908
rect 14220 10852 14276 10908
rect 14276 10852 14280 10908
rect 14216 10848 14280 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 44216 10908 44280 10912
rect 44216 10852 44220 10908
rect 44220 10852 44276 10908
rect 44276 10852 44280 10908
rect 44216 10848 44280 10852
rect 44296 10908 44360 10912
rect 44296 10852 44300 10908
rect 44300 10852 44356 10908
rect 44356 10852 44360 10908
rect 44296 10848 44360 10852
rect 44376 10908 44440 10912
rect 44376 10852 44380 10908
rect 44380 10852 44436 10908
rect 44436 10852 44440 10908
rect 44376 10848 44440 10852
rect 44456 10908 44520 10912
rect 44456 10852 44460 10908
rect 44460 10852 44516 10908
rect 44516 10852 44520 10908
rect 44456 10848 44520 10852
rect 54216 10908 54280 10912
rect 54216 10852 54220 10908
rect 54220 10852 54276 10908
rect 54276 10852 54280 10908
rect 54216 10848 54280 10852
rect 54296 10908 54360 10912
rect 54296 10852 54300 10908
rect 54300 10852 54356 10908
rect 54356 10852 54360 10908
rect 54296 10848 54360 10852
rect 54376 10908 54440 10912
rect 54376 10852 54380 10908
rect 54380 10852 54436 10908
rect 54436 10852 54440 10908
rect 54376 10848 54440 10852
rect 54456 10908 54520 10912
rect 54456 10852 54460 10908
rect 54460 10852 54516 10908
rect 54516 10852 54520 10908
rect 54456 10848 54520 10852
rect 64216 10908 64280 10912
rect 64216 10852 64220 10908
rect 64220 10852 64276 10908
rect 64276 10852 64280 10908
rect 64216 10848 64280 10852
rect 64296 10908 64360 10912
rect 64296 10852 64300 10908
rect 64300 10852 64356 10908
rect 64356 10852 64360 10908
rect 64296 10848 64360 10852
rect 64376 10908 64440 10912
rect 64376 10852 64380 10908
rect 64380 10852 64436 10908
rect 64436 10852 64440 10908
rect 64376 10848 64440 10852
rect 64456 10908 64520 10912
rect 64456 10852 64460 10908
rect 64460 10852 64516 10908
rect 64516 10852 64520 10908
rect 64456 10848 64520 10852
rect 14780 10508 14844 10572
rect 29216 10569 29280 10633
rect 29296 10569 29360 10633
rect 29376 10569 29440 10633
rect 29456 10569 29520 10633
rect 29216 10489 29280 10553
rect 29296 10489 29360 10553
rect 29376 10489 29440 10553
rect 29456 10489 29520 10553
rect 40356 10508 40420 10572
rect 29216 10409 29280 10473
rect 29296 10409 29360 10473
rect 29376 10409 29440 10473
rect 29456 10409 29520 10473
rect 9216 10364 9280 10368
rect 9216 10308 9220 10364
rect 9220 10308 9276 10364
rect 9276 10308 9280 10364
rect 9216 10304 9280 10308
rect 9296 10364 9360 10368
rect 9296 10308 9300 10364
rect 9300 10308 9356 10364
rect 9356 10308 9360 10364
rect 9296 10304 9360 10308
rect 9376 10364 9440 10368
rect 9376 10308 9380 10364
rect 9380 10308 9436 10364
rect 9436 10308 9440 10364
rect 9376 10304 9440 10308
rect 9456 10364 9520 10368
rect 9456 10308 9460 10364
rect 9460 10308 9516 10364
rect 9516 10308 9520 10364
rect 9456 10304 9520 10308
rect 29216 10329 29280 10393
rect 29296 10329 29360 10393
rect 29376 10329 29440 10393
rect 29456 10329 29520 10393
rect 39216 10364 39280 10368
rect 39216 10308 39220 10364
rect 39220 10308 39276 10364
rect 39276 10308 39280 10364
rect 39216 10304 39280 10308
rect 39296 10364 39360 10368
rect 39296 10308 39300 10364
rect 39300 10308 39356 10364
rect 39356 10308 39360 10364
rect 39296 10304 39360 10308
rect 39376 10364 39440 10368
rect 39376 10308 39380 10364
rect 39380 10308 39436 10364
rect 39436 10308 39440 10364
rect 39376 10304 39440 10308
rect 39456 10364 39520 10368
rect 39456 10308 39460 10364
rect 39460 10308 39516 10364
rect 39516 10308 39520 10364
rect 39456 10304 39520 10308
rect 49216 10364 49280 10368
rect 49216 10308 49220 10364
rect 49220 10308 49276 10364
rect 49276 10308 49280 10364
rect 49216 10304 49280 10308
rect 49296 10364 49360 10368
rect 49296 10308 49300 10364
rect 49300 10308 49356 10364
rect 49356 10308 49360 10364
rect 49296 10304 49360 10308
rect 49376 10364 49440 10368
rect 49376 10308 49380 10364
rect 49380 10308 49436 10364
rect 49436 10308 49440 10364
rect 49376 10304 49440 10308
rect 49456 10364 49520 10368
rect 49456 10308 49460 10364
rect 49460 10308 49516 10364
rect 49516 10308 49520 10364
rect 49456 10304 49520 10308
rect 59216 10364 59280 10368
rect 59216 10308 59220 10364
rect 59220 10308 59276 10364
rect 59276 10308 59280 10364
rect 59216 10304 59280 10308
rect 59296 10364 59360 10368
rect 59296 10308 59300 10364
rect 59300 10308 59356 10364
rect 59356 10308 59360 10364
rect 59296 10304 59360 10308
rect 59376 10364 59440 10368
rect 59376 10308 59380 10364
rect 59380 10308 59436 10364
rect 59436 10308 59440 10364
rect 59376 10304 59440 10308
rect 59456 10364 59520 10368
rect 59456 10308 59460 10364
rect 59460 10308 59516 10364
rect 59516 10308 59520 10364
rect 59456 10304 59520 10308
rect 11652 10024 11716 10028
rect 11652 9968 11666 10024
rect 11666 9968 11716 10024
rect 11652 9964 11716 9968
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 14216 9820 14280 9824
rect 14216 9764 14220 9820
rect 14220 9764 14276 9820
rect 14276 9764 14280 9820
rect 14216 9760 14280 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 38884 9420 38948 9484
rect 14780 9284 14844 9348
rect 9216 9276 9280 9280
rect 9216 9220 9220 9276
rect 9220 9220 9276 9276
rect 9276 9220 9280 9276
rect 9216 9216 9280 9220
rect 9296 9276 9360 9280
rect 9296 9220 9300 9276
rect 9300 9220 9356 9276
rect 9356 9220 9360 9276
rect 9296 9216 9360 9220
rect 9376 9276 9440 9280
rect 9376 9220 9380 9276
rect 9380 9220 9436 9276
rect 9436 9220 9440 9276
rect 9376 9216 9440 9220
rect 9456 9276 9520 9280
rect 9456 9220 9460 9276
rect 9460 9220 9516 9276
rect 9516 9220 9520 9276
rect 9456 9216 9520 9220
rect 14044 9072 14108 9076
rect 14044 9016 14094 9072
rect 14094 9016 14108 9072
rect 14044 9012 14108 9016
rect 14596 8876 14660 8940
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 14216 8732 14280 8736
rect 14216 8676 14220 8732
rect 14220 8676 14276 8732
rect 14276 8676 14280 8732
rect 14216 8672 14280 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 12204 8528 12268 8532
rect 12204 8472 12254 8528
rect 12254 8472 12268 8528
rect 12204 8468 12268 8472
rect 24216 9294 24280 9358
rect 24296 9294 24360 9358
rect 24376 9294 24440 9358
rect 24456 9294 24520 9358
rect 24216 9214 24280 9278
rect 24296 9214 24360 9278
rect 24376 9214 24440 9278
rect 24456 9214 24520 9278
rect 24216 9134 24280 9198
rect 24296 9134 24360 9198
rect 24376 9134 24440 9198
rect 24456 9134 24520 9198
rect 24216 9054 24280 9118
rect 24296 9054 24360 9118
rect 24376 9054 24440 9118
rect 24456 9054 24520 9118
rect 34216 9294 34280 9358
rect 34296 9294 34360 9358
rect 34376 9294 34440 9358
rect 34456 9294 34520 9358
rect 34216 9214 34280 9278
rect 34296 9214 34360 9278
rect 34376 9214 34440 9278
rect 34456 9214 34520 9278
rect 39216 9276 39280 9280
rect 39216 9220 39220 9276
rect 39220 9220 39276 9276
rect 39276 9220 39280 9276
rect 39216 9216 39280 9220
rect 39296 9276 39360 9280
rect 39296 9220 39300 9276
rect 39300 9220 39356 9276
rect 39356 9220 39360 9276
rect 39296 9216 39360 9220
rect 39376 9276 39440 9280
rect 39376 9220 39380 9276
rect 39380 9220 39436 9276
rect 39436 9220 39440 9276
rect 39376 9216 39440 9220
rect 39456 9276 39520 9280
rect 39456 9220 39460 9276
rect 39460 9220 39516 9276
rect 39516 9220 39520 9276
rect 39456 9216 39520 9220
rect 44216 9820 44280 9824
rect 44216 9764 44220 9820
rect 44220 9764 44276 9820
rect 44276 9764 44280 9820
rect 44216 9760 44280 9764
rect 44296 9820 44360 9824
rect 44296 9764 44300 9820
rect 44300 9764 44356 9820
rect 44356 9764 44360 9820
rect 44296 9760 44360 9764
rect 44376 9820 44440 9824
rect 44376 9764 44380 9820
rect 44380 9764 44436 9820
rect 44436 9764 44440 9820
rect 44376 9760 44440 9764
rect 44456 9820 44520 9824
rect 44456 9764 44460 9820
rect 44460 9764 44516 9820
rect 44516 9764 44520 9820
rect 44456 9760 44520 9764
rect 54216 9820 54280 9824
rect 54216 9764 54220 9820
rect 54220 9764 54276 9820
rect 54276 9764 54280 9820
rect 54216 9760 54280 9764
rect 54296 9820 54360 9824
rect 54296 9764 54300 9820
rect 54300 9764 54356 9820
rect 54356 9764 54360 9820
rect 54296 9760 54360 9764
rect 54376 9820 54440 9824
rect 54376 9764 54380 9820
rect 54380 9764 54436 9820
rect 54436 9764 54440 9820
rect 54376 9760 54440 9764
rect 54456 9820 54520 9824
rect 54456 9764 54460 9820
rect 54460 9764 54516 9820
rect 54516 9764 54520 9820
rect 54456 9760 54520 9764
rect 64216 9820 64280 9824
rect 64216 9764 64220 9820
rect 64220 9764 64276 9820
rect 64276 9764 64280 9820
rect 64216 9760 64280 9764
rect 64296 9820 64360 9824
rect 64296 9764 64300 9820
rect 64300 9764 64356 9820
rect 64356 9764 64360 9820
rect 64296 9760 64360 9764
rect 64376 9820 64440 9824
rect 64376 9764 64380 9820
rect 64380 9764 64436 9820
rect 64436 9764 64440 9820
rect 64376 9760 64440 9764
rect 64456 9820 64520 9824
rect 64456 9764 64460 9820
rect 64460 9764 64516 9820
rect 64516 9764 64520 9820
rect 64456 9760 64520 9764
rect 43852 9420 43916 9484
rect 49216 9276 49280 9280
rect 49216 9220 49220 9276
rect 49220 9220 49276 9276
rect 49276 9220 49280 9276
rect 49216 9216 49280 9220
rect 49296 9276 49360 9280
rect 49296 9220 49300 9276
rect 49300 9220 49356 9276
rect 49356 9220 49360 9276
rect 49296 9216 49360 9220
rect 49376 9276 49440 9280
rect 49376 9220 49380 9276
rect 49380 9220 49436 9276
rect 49436 9220 49440 9276
rect 49376 9216 49440 9220
rect 49456 9276 49520 9280
rect 49456 9220 49460 9276
rect 49460 9220 49516 9276
rect 49516 9220 49520 9276
rect 49456 9216 49520 9220
rect 59216 9276 59280 9280
rect 59216 9220 59220 9276
rect 59220 9220 59276 9276
rect 59276 9220 59280 9276
rect 59216 9216 59280 9220
rect 59296 9276 59360 9280
rect 59296 9220 59300 9276
rect 59300 9220 59356 9276
rect 59356 9220 59360 9276
rect 59296 9216 59360 9220
rect 59376 9276 59440 9280
rect 59376 9220 59380 9276
rect 59380 9220 59436 9276
rect 59436 9220 59440 9276
rect 59376 9216 59440 9220
rect 59456 9276 59520 9280
rect 59456 9220 59460 9276
rect 59460 9220 59516 9276
rect 59516 9220 59520 9276
rect 59456 9216 59520 9220
rect 34216 9134 34280 9198
rect 34296 9134 34360 9198
rect 34376 9134 34440 9198
rect 34456 9134 34520 9198
rect 40908 9148 40972 9212
rect 34216 9054 34280 9118
rect 34296 9054 34360 9118
rect 34376 9054 34440 9118
rect 34456 9054 34520 9118
rect 40172 9012 40236 9076
rect 41460 9012 41524 9076
rect 39988 8876 40052 8940
rect 42380 8936 42444 8940
rect 42380 8880 42394 8936
rect 42394 8880 42444 8936
rect 42380 8876 42444 8880
rect 44036 8876 44100 8940
rect 44216 8732 44280 8736
rect 44216 8676 44220 8732
rect 44220 8676 44276 8732
rect 44276 8676 44280 8732
rect 44216 8672 44280 8676
rect 44296 8732 44360 8736
rect 44296 8676 44300 8732
rect 44300 8676 44356 8732
rect 44356 8676 44360 8732
rect 44296 8672 44360 8676
rect 44376 8732 44440 8736
rect 44376 8676 44380 8732
rect 44380 8676 44436 8732
rect 44436 8676 44440 8732
rect 44376 8672 44440 8676
rect 44456 8732 44520 8736
rect 44456 8676 44460 8732
rect 44460 8676 44516 8732
rect 44516 8676 44520 8732
rect 44456 8672 44520 8676
rect 54216 8732 54280 8736
rect 54216 8676 54220 8732
rect 54220 8676 54276 8732
rect 54276 8676 54280 8732
rect 54216 8672 54280 8676
rect 54296 8732 54360 8736
rect 54296 8676 54300 8732
rect 54300 8676 54356 8732
rect 54356 8676 54360 8732
rect 54296 8672 54360 8676
rect 54376 8732 54440 8736
rect 54376 8676 54380 8732
rect 54380 8676 54436 8732
rect 54436 8676 54440 8732
rect 54376 8672 54440 8676
rect 54456 8732 54520 8736
rect 54456 8676 54460 8732
rect 54460 8676 54516 8732
rect 54516 8676 54520 8732
rect 54456 8672 54520 8676
rect 64216 8732 64280 8736
rect 64216 8676 64220 8732
rect 64220 8676 64276 8732
rect 64276 8676 64280 8732
rect 64216 8672 64280 8676
rect 64296 8732 64360 8736
rect 64296 8676 64300 8732
rect 64300 8676 64356 8732
rect 64356 8676 64360 8732
rect 64296 8672 64360 8676
rect 64376 8732 64440 8736
rect 64376 8676 64380 8732
rect 64380 8676 64436 8732
rect 64436 8676 64440 8732
rect 64376 8672 64440 8676
rect 64456 8732 64520 8736
rect 64456 8676 64460 8732
rect 64460 8676 64516 8732
rect 64516 8676 64520 8732
rect 64456 8672 64520 8676
rect 40356 8468 40420 8532
rect 44956 8468 45020 8532
rect 41276 8256 41340 8260
rect 41276 8200 41326 8256
rect 41326 8200 41340 8256
rect 41276 8196 41340 8200
rect 9216 8188 9280 8192
rect 9216 8132 9220 8188
rect 9220 8132 9276 8188
rect 9276 8132 9280 8188
rect 9216 8128 9280 8132
rect 9296 8188 9360 8192
rect 9296 8132 9300 8188
rect 9300 8132 9356 8188
rect 9356 8132 9360 8188
rect 9296 8128 9360 8132
rect 9376 8188 9440 8192
rect 9376 8132 9380 8188
rect 9380 8132 9436 8188
rect 9436 8132 9440 8188
rect 9376 8128 9440 8132
rect 9456 8188 9520 8192
rect 9456 8132 9460 8188
rect 9460 8132 9516 8188
rect 9516 8132 9520 8188
rect 9456 8128 9520 8132
rect 39216 8188 39280 8192
rect 39216 8132 39220 8188
rect 39220 8132 39276 8188
rect 39276 8132 39280 8188
rect 39216 8128 39280 8132
rect 39296 8188 39360 8192
rect 39296 8132 39300 8188
rect 39300 8132 39356 8188
rect 39356 8132 39360 8188
rect 39296 8128 39360 8132
rect 39376 8188 39440 8192
rect 39376 8132 39380 8188
rect 39380 8132 39436 8188
rect 39436 8132 39440 8188
rect 39376 8128 39440 8132
rect 39456 8188 39520 8192
rect 39456 8132 39460 8188
rect 39460 8132 39516 8188
rect 39516 8132 39520 8188
rect 39456 8128 39520 8132
rect 49216 8188 49280 8192
rect 49216 8132 49220 8188
rect 49220 8132 49276 8188
rect 49276 8132 49280 8188
rect 49216 8128 49280 8132
rect 49296 8188 49360 8192
rect 49296 8132 49300 8188
rect 49300 8132 49356 8188
rect 49356 8132 49360 8188
rect 49296 8128 49360 8132
rect 49376 8188 49440 8192
rect 49376 8132 49380 8188
rect 49380 8132 49436 8188
rect 49436 8132 49440 8188
rect 49376 8128 49440 8132
rect 49456 8188 49520 8192
rect 49456 8132 49460 8188
rect 49460 8132 49516 8188
rect 49516 8132 49520 8188
rect 49456 8128 49520 8132
rect 59216 8188 59280 8192
rect 59216 8132 59220 8188
rect 59220 8132 59276 8188
rect 59276 8132 59280 8188
rect 59216 8128 59280 8132
rect 59296 8188 59360 8192
rect 59296 8132 59300 8188
rect 59300 8132 59356 8188
rect 59356 8132 59360 8188
rect 59296 8128 59360 8132
rect 59376 8188 59440 8192
rect 59376 8132 59380 8188
rect 59380 8132 59436 8188
rect 59436 8132 59440 8188
rect 59376 8128 59440 8132
rect 59456 8188 59520 8192
rect 59456 8132 59460 8188
rect 59460 8132 59516 8188
rect 59516 8132 59520 8188
rect 59456 8128 59520 8132
rect 29216 8019 29280 8083
rect 29296 8019 29360 8083
rect 29376 8019 29440 8083
rect 29456 8019 29520 8083
rect 29216 7939 29280 8003
rect 29296 7939 29360 8003
rect 29376 7939 29440 8003
rect 29456 7939 29520 8003
rect 29216 7859 29280 7923
rect 29296 7859 29360 7923
rect 29376 7859 29440 7923
rect 29456 7859 29520 7923
rect 29216 7779 29280 7843
rect 29296 7779 29360 7843
rect 29376 7779 29440 7843
rect 29456 7779 29520 7843
rect 46796 7848 46860 7852
rect 46796 7792 46846 7848
rect 46846 7792 46860 7848
rect 46796 7788 46860 7792
rect 13676 7712 13740 7716
rect 13676 7656 13690 7712
rect 13690 7656 13740 7712
rect 13676 7652 13740 7656
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 14216 7644 14280 7648
rect 14216 7588 14220 7644
rect 14220 7588 14276 7644
rect 14276 7588 14280 7644
rect 14216 7584 14280 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 44216 7644 44280 7648
rect 44216 7588 44220 7644
rect 44220 7588 44276 7644
rect 44276 7588 44280 7644
rect 44216 7584 44280 7588
rect 44296 7644 44360 7648
rect 44296 7588 44300 7644
rect 44300 7588 44356 7644
rect 44356 7588 44360 7644
rect 44296 7584 44360 7588
rect 44376 7644 44440 7648
rect 44376 7588 44380 7644
rect 44380 7588 44436 7644
rect 44436 7588 44440 7644
rect 44376 7584 44440 7588
rect 44456 7644 44520 7648
rect 44456 7588 44460 7644
rect 44460 7588 44516 7644
rect 44516 7588 44520 7644
rect 44456 7584 44520 7588
rect 54216 7644 54280 7648
rect 54216 7588 54220 7644
rect 54220 7588 54276 7644
rect 54276 7588 54280 7644
rect 54216 7584 54280 7588
rect 54296 7644 54360 7648
rect 54296 7588 54300 7644
rect 54300 7588 54356 7644
rect 54356 7588 54360 7644
rect 54296 7584 54360 7588
rect 54376 7644 54440 7648
rect 54376 7588 54380 7644
rect 54380 7588 54436 7644
rect 54436 7588 54440 7644
rect 54376 7584 54440 7588
rect 54456 7644 54520 7648
rect 54456 7588 54460 7644
rect 54460 7588 54516 7644
rect 54516 7588 54520 7644
rect 54456 7584 54520 7588
rect 64216 7644 64280 7648
rect 64216 7588 64220 7644
rect 64220 7588 64276 7644
rect 64276 7588 64280 7644
rect 64216 7584 64280 7588
rect 64296 7644 64360 7648
rect 64296 7588 64300 7644
rect 64300 7588 64356 7644
rect 64356 7588 64360 7644
rect 64296 7584 64360 7588
rect 64376 7644 64440 7648
rect 64376 7588 64380 7644
rect 64380 7588 64436 7644
rect 64436 7588 64440 7644
rect 64376 7584 64440 7588
rect 64456 7644 64520 7648
rect 64456 7588 64460 7644
rect 64460 7588 64516 7644
rect 64516 7588 64520 7644
rect 64456 7584 64520 7588
rect 38884 7380 38948 7444
rect 5396 7108 5460 7172
rect 9216 7100 9280 7104
rect 9216 7044 9220 7100
rect 9220 7044 9276 7100
rect 9276 7044 9280 7100
rect 9216 7040 9280 7044
rect 9296 7100 9360 7104
rect 9296 7044 9300 7100
rect 9300 7044 9356 7100
rect 9356 7044 9360 7100
rect 9296 7040 9360 7044
rect 9376 7100 9440 7104
rect 9376 7044 9380 7100
rect 9380 7044 9436 7100
rect 9436 7044 9440 7100
rect 9376 7040 9440 7044
rect 9456 7100 9520 7104
rect 9456 7044 9460 7100
rect 9460 7044 9516 7100
rect 9516 7044 9520 7100
rect 9456 7040 9520 7044
rect 39216 7100 39280 7104
rect 39216 7044 39220 7100
rect 39220 7044 39276 7100
rect 39276 7044 39280 7100
rect 39216 7040 39280 7044
rect 39296 7100 39360 7104
rect 39296 7044 39300 7100
rect 39300 7044 39356 7100
rect 39356 7044 39360 7100
rect 39296 7040 39360 7044
rect 39376 7100 39440 7104
rect 39376 7044 39380 7100
rect 39380 7044 39436 7100
rect 39436 7044 39440 7100
rect 39376 7040 39440 7044
rect 39456 7100 39520 7104
rect 39456 7044 39460 7100
rect 39460 7044 39516 7100
rect 39516 7044 39520 7100
rect 39456 7040 39520 7044
rect 49216 7100 49280 7104
rect 49216 7044 49220 7100
rect 49220 7044 49276 7100
rect 49276 7044 49280 7100
rect 49216 7040 49280 7044
rect 49296 7100 49360 7104
rect 49296 7044 49300 7100
rect 49300 7044 49356 7100
rect 49356 7044 49360 7100
rect 49296 7040 49360 7044
rect 49376 7100 49440 7104
rect 49376 7044 49380 7100
rect 49380 7044 49436 7100
rect 49436 7044 49440 7100
rect 49376 7040 49440 7044
rect 49456 7100 49520 7104
rect 49456 7044 49460 7100
rect 49460 7044 49516 7100
rect 49516 7044 49520 7100
rect 49456 7040 49520 7044
rect 59216 7100 59280 7104
rect 59216 7044 59220 7100
rect 59220 7044 59276 7100
rect 59276 7044 59280 7100
rect 59216 7040 59280 7044
rect 59296 7100 59360 7104
rect 59296 7044 59300 7100
rect 59300 7044 59356 7100
rect 59356 7044 59360 7100
rect 59296 7040 59360 7044
rect 59376 7100 59440 7104
rect 59376 7044 59380 7100
rect 59380 7044 59436 7100
rect 59436 7044 59440 7100
rect 59376 7040 59440 7044
rect 59456 7100 59520 7104
rect 59456 7044 59460 7100
rect 59460 7044 59516 7100
rect 59516 7044 59520 7100
rect 59456 7040 59520 7044
rect 39620 7032 39684 7036
rect 39620 6976 39670 7032
rect 39670 6976 39684 7032
rect 39620 6972 39684 6976
rect 24216 6745 24280 6809
rect 24296 6745 24360 6809
rect 24376 6745 24440 6809
rect 24456 6745 24520 6809
rect 24216 6665 24280 6729
rect 24296 6665 24360 6729
rect 24376 6665 24440 6729
rect 24456 6665 24520 6729
rect 24216 6585 24280 6649
rect 24296 6585 24360 6649
rect 24376 6585 24440 6649
rect 24456 6585 24520 6649
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 14216 6556 14280 6560
rect 14216 6500 14220 6556
rect 14220 6500 14276 6556
rect 14276 6500 14280 6556
rect 14216 6496 14280 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 24216 6505 24280 6569
rect 24296 6505 24360 6569
rect 24376 6505 24440 6569
rect 24456 6505 24520 6569
rect 34216 6745 34280 6809
rect 34296 6745 34360 6809
rect 34376 6745 34440 6809
rect 34456 6745 34520 6809
rect 34216 6665 34280 6729
rect 34296 6665 34360 6729
rect 34376 6665 34440 6729
rect 34456 6665 34520 6729
rect 34216 6585 34280 6649
rect 34296 6585 34360 6649
rect 34376 6585 34440 6649
rect 34456 6585 34520 6649
rect 34216 6505 34280 6569
rect 34296 6505 34360 6569
rect 34376 6505 34440 6569
rect 34456 6505 34520 6569
rect 44216 6556 44280 6560
rect 44216 6500 44220 6556
rect 44220 6500 44276 6556
rect 44276 6500 44280 6556
rect 44216 6496 44280 6500
rect 44296 6556 44360 6560
rect 44296 6500 44300 6556
rect 44300 6500 44356 6556
rect 44356 6500 44360 6556
rect 44296 6496 44360 6500
rect 44376 6556 44440 6560
rect 44376 6500 44380 6556
rect 44380 6500 44436 6556
rect 44436 6500 44440 6556
rect 44376 6496 44440 6500
rect 44456 6556 44520 6560
rect 44456 6500 44460 6556
rect 44460 6500 44516 6556
rect 44516 6500 44520 6556
rect 44456 6496 44520 6500
rect 54216 6556 54280 6560
rect 54216 6500 54220 6556
rect 54220 6500 54276 6556
rect 54276 6500 54280 6556
rect 54216 6496 54280 6500
rect 54296 6556 54360 6560
rect 54296 6500 54300 6556
rect 54300 6500 54356 6556
rect 54356 6500 54360 6556
rect 54296 6496 54360 6500
rect 54376 6556 54440 6560
rect 54376 6500 54380 6556
rect 54380 6500 54436 6556
rect 54436 6500 54440 6556
rect 54376 6496 54440 6500
rect 54456 6556 54520 6560
rect 54456 6500 54460 6556
rect 54460 6500 54516 6556
rect 54516 6500 54520 6556
rect 54456 6496 54520 6500
rect 64216 6556 64280 6560
rect 64216 6500 64220 6556
rect 64220 6500 64276 6556
rect 64276 6500 64280 6556
rect 64216 6496 64280 6500
rect 64296 6556 64360 6560
rect 64296 6500 64300 6556
rect 64300 6500 64356 6556
rect 64356 6500 64360 6556
rect 64296 6496 64360 6500
rect 64376 6556 64440 6560
rect 64376 6500 64380 6556
rect 64380 6500 64436 6556
rect 64436 6500 64440 6556
rect 64376 6496 64440 6500
rect 64456 6556 64520 6560
rect 64456 6500 64460 6556
rect 64460 6500 64516 6556
rect 64516 6500 64520 6556
rect 64456 6496 64520 6500
rect 14596 6292 14660 6356
rect 30420 6020 30484 6084
rect 42012 6020 42076 6084
rect 9216 6012 9280 6016
rect 9216 5956 9220 6012
rect 9220 5956 9276 6012
rect 9276 5956 9280 6012
rect 9216 5952 9280 5956
rect 9296 6012 9360 6016
rect 9296 5956 9300 6012
rect 9300 5956 9356 6012
rect 9356 5956 9360 6012
rect 9296 5952 9360 5956
rect 9376 6012 9440 6016
rect 9376 5956 9380 6012
rect 9380 5956 9436 6012
rect 9436 5956 9440 6012
rect 9376 5952 9440 5956
rect 9456 6012 9520 6016
rect 9456 5956 9460 6012
rect 9460 5956 9516 6012
rect 9516 5956 9520 6012
rect 9456 5952 9520 5956
rect 39216 6012 39280 6016
rect 39216 5956 39220 6012
rect 39220 5956 39276 6012
rect 39276 5956 39280 6012
rect 39216 5952 39280 5956
rect 39296 6012 39360 6016
rect 39296 5956 39300 6012
rect 39300 5956 39356 6012
rect 39356 5956 39360 6012
rect 39296 5952 39360 5956
rect 39376 6012 39440 6016
rect 39376 5956 39380 6012
rect 39380 5956 39436 6012
rect 39436 5956 39440 6012
rect 39376 5952 39440 5956
rect 39456 6012 39520 6016
rect 39456 5956 39460 6012
rect 39460 5956 39516 6012
rect 39516 5956 39520 6012
rect 39456 5952 39520 5956
rect 49216 6012 49280 6016
rect 49216 5956 49220 6012
rect 49220 5956 49276 6012
rect 49276 5956 49280 6012
rect 49216 5952 49280 5956
rect 49296 6012 49360 6016
rect 49296 5956 49300 6012
rect 49300 5956 49356 6012
rect 49356 5956 49360 6012
rect 49296 5952 49360 5956
rect 49376 6012 49440 6016
rect 49376 5956 49380 6012
rect 49380 5956 49436 6012
rect 49436 5956 49440 6012
rect 49376 5952 49440 5956
rect 49456 6012 49520 6016
rect 49456 5956 49460 6012
rect 49460 5956 49516 6012
rect 49516 5956 49520 6012
rect 49456 5952 49520 5956
rect 59216 6012 59280 6016
rect 59216 5956 59220 6012
rect 59220 5956 59276 6012
rect 59276 5956 59280 6012
rect 59216 5952 59280 5956
rect 59296 6012 59360 6016
rect 59296 5956 59300 6012
rect 59300 5956 59356 6012
rect 59356 5956 59360 6012
rect 59296 5952 59360 5956
rect 59376 6012 59440 6016
rect 59376 5956 59380 6012
rect 59380 5956 59436 6012
rect 59436 5956 59440 6012
rect 59376 5952 59440 5956
rect 59456 6012 59520 6016
rect 59456 5956 59460 6012
rect 59460 5956 59516 6012
rect 59516 5956 59520 6012
rect 59456 5952 59520 5956
rect 27660 5884 27724 5948
rect 46612 5808 46676 5812
rect 46612 5752 46662 5808
rect 46662 5752 46676 5808
rect 46612 5748 46676 5752
rect 30604 5476 30668 5540
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 14216 5468 14280 5472
rect 14216 5412 14220 5468
rect 14220 5412 14276 5468
rect 14276 5412 14280 5468
rect 14216 5408 14280 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 44216 5468 44280 5472
rect 44216 5412 44220 5468
rect 44220 5412 44276 5468
rect 44276 5412 44280 5468
rect 44216 5408 44280 5412
rect 44296 5468 44360 5472
rect 44296 5412 44300 5468
rect 44300 5412 44356 5468
rect 44356 5412 44360 5468
rect 44296 5408 44360 5412
rect 44376 5468 44440 5472
rect 44376 5412 44380 5468
rect 44380 5412 44436 5468
rect 44436 5412 44440 5468
rect 44376 5408 44440 5412
rect 44456 5468 44520 5472
rect 44456 5412 44460 5468
rect 44460 5412 44516 5468
rect 44516 5412 44520 5468
rect 44456 5408 44520 5412
rect 54216 5468 54280 5472
rect 54216 5412 54220 5468
rect 54220 5412 54276 5468
rect 54276 5412 54280 5468
rect 54216 5408 54280 5412
rect 54296 5468 54360 5472
rect 54296 5412 54300 5468
rect 54300 5412 54356 5468
rect 54356 5412 54360 5468
rect 54296 5408 54360 5412
rect 54376 5468 54440 5472
rect 54376 5412 54380 5468
rect 54380 5412 54436 5468
rect 54436 5412 54440 5468
rect 54376 5408 54440 5412
rect 54456 5468 54520 5472
rect 54456 5412 54460 5468
rect 54460 5412 54516 5468
rect 54516 5412 54520 5468
rect 54456 5408 54520 5412
rect 64216 5468 64280 5472
rect 64216 5412 64220 5468
rect 64220 5412 64276 5468
rect 64276 5412 64280 5468
rect 64216 5408 64280 5412
rect 64296 5468 64360 5472
rect 64296 5412 64300 5468
rect 64300 5412 64356 5468
rect 64356 5412 64360 5468
rect 64296 5408 64360 5412
rect 64376 5468 64440 5472
rect 64376 5412 64380 5468
rect 64380 5412 64436 5468
rect 64436 5412 64440 5468
rect 64376 5408 64440 5412
rect 64456 5468 64520 5472
rect 64456 5412 64460 5468
rect 64460 5412 64516 5468
rect 64516 5412 64520 5468
rect 64456 5408 64520 5412
rect 31892 5340 31956 5404
rect 30052 5204 30116 5268
rect 55996 5264 56060 5268
rect 55996 5208 56010 5264
rect 56010 5208 56060 5264
rect 55996 5204 56060 5208
rect 5396 5128 5460 5132
rect 5396 5072 5446 5128
rect 5446 5072 5460 5128
rect 5396 5068 5460 5072
rect 53604 4932 53668 4996
rect 54892 4992 54956 4996
rect 54892 4936 54942 4992
rect 54942 4936 54956 4992
rect 54892 4932 54956 4936
rect 9216 4924 9280 4928
rect 9216 4868 9220 4924
rect 9220 4868 9276 4924
rect 9276 4868 9280 4924
rect 9216 4864 9280 4868
rect 9296 4924 9360 4928
rect 9296 4868 9300 4924
rect 9300 4868 9356 4924
rect 9356 4868 9360 4924
rect 9296 4864 9360 4868
rect 9376 4924 9440 4928
rect 9376 4868 9380 4924
rect 9380 4868 9436 4924
rect 9436 4868 9440 4924
rect 9376 4864 9440 4868
rect 9456 4924 9520 4928
rect 9456 4868 9460 4924
rect 9460 4868 9516 4924
rect 9516 4868 9520 4924
rect 9456 4864 9520 4868
rect 39216 4924 39280 4928
rect 39216 4868 39220 4924
rect 39220 4868 39276 4924
rect 39276 4868 39280 4924
rect 39216 4864 39280 4868
rect 39296 4924 39360 4928
rect 39296 4868 39300 4924
rect 39300 4868 39356 4924
rect 39356 4868 39360 4924
rect 39296 4864 39360 4868
rect 39376 4924 39440 4928
rect 39376 4868 39380 4924
rect 39380 4868 39436 4924
rect 39436 4868 39440 4924
rect 39376 4864 39440 4868
rect 39456 4924 39520 4928
rect 39456 4868 39460 4924
rect 39460 4868 39516 4924
rect 39516 4868 39520 4924
rect 39456 4864 39520 4868
rect 49216 4924 49280 4928
rect 49216 4868 49220 4924
rect 49220 4868 49276 4924
rect 49276 4868 49280 4924
rect 49216 4864 49280 4868
rect 49296 4924 49360 4928
rect 49296 4868 49300 4924
rect 49300 4868 49356 4924
rect 49356 4868 49360 4924
rect 49296 4864 49360 4868
rect 49376 4924 49440 4928
rect 49376 4868 49380 4924
rect 49380 4868 49436 4924
rect 49436 4868 49440 4924
rect 49376 4864 49440 4868
rect 49456 4924 49520 4928
rect 49456 4868 49460 4924
rect 49460 4868 49516 4924
rect 49516 4868 49520 4924
rect 49456 4864 49520 4868
rect 59216 4924 59280 4928
rect 59216 4868 59220 4924
rect 59220 4868 59276 4924
rect 59276 4868 59280 4924
rect 59216 4864 59280 4868
rect 59296 4924 59360 4928
rect 59296 4868 59300 4924
rect 59300 4868 59356 4924
rect 59356 4868 59360 4924
rect 59296 4864 59360 4868
rect 59376 4924 59440 4928
rect 59376 4868 59380 4924
rect 59380 4868 59436 4924
rect 59436 4868 59440 4924
rect 59376 4864 59440 4868
rect 59456 4924 59520 4928
rect 59456 4868 59460 4924
rect 59460 4868 59516 4924
rect 59516 4868 59520 4924
rect 59456 4864 59520 4868
rect 31156 4660 31220 4724
rect 40908 4660 40972 4724
rect 39988 4524 40052 4588
rect 64644 4584 64708 4588
rect 64644 4528 64694 4584
rect 64694 4528 64708 4584
rect 64644 4524 64708 4528
rect 38884 4388 38948 4452
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 14216 4380 14280 4384
rect 14216 4324 14220 4380
rect 14220 4324 14276 4380
rect 14276 4324 14280 4380
rect 14216 4320 14280 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 44216 4380 44280 4384
rect 44216 4324 44220 4380
rect 44220 4324 44276 4380
rect 44276 4324 44280 4380
rect 44216 4320 44280 4324
rect 44296 4380 44360 4384
rect 44296 4324 44300 4380
rect 44300 4324 44356 4380
rect 44356 4324 44360 4380
rect 44296 4320 44360 4324
rect 44376 4380 44440 4384
rect 44376 4324 44380 4380
rect 44380 4324 44436 4380
rect 44436 4324 44440 4380
rect 44376 4320 44440 4324
rect 44456 4380 44520 4384
rect 44456 4324 44460 4380
rect 44460 4324 44516 4380
rect 44516 4324 44520 4380
rect 44456 4320 44520 4324
rect 54216 4380 54280 4384
rect 54216 4324 54220 4380
rect 54220 4324 54276 4380
rect 54276 4324 54280 4380
rect 54216 4320 54280 4324
rect 54296 4380 54360 4384
rect 54296 4324 54300 4380
rect 54300 4324 54356 4380
rect 54356 4324 54360 4380
rect 54296 4320 54360 4324
rect 54376 4380 54440 4384
rect 54376 4324 54380 4380
rect 54380 4324 54436 4380
rect 54436 4324 54440 4380
rect 54376 4320 54440 4324
rect 54456 4380 54520 4384
rect 54456 4324 54460 4380
rect 54460 4324 54516 4380
rect 54516 4324 54520 4380
rect 54456 4320 54520 4324
rect 64216 4380 64280 4384
rect 64216 4324 64220 4380
rect 64220 4324 64276 4380
rect 64276 4324 64280 4380
rect 64216 4320 64280 4324
rect 64296 4380 64360 4384
rect 64296 4324 64300 4380
rect 64300 4324 64356 4380
rect 64356 4324 64360 4380
rect 64296 4320 64360 4324
rect 64376 4380 64440 4384
rect 64376 4324 64380 4380
rect 64380 4324 64436 4380
rect 64436 4324 64440 4380
rect 64376 4320 64440 4324
rect 64456 4380 64520 4384
rect 64456 4324 64460 4380
rect 64460 4324 64516 4380
rect 64516 4324 64520 4380
rect 64456 4320 64520 4324
rect 11652 3980 11716 4044
rect 13676 3980 13740 4044
rect 16252 4040 16316 4044
rect 16252 3984 16266 4040
rect 16266 3984 16316 4040
rect 16252 3980 16316 3984
rect 14044 3904 14108 3908
rect 49740 3980 49804 4044
rect 14044 3848 14058 3904
rect 14058 3848 14108 3904
rect 14044 3844 14108 3848
rect 9216 3836 9280 3840
rect 9216 3780 9220 3836
rect 9220 3780 9276 3836
rect 9276 3780 9280 3836
rect 9216 3776 9280 3780
rect 9296 3836 9360 3840
rect 9296 3780 9300 3836
rect 9300 3780 9356 3836
rect 9356 3780 9360 3836
rect 9296 3776 9360 3780
rect 9376 3836 9440 3840
rect 9376 3780 9380 3836
rect 9380 3780 9436 3836
rect 9436 3780 9440 3836
rect 9376 3776 9440 3780
rect 9456 3836 9520 3840
rect 9456 3780 9460 3836
rect 9460 3780 9516 3836
rect 9516 3780 9520 3836
rect 9456 3776 9520 3780
rect 9628 3708 9692 3772
rect 12204 3708 12268 3772
rect 13492 3708 13556 3772
rect 38884 3844 38948 3908
rect 39216 3836 39280 3840
rect 39216 3780 39220 3836
rect 39220 3780 39276 3836
rect 39276 3780 39280 3836
rect 39216 3776 39280 3780
rect 39296 3836 39360 3840
rect 39296 3780 39300 3836
rect 39300 3780 39356 3836
rect 39356 3780 39360 3836
rect 39296 3776 39360 3780
rect 39376 3836 39440 3840
rect 39376 3780 39380 3836
rect 39380 3780 39436 3836
rect 39436 3780 39440 3836
rect 39376 3776 39440 3780
rect 39456 3836 39520 3840
rect 39456 3780 39460 3836
rect 39460 3780 39516 3836
rect 39516 3780 39520 3836
rect 39456 3776 39520 3780
rect 49216 3836 49280 3840
rect 49216 3780 49220 3836
rect 49220 3780 49276 3836
rect 49276 3780 49280 3836
rect 49216 3776 49280 3780
rect 49296 3836 49360 3840
rect 49296 3780 49300 3836
rect 49300 3780 49356 3836
rect 49356 3780 49360 3836
rect 49296 3776 49360 3780
rect 49376 3836 49440 3840
rect 49376 3780 49380 3836
rect 49380 3780 49436 3836
rect 49436 3780 49440 3836
rect 49376 3776 49440 3780
rect 49456 3836 49520 3840
rect 49456 3780 49460 3836
rect 49460 3780 49516 3836
rect 49516 3780 49520 3836
rect 49456 3776 49520 3780
rect 59216 3836 59280 3840
rect 59216 3780 59220 3836
rect 59220 3780 59276 3836
rect 59276 3780 59280 3836
rect 59216 3776 59280 3780
rect 59296 3836 59360 3840
rect 59296 3780 59300 3836
rect 59300 3780 59356 3836
rect 59356 3780 59360 3836
rect 59296 3776 59360 3780
rect 59376 3836 59440 3840
rect 59376 3780 59380 3836
rect 59380 3780 59436 3836
rect 59436 3780 59440 3836
rect 59376 3776 59440 3780
rect 59456 3836 59520 3840
rect 59456 3780 59460 3836
rect 59460 3780 59516 3836
rect 59516 3780 59520 3836
rect 59456 3776 59520 3780
rect 28212 3708 28276 3772
rect 33732 3708 33796 3772
rect 28028 3572 28092 3636
rect 44036 3708 44100 3772
rect 55996 3768 56060 3772
rect 55996 3712 56010 3768
rect 56010 3712 56060 3768
rect 55996 3708 56060 3712
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 39068 3300 39132 3364
rect 39804 3300 39868 3364
rect 46796 3300 46860 3364
rect 14216 3292 14280 3296
rect 14216 3236 14220 3292
rect 14220 3236 14276 3292
rect 14276 3236 14280 3292
rect 14216 3232 14280 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 44216 3292 44280 3296
rect 44216 3236 44220 3292
rect 44220 3236 44276 3292
rect 44276 3236 44280 3292
rect 44216 3232 44280 3236
rect 44296 3292 44360 3296
rect 44296 3236 44300 3292
rect 44300 3236 44356 3292
rect 44356 3236 44360 3292
rect 44296 3232 44360 3236
rect 44376 3292 44440 3296
rect 44376 3236 44380 3292
rect 44380 3236 44436 3292
rect 44436 3236 44440 3292
rect 44376 3232 44440 3236
rect 44456 3292 44520 3296
rect 44456 3236 44460 3292
rect 44460 3236 44516 3292
rect 44516 3236 44520 3292
rect 44456 3232 44520 3236
rect 54216 3292 54280 3296
rect 54216 3236 54220 3292
rect 54220 3236 54276 3292
rect 54276 3236 54280 3292
rect 54216 3232 54280 3236
rect 54296 3292 54360 3296
rect 54296 3236 54300 3292
rect 54300 3236 54356 3292
rect 54356 3236 54360 3292
rect 54296 3232 54360 3236
rect 54376 3292 54440 3296
rect 54376 3236 54380 3292
rect 54380 3236 54436 3292
rect 54436 3236 54440 3292
rect 54376 3232 54440 3236
rect 54456 3292 54520 3296
rect 54456 3236 54460 3292
rect 54460 3236 54516 3292
rect 54516 3236 54520 3292
rect 54456 3232 54520 3236
rect 64216 3292 64280 3296
rect 64216 3236 64220 3292
rect 64220 3236 64276 3292
rect 64276 3236 64280 3292
rect 64216 3232 64280 3236
rect 64296 3292 64360 3296
rect 64296 3236 64300 3292
rect 64300 3236 64356 3292
rect 64356 3236 64360 3292
rect 64296 3232 64360 3236
rect 64376 3292 64440 3296
rect 64376 3236 64380 3292
rect 64380 3236 64436 3292
rect 64436 3236 64440 3292
rect 64376 3232 64440 3236
rect 64456 3292 64520 3296
rect 64456 3236 64460 3292
rect 64460 3236 64516 3292
rect 64516 3236 64520 3292
rect 64456 3232 64520 3236
rect 24216 3158 24280 3222
rect 24296 3158 24360 3222
rect 24376 3158 24440 3222
rect 24456 3158 24520 3222
rect 15700 3028 15764 3092
rect 24216 3078 24280 3142
rect 24296 3078 24360 3142
rect 24376 3078 24440 3142
rect 24456 3078 24520 3142
rect 24216 2998 24280 3062
rect 24296 2998 24360 3062
rect 24376 2998 24440 3062
rect 24456 2998 24520 3062
rect 40724 3088 40788 3092
rect 40724 3032 40738 3088
rect 40738 3032 40788 3088
rect 40724 3028 40788 3032
rect 41460 3088 41524 3092
rect 41460 3032 41474 3088
rect 41474 3032 41524 3088
rect 41460 3028 41524 3032
rect 42380 3028 42444 3092
rect 43852 3028 43916 3092
rect 9216 2748 9280 2752
rect 9216 2692 9220 2748
rect 9220 2692 9276 2748
rect 9276 2692 9280 2748
rect 9216 2688 9280 2692
rect 9296 2748 9360 2752
rect 9296 2692 9300 2748
rect 9300 2692 9356 2748
rect 9356 2692 9360 2748
rect 9296 2688 9360 2692
rect 9376 2748 9440 2752
rect 9376 2692 9380 2748
rect 9380 2692 9436 2748
rect 9436 2692 9440 2748
rect 9376 2688 9440 2692
rect 9456 2748 9520 2752
rect 9456 2692 9460 2748
rect 9460 2692 9516 2748
rect 9516 2692 9520 2748
rect 9456 2688 9520 2692
rect 13124 2680 13188 2684
rect 13124 2624 13138 2680
rect 13138 2624 13188 2680
rect 13124 2620 13188 2624
rect 13860 2680 13924 2684
rect 24216 2918 24280 2982
rect 24296 2918 24360 2982
rect 24376 2918 24440 2982
rect 24456 2918 24520 2982
rect 24216 2838 24280 2902
rect 24296 2838 24360 2902
rect 24376 2838 24440 2902
rect 24456 2838 24520 2902
rect 33916 2892 33980 2956
rect 44956 2756 45020 2820
rect 39216 2748 39280 2752
rect 39216 2692 39220 2748
rect 39220 2692 39276 2748
rect 39276 2692 39280 2748
rect 39216 2688 39280 2692
rect 39296 2748 39360 2752
rect 39296 2692 39300 2748
rect 39300 2692 39356 2748
rect 39356 2692 39360 2748
rect 39296 2688 39360 2692
rect 39376 2748 39440 2752
rect 39376 2692 39380 2748
rect 39380 2692 39436 2748
rect 39436 2692 39440 2748
rect 39376 2688 39440 2692
rect 39456 2748 39520 2752
rect 39456 2692 39460 2748
rect 39460 2692 39516 2748
rect 39516 2692 39520 2748
rect 39456 2688 39520 2692
rect 13860 2624 13874 2680
rect 13874 2624 13924 2680
rect 13860 2620 13924 2624
rect 42564 2620 42628 2684
rect 49216 2748 49280 2752
rect 49216 2692 49220 2748
rect 49220 2692 49276 2748
rect 49276 2692 49280 2748
rect 49216 2688 49280 2692
rect 49296 2748 49360 2752
rect 49296 2692 49300 2748
rect 49300 2692 49356 2748
rect 49356 2692 49360 2748
rect 49296 2688 49360 2692
rect 49376 2748 49440 2752
rect 49376 2692 49380 2748
rect 49380 2692 49436 2748
rect 49436 2692 49440 2748
rect 49376 2688 49440 2692
rect 49456 2748 49520 2752
rect 49456 2692 49460 2748
rect 49460 2692 49516 2748
rect 49516 2692 49520 2748
rect 49456 2688 49520 2692
rect 29216 2366 29280 2430
rect 29296 2366 29360 2430
rect 29376 2366 29440 2430
rect 29456 2366 29520 2430
rect 29216 2286 29280 2350
rect 29296 2286 29360 2350
rect 29376 2286 29440 2350
rect 29456 2286 29520 2350
rect 59216 2748 59280 2752
rect 59216 2692 59220 2748
rect 59220 2692 59276 2748
rect 59276 2692 59280 2748
rect 59216 2688 59280 2692
rect 59296 2748 59360 2752
rect 59296 2692 59300 2748
rect 59300 2692 59356 2748
rect 59356 2692 59360 2748
rect 59296 2688 59360 2692
rect 59376 2748 59440 2752
rect 59376 2692 59380 2748
rect 59380 2692 59436 2748
rect 59436 2692 59440 2748
rect 59376 2688 59440 2692
rect 59456 2748 59520 2752
rect 59456 2692 59460 2748
rect 59460 2692 59516 2748
rect 59516 2692 59520 2748
rect 59456 2688 59520 2692
rect 53604 2484 53668 2548
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 14216 2204 14280 2208
rect 14216 2148 14220 2204
rect 14220 2148 14276 2204
rect 14276 2148 14280 2204
rect 14216 2144 14280 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 29216 2206 29280 2270
rect 29296 2206 29360 2270
rect 29376 2206 29440 2270
rect 29456 2206 29520 2270
rect 42012 2212 42076 2276
rect 49740 2212 49804 2276
rect 44216 2204 44280 2208
rect 44216 2148 44220 2204
rect 44220 2148 44276 2204
rect 44276 2148 44280 2204
rect 44216 2144 44280 2148
rect 44296 2204 44360 2208
rect 44296 2148 44300 2204
rect 44300 2148 44356 2204
rect 44356 2148 44360 2204
rect 44296 2144 44360 2148
rect 44376 2204 44440 2208
rect 44376 2148 44380 2204
rect 44380 2148 44436 2204
rect 44436 2148 44440 2204
rect 44376 2144 44440 2148
rect 44456 2204 44520 2208
rect 44456 2148 44460 2204
rect 44460 2148 44516 2204
rect 44516 2148 44520 2204
rect 44456 2144 44520 2148
rect 54216 2204 54280 2208
rect 54216 2148 54220 2204
rect 54220 2148 54276 2204
rect 54276 2148 54280 2204
rect 54216 2144 54280 2148
rect 54296 2204 54360 2208
rect 54296 2148 54300 2204
rect 54300 2148 54356 2204
rect 54356 2148 54360 2204
rect 54296 2144 54360 2148
rect 54376 2204 54440 2208
rect 54376 2148 54380 2204
rect 54380 2148 54436 2204
rect 54436 2148 54440 2204
rect 54376 2144 54440 2148
rect 54456 2204 54520 2208
rect 54456 2148 54460 2204
rect 54460 2148 54516 2204
rect 54516 2148 54520 2204
rect 54456 2144 54520 2148
rect 64216 2204 64280 2208
rect 64216 2148 64220 2204
rect 64220 2148 64276 2204
rect 64276 2148 64280 2204
rect 64216 2144 64280 2148
rect 64296 2204 64360 2208
rect 64296 2148 64300 2204
rect 64300 2148 64356 2204
rect 64356 2148 64360 2204
rect 64296 2144 64360 2148
rect 64376 2204 64440 2208
rect 64376 2148 64380 2204
rect 64380 2148 64436 2204
rect 64436 2148 64440 2204
rect 64376 2144 64440 2148
rect 64456 2204 64520 2208
rect 64456 2148 64460 2204
rect 64460 2148 64516 2204
rect 64516 2148 64520 2204
rect 64456 2144 64520 2148
rect 5396 1940 5460 2004
rect 46612 1940 46676 2004
rect 54892 1940 54956 2004
rect 64644 1940 64708 2004
rect 27660 1864 27724 1868
rect 27660 1808 27710 1864
rect 27710 1808 27724 1864
rect 27660 1804 27724 1808
rect 28028 1864 28092 1868
rect 28028 1808 28078 1864
rect 28078 1808 28092 1864
rect 28028 1804 28092 1808
rect 30052 1804 30116 1868
rect 30420 1804 30484 1868
rect 31156 1804 31220 1868
rect 28212 1728 28276 1732
rect 28212 1672 28226 1728
rect 28226 1672 28276 1728
rect 28212 1668 28276 1672
rect 30604 1668 30668 1732
rect 41276 1260 41340 1324
rect 31892 1184 31956 1188
rect 31892 1128 31906 1184
rect 31906 1128 31956 1184
rect 31892 1124 31956 1128
<< metal4 >>
rect 4208 67488 4528 67504
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66400 4528 67424
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 9208 66944 9528 67504
rect 9208 66880 9216 66944
rect 9280 66880 9296 66944
rect 9360 66880 9376 66944
rect 9440 66880 9456 66944
rect 9520 66880 9528 66944
rect 9208 65856 9528 66880
rect 9208 65792 9216 65856
rect 9280 65792 9296 65856
rect 9360 65792 9376 65856
rect 9440 65792 9456 65856
rect 9520 65792 9528 65856
rect 9208 64768 9528 65792
rect 9208 64704 9216 64768
rect 9280 64704 9296 64768
rect 9360 64704 9376 64768
rect 9440 64704 9456 64768
rect 9520 64704 9528 64768
rect 9208 63680 9528 64704
rect 9208 63616 9216 63680
rect 9280 63616 9296 63680
rect 9360 63616 9376 63680
rect 9440 63616 9456 63680
rect 9520 63616 9528 63680
rect 9208 62592 9528 63616
rect 9208 62528 9216 62592
rect 9280 62528 9296 62592
rect 9360 62528 9376 62592
rect 9440 62528 9456 62592
rect 9520 62528 9528 62592
rect 9208 61504 9528 62528
rect 9208 61440 9216 61504
rect 9280 61440 9296 61504
rect 9360 61440 9376 61504
rect 9440 61440 9456 61504
rect 9520 61440 9528 61504
rect 9208 60416 9528 61440
rect 9208 60352 9216 60416
rect 9280 60352 9296 60416
rect 9360 60352 9376 60416
rect 9440 60352 9456 60416
rect 9520 60352 9528 60416
rect 9208 59328 9528 60352
rect 9208 59264 9216 59328
rect 9280 59264 9296 59328
rect 9360 59264 9376 59328
rect 9440 59264 9456 59328
rect 9520 59264 9528 59328
rect 9208 58240 9528 59264
rect 9208 58176 9216 58240
rect 9280 58176 9296 58240
rect 9360 58176 9376 58240
rect 9440 58176 9456 58240
rect 9520 58176 9528 58240
rect 9208 57152 9528 58176
rect 9208 57088 9216 57152
rect 9280 57088 9296 57152
rect 9360 57088 9376 57152
rect 9440 57088 9456 57152
rect 9520 57088 9528 57152
rect 9208 56064 9528 57088
rect 9208 56000 9216 56064
rect 9280 56000 9296 56064
rect 9360 56000 9376 56064
rect 9440 56000 9456 56064
rect 9520 56000 9528 56064
rect 9208 54976 9528 56000
rect 9208 54912 9216 54976
rect 9280 54912 9296 54976
rect 9360 54912 9376 54976
rect 9440 54912 9456 54976
rect 9520 54912 9528 54976
rect 9208 53888 9528 54912
rect 9208 53824 9216 53888
rect 9280 53824 9296 53888
rect 9360 53824 9376 53888
rect 9440 53824 9456 53888
rect 9520 53824 9528 53888
rect 9208 52800 9528 53824
rect 9208 52736 9216 52800
rect 9280 52736 9296 52800
rect 9360 52736 9376 52800
rect 9440 52736 9456 52800
rect 9520 52736 9528 52800
rect 9208 51712 9528 52736
rect 9208 51648 9216 51712
rect 9280 51648 9296 51712
rect 9360 51648 9376 51712
rect 9440 51648 9456 51712
rect 9520 51648 9528 51712
rect 9208 50624 9528 51648
rect 9208 50560 9216 50624
rect 9280 50560 9296 50624
rect 9360 50560 9376 50624
rect 9440 50560 9456 50624
rect 9520 50560 9528 50624
rect 9208 49536 9528 50560
rect 9208 49472 9216 49536
rect 9280 49472 9296 49536
rect 9360 49472 9376 49536
rect 9440 49472 9456 49536
rect 9520 49472 9528 49536
rect 9208 48448 9528 49472
rect 9208 48384 9216 48448
rect 9280 48384 9296 48448
rect 9360 48384 9376 48448
rect 9440 48384 9456 48448
rect 9520 48384 9528 48448
rect 9208 47360 9528 48384
rect 9208 47296 9216 47360
rect 9280 47296 9296 47360
rect 9360 47296 9376 47360
rect 9440 47296 9456 47360
rect 9520 47296 9528 47360
rect 9208 46272 9528 47296
rect 9208 46208 9216 46272
rect 9280 46208 9296 46272
rect 9360 46208 9376 46272
rect 9440 46208 9456 46272
rect 9520 46208 9528 46272
rect 9208 45184 9528 46208
rect 9208 45120 9216 45184
rect 9280 45120 9296 45184
rect 9360 45120 9376 45184
rect 9440 45120 9456 45184
rect 9520 45120 9528 45184
rect 9208 44096 9528 45120
rect 9208 44032 9216 44096
rect 9280 44032 9296 44096
rect 9360 44032 9376 44096
rect 9440 44032 9456 44096
rect 9520 44032 9528 44096
rect 9208 43008 9528 44032
rect 9208 42944 9216 43008
rect 9280 42944 9296 43008
rect 9360 42944 9376 43008
rect 9440 42944 9456 43008
rect 9520 42944 9528 43008
rect 9208 41920 9528 42944
rect 9208 41856 9216 41920
rect 9280 41856 9296 41920
rect 9360 41856 9376 41920
rect 9440 41856 9456 41920
rect 9520 41856 9528 41920
rect 9208 40832 9528 41856
rect 9208 40768 9216 40832
rect 9280 40768 9296 40832
rect 9360 40768 9376 40832
rect 9440 40768 9456 40832
rect 9520 40768 9528 40832
rect 9208 39744 9528 40768
rect 9208 39680 9216 39744
rect 9280 39680 9296 39744
rect 9360 39680 9376 39744
rect 9440 39680 9456 39744
rect 9520 39680 9528 39744
rect 9208 38656 9528 39680
rect 9208 38592 9216 38656
rect 9280 38592 9296 38656
rect 9360 38592 9376 38656
rect 9440 38592 9456 38656
rect 9520 38592 9528 38656
rect 9208 37568 9528 38592
rect 9208 37504 9216 37568
rect 9280 37504 9296 37568
rect 9360 37504 9376 37568
rect 9440 37504 9456 37568
rect 9520 37504 9528 37568
rect 9208 36480 9528 37504
rect 9208 36416 9216 36480
rect 9280 36416 9296 36480
rect 9360 36416 9376 36480
rect 9440 36416 9456 36480
rect 9520 36416 9528 36480
rect 9208 35392 9528 36416
rect 9208 35328 9216 35392
rect 9280 35328 9296 35392
rect 9360 35328 9376 35392
rect 9440 35328 9456 35392
rect 9520 35328 9528 35392
rect 9208 34304 9528 35328
rect 9208 34240 9216 34304
rect 9280 34240 9296 34304
rect 9360 34240 9376 34304
rect 9440 34240 9456 34304
rect 9520 34240 9528 34304
rect 9208 33216 9528 34240
rect 9208 33152 9216 33216
rect 9280 33152 9296 33216
rect 9360 33152 9376 33216
rect 9440 33152 9456 33216
rect 9520 33152 9528 33216
rect 9208 32128 9528 33152
rect 9208 32064 9216 32128
rect 9280 32064 9296 32128
rect 9360 32064 9376 32128
rect 9440 32064 9456 32128
rect 9520 32064 9528 32128
rect 9208 31040 9528 32064
rect 9208 30976 9216 31040
rect 9280 30976 9296 31040
rect 9360 30976 9376 31040
rect 9440 30976 9456 31040
rect 9520 30976 9528 31040
rect 9208 29952 9528 30976
rect 9208 29888 9216 29952
rect 9280 29888 9296 29952
rect 9360 29888 9376 29952
rect 9440 29888 9456 29952
rect 9520 29888 9528 29952
rect 9208 28864 9528 29888
rect 9208 28800 9216 28864
rect 9280 28800 9296 28864
rect 9360 28800 9376 28864
rect 9440 28800 9456 28864
rect 9520 28800 9528 28864
rect 9208 27776 9528 28800
rect 9208 27712 9216 27776
rect 9280 27712 9296 27776
rect 9360 27712 9376 27776
rect 9440 27712 9456 27776
rect 9520 27712 9528 27776
rect 9208 26688 9528 27712
rect 9208 26624 9216 26688
rect 9280 26624 9296 26688
rect 9360 26624 9376 26688
rect 9440 26624 9456 26688
rect 9520 26624 9528 26688
rect 9208 25600 9528 26624
rect 9208 25536 9216 25600
rect 9280 25536 9296 25600
rect 9360 25536 9376 25600
rect 9440 25536 9456 25600
rect 9520 25536 9528 25600
rect 9208 24512 9528 25536
rect 9208 24448 9216 24512
rect 9280 24448 9296 24512
rect 9360 24448 9376 24512
rect 9440 24448 9456 24512
rect 9520 24448 9528 24512
rect 9208 23424 9528 24448
rect 9208 23360 9216 23424
rect 9280 23360 9296 23424
rect 9360 23360 9376 23424
rect 9440 23360 9456 23424
rect 9520 23360 9528 23424
rect 9208 22336 9528 23360
rect 9208 22272 9216 22336
rect 9280 22272 9296 22336
rect 9360 22272 9376 22336
rect 9440 22272 9456 22336
rect 9520 22272 9528 22336
rect 9208 21248 9528 22272
rect 9208 21184 9216 21248
rect 9280 21184 9296 21248
rect 9360 21184 9376 21248
rect 9440 21184 9456 21248
rect 9520 21184 9528 21248
rect 9208 20160 9528 21184
rect 9208 20096 9216 20160
rect 9280 20096 9296 20160
rect 9360 20096 9376 20160
rect 9440 20096 9456 20160
rect 9520 20096 9528 20160
rect 9208 19072 9528 20096
rect 9208 19008 9216 19072
rect 9280 19008 9296 19072
rect 9360 19008 9376 19072
rect 9440 19008 9456 19072
rect 9520 19008 9528 19072
rect 9208 17984 9528 19008
rect 9208 17920 9216 17984
rect 9280 17920 9296 17984
rect 9360 17920 9376 17984
rect 9440 17920 9456 17984
rect 9520 17920 9528 17984
rect 9208 16896 9528 17920
rect 9208 16832 9216 16896
rect 9280 16832 9296 16896
rect 9360 16832 9376 16896
rect 9440 16832 9456 16896
rect 9520 16832 9528 16896
rect 9208 15808 9528 16832
rect 9208 15744 9216 15808
rect 9280 15744 9296 15808
rect 9360 15744 9376 15808
rect 9440 15744 9456 15808
rect 9520 15744 9528 15808
rect 9208 14720 9528 15744
rect 9208 14656 9216 14720
rect 9280 14656 9296 14720
rect 9360 14656 9376 14720
rect 9440 14656 9456 14720
rect 9520 14656 9528 14720
rect 9208 13632 9528 14656
rect 9208 13568 9216 13632
rect 9280 13568 9296 13632
rect 9360 13568 9376 13632
rect 9440 13568 9456 13632
rect 9520 13568 9528 13632
rect 9208 12544 9528 13568
rect 14208 67488 14528 67504
rect 14208 67424 14216 67488
rect 14280 67424 14296 67488
rect 14360 67424 14376 67488
rect 14440 67424 14456 67488
rect 14520 67424 14528 67488
rect 14208 66400 14528 67424
rect 14208 66336 14216 66400
rect 14280 66336 14296 66400
rect 14360 66336 14376 66400
rect 14440 66336 14456 66400
rect 14520 66336 14528 66400
rect 14208 65312 14528 66336
rect 14208 65248 14216 65312
rect 14280 65248 14296 65312
rect 14360 65248 14376 65312
rect 14440 65248 14456 65312
rect 14520 65248 14528 65312
rect 14208 64224 14528 65248
rect 14208 64160 14216 64224
rect 14280 64160 14296 64224
rect 14360 64160 14376 64224
rect 14440 64160 14456 64224
rect 14520 64160 14528 64224
rect 14208 63136 14528 64160
rect 14208 63072 14216 63136
rect 14280 63072 14296 63136
rect 14360 63072 14376 63136
rect 14440 63072 14456 63136
rect 14520 63072 14528 63136
rect 14208 62048 14528 63072
rect 14208 61984 14216 62048
rect 14280 61984 14296 62048
rect 14360 61984 14376 62048
rect 14440 61984 14456 62048
rect 14520 61984 14528 62048
rect 14208 60960 14528 61984
rect 14208 60896 14216 60960
rect 14280 60896 14296 60960
rect 14360 60896 14376 60960
rect 14440 60896 14456 60960
rect 14520 60896 14528 60960
rect 14208 59872 14528 60896
rect 14208 59808 14216 59872
rect 14280 59808 14296 59872
rect 14360 59808 14376 59872
rect 14440 59808 14456 59872
rect 14520 59808 14528 59872
rect 14208 58784 14528 59808
rect 14208 58720 14216 58784
rect 14280 58720 14296 58784
rect 14360 58720 14376 58784
rect 14440 58720 14456 58784
rect 14520 58720 14528 58784
rect 14208 57696 14528 58720
rect 14208 57632 14216 57696
rect 14280 57632 14296 57696
rect 14360 57632 14376 57696
rect 14440 57632 14456 57696
rect 14520 57632 14528 57696
rect 14208 56608 14528 57632
rect 14208 56544 14216 56608
rect 14280 56544 14296 56608
rect 14360 56544 14376 56608
rect 14440 56544 14456 56608
rect 14520 56544 14528 56608
rect 14208 55520 14528 56544
rect 14208 55456 14216 55520
rect 14280 55456 14296 55520
rect 14360 55456 14376 55520
rect 14440 55456 14456 55520
rect 14520 55456 14528 55520
rect 14208 54432 14528 55456
rect 14208 54368 14216 54432
rect 14280 54368 14296 54432
rect 14360 54368 14376 54432
rect 14440 54368 14456 54432
rect 14520 54368 14528 54432
rect 14208 53344 14528 54368
rect 14208 53280 14216 53344
rect 14280 53280 14296 53344
rect 14360 53280 14376 53344
rect 14440 53280 14456 53344
rect 14520 53280 14528 53344
rect 14208 52256 14528 53280
rect 14208 52192 14216 52256
rect 14280 52192 14296 52256
rect 14360 52192 14376 52256
rect 14440 52192 14456 52256
rect 14520 52192 14528 52256
rect 14208 51168 14528 52192
rect 14208 51104 14216 51168
rect 14280 51104 14296 51168
rect 14360 51104 14376 51168
rect 14440 51104 14456 51168
rect 14520 51104 14528 51168
rect 14208 50080 14528 51104
rect 14208 50016 14216 50080
rect 14280 50016 14296 50080
rect 14360 50016 14376 50080
rect 14440 50016 14456 50080
rect 14520 50016 14528 50080
rect 14208 48992 14528 50016
rect 14208 48928 14216 48992
rect 14280 48928 14296 48992
rect 14360 48928 14376 48992
rect 14440 48928 14456 48992
rect 14520 48928 14528 48992
rect 14208 47904 14528 48928
rect 14208 47840 14216 47904
rect 14280 47840 14296 47904
rect 14360 47840 14376 47904
rect 14440 47840 14456 47904
rect 14520 47840 14528 47904
rect 14208 46816 14528 47840
rect 14208 46752 14216 46816
rect 14280 46752 14296 46816
rect 14360 46752 14376 46816
rect 14440 46752 14456 46816
rect 14520 46752 14528 46816
rect 14208 45728 14528 46752
rect 14208 45664 14216 45728
rect 14280 45664 14296 45728
rect 14360 45664 14376 45728
rect 14440 45664 14456 45728
rect 14520 45664 14528 45728
rect 14208 44640 14528 45664
rect 14208 44576 14216 44640
rect 14280 44576 14296 44640
rect 14360 44576 14376 44640
rect 14440 44576 14456 44640
rect 14520 44576 14528 44640
rect 14208 43552 14528 44576
rect 14208 43488 14216 43552
rect 14280 43488 14296 43552
rect 14360 43488 14376 43552
rect 14440 43488 14456 43552
rect 14520 43488 14528 43552
rect 14208 42464 14528 43488
rect 14208 42400 14216 42464
rect 14280 42400 14296 42464
rect 14360 42400 14376 42464
rect 14440 42400 14456 42464
rect 14520 42400 14528 42464
rect 14208 41376 14528 42400
rect 14208 41312 14216 41376
rect 14280 41312 14296 41376
rect 14360 41312 14376 41376
rect 14440 41312 14456 41376
rect 14520 41312 14528 41376
rect 14208 40288 14528 41312
rect 14208 40224 14216 40288
rect 14280 40224 14296 40288
rect 14360 40224 14376 40288
rect 14440 40224 14456 40288
rect 14520 40224 14528 40288
rect 14208 39200 14528 40224
rect 14208 39136 14216 39200
rect 14280 39136 14296 39200
rect 14360 39136 14376 39200
rect 14440 39136 14456 39200
rect 14520 39136 14528 39200
rect 14208 38112 14528 39136
rect 14208 38048 14216 38112
rect 14280 38048 14296 38112
rect 14360 38048 14376 38112
rect 14440 38048 14456 38112
rect 14520 38048 14528 38112
rect 14208 37024 14528 38048
rect 14208 36960 14216 37024
rect 14280 36960 14296 37024
rect 14360 36960 14376 37024
rect 14440 36960 14456 37024
rect 14520 36960 14528 37024
rect 14208 35936 14528 36960
rect 14208 35872 14216 35936
rect 14280 35872 14296 35936
rect 14360 35872 14376 35936
rect 14440 35872 14456 35936
rect 14520 35872 14528 35936
rect 14208 34848 14528 35872
rect 14208 34784 14216 34848
rect 14280 34784 14296 34848
rect 14360 34784 14376 34848
rect 14440 34784 14456 34848
rect 14520 34784 14528 34848
rect 14208 33760 14528 34784
rect 14208 33696 14216 33760
rect 14280 33696 14296 33760
rect 14360 33696 14376 33760
rect 14440 33696 14456 33760
rect 14520 33696 14528 33760
rect 14208 32672 14528 33696
rect 14208 32608 14216 32672
rect 14280 32608 14296 32672
rect 14360 32608 14376 32672
rect 14440 32608 14456 32672
rect 14520 32608 14528 32672
rect 14208 31584 14528 32608
rect 14208 31520 14216 31584
rect 14280 31520 14296 31584
rect 14360 31520 14376 31584
rect 14440 31520 14456 31584
rect 14520 31520 14528 31584
rect 14208 30496 14528 31520
rect 14208 30432 14216 30496
rect 14280 30432 14296 30496
rect 14360 30432 14376 30496
rect 14440 30432 14456 30496
rect 14520 30432 14528 30496
rect 14208 29408 14528 30432
rect 14208 29344 14216 29408
rect 14280 29344 14296 29408
rect 14360 29344 14376 29408
rect 14440 29344 14456 29408
rect 14520 29344 14528 29408
rect 14208 28320 14528 29344
rect 14208 28256 14216 28320
rect 14280 28256 14296 28320
rect 14360 28256 14376 28320
rect 14440 28256 14456 28320
rect 14520 28256 14528 28320
rect 14208 27232 14528 28256
rect 14208 27168 14216 27232
rect 14280 27168 14296 27232
rect 14360 27168 14376 27232
rect 14440 27168 14456 27232
rect 14520 27168 14528 27232
rect 14208 26144 14528 27168
rect 14208 26080 14216 26144
rect 14280 26080 14296 26144
rect 14360 26080 14376 26144
rect 14440 26080 14456 26144
rect 14520 26080 14528 26144
rect 14208 25056 14528 26080
rect 14208 24992 14216 25056
rect 14280 24992 14296 25056
rect 14360 24992 14376 25056
rect 14440 24992 14456 25056
rect 14520 24992 14528 25056
rect 14208 23968 14528 24992
rect 14208 23904 14216 23968
rect 14280 23904 14296 23968
rect 14360 23904 14376 23968
rect 14440 23904 14456 23968
rect 14520 23904 14528 23968
rect 14208 22880 14528 23904
rect 14208 22816 14216 22880
rect 14280 22816 14296 22880
rect 14360 22816 14376 22880
rect 14440 22816 14456 22880
rect 14520 22816 14528 22880
rect 14208 21792 14528 22816
rect 14208 21728 14216 21792
rect 14280 21728 14296 21792
rect 14360 21728 14376 21792
rect 14440 21728 14456 21792
rect 14520 21728 14528 21792
rect 14208 20704 14528 21728
rect 14208 20640 14216 20704
rect 14280 20640 14296 20704
rect 14360 20640 14376 20704
rect 14440 20640 14456 20704
rect 14520 20640 14528 20704
rect 14208 19616 14528 20640
rect 14208 19552 14216 19616
rect 14280 19552 14296 19616
rect 14360 19552 14376 19616
rect 14440 19552 14456 19616
rect 14520 19552 14528 19616
rect 14208 18528 14528 19552
rect 14208 18464 14216 18528
rect 14280 18464 14296 18528
rect 14360 18464 14376 18528
rect 14440 18464 14456 18528
rect 14520 18464 14528 18528
rect 14208 17440 14528 18464
rect 14208 17376 14216 17440
rect 14280 17376 14296 17440
rect 14360 17376 14376 17440
rect 14440 17376 14456 17440
rect 14520 17376 14528 17440
rect 14208 16352 14528 17376
rect 14208 16288 14216 16352
rect 14280 16288 14296 16352
rect 14360 16288 14376 16352
rect 14440 16288 14456 16352
rect 14520 16288 14528 16352
rect 14208 15264 14528 16288
rect 14208 15200 14216 15264
rect 14280 15200 14296 15264
rect 14360 15200 14376 15264
rect 14440 15200 14456 15264
rect 14520 15200 14528 15264
rect 14208 14176 14528 15200
rect 14208 14112 14216 14176
rect 14280 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14528 14176
rect 13491 13156 13557 13157
rect 13491 13092 13492 13156
rect 13556 13092 13557 13156
rect 13491 13091 13557 13092
rect 13123 12612 13189 12613
rect 13123 12548 13124 12612
rect 13188 12548 13189 12612
rect 13123 12547 13189 12548
rect 9208 12480 9216 12544
rect 9280 12480 9296 12544
rect 9360 12480 9376 12544
rect 9440 12480 9456 12544
rect 9520 12480 9528 12544
rect 9208 11456 9528 12480
rect 9208 11392 9216 11456
rect 9280 11392 9296 11456
rect 9360 11392 9376 11456
rect 9440 11392 9456 11456
rect 9520 11392 9528 11456
rect 9208 10368 9528 11392
rect 9627 11252 9693 11253
rect 9627 11188 9628 11252
rect 9692 11188 9693 11252
rect 9627 11187 9693 11188
rect 9208 10304 9216 10368
rect 9280 10304 9296 10368
rect 9360 10304 9376 10368
rect 9440 10304 9456 10368
rect 9520 10304 9528 10368
rect 9208 9280 9528 10304
rect 9208 9216 9216 9280
rect 9280 9216 9296 9280
rect 9360 9216 9376 9280
rect 9440 9216 9456 9280
rect 9520 9216 9528 9280
rect 9208 8192 9528 9216
rect 9208 8128 9216 8192
rect 9280 8128 9296 8192
rect 9360 8128 9376 8192
rect 9440 8128 9456 8192
rect 9520 8128 9528 8192
rect 5395 7172 5461 7173
rect 5395 7108 5396 7172
rect 5460 7108 5461 7172
rect 5395 7107 5461 7108
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 5398 5133 5458 7107
rect 9208 7104 9528 8128
rect 9208 7040 9216 7104
rect 9280 7040 9296 7104
rect 9360 7040 9376 7104
rect 9440 7040 9456 7104
rect 9520 7040 9528 7104
rect 9208 6016 9528 7040
rect 9208 5952 9216 6016
rect 9280 5952 9296 6016
rect 9360 5952 9376 6016
rect 9440 5952 9456 6016
rect 9520 5952 9528 6016
rect 5395 5132 5461 5133
rect 5395 5068 5396 5132
rect 5460 5068 5461 5132
rect 5395 5067 5461 5068
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 5398 2005 5458 5067
rect 9208 4928 9528 5952
rect 9208 4864 9216 4928
rect 9280 4864 9296 4928
rect 9360 4864 9376 4928
rect 9440 4864 9456 4928
rect 9520 4864 9528 4928
rect 9208 3840 9528 4864
rect 9208 3776 9216 3840
rect 9280 3776 9296 3840
rect 9360 3776 9376 3840
rect 9440 3776 9456 3840
rect 9520 3776 9528 3840
rect 9208 2752 9528 3776
rect 9630 3773 9690 11187
rect 11651 10028 11717 10029
rect 11651 9964 11652 10028
rect 11716 9964 11717 10028
rect 11651 9963 11717 9964
rect 11654 4045 11714 9963
rect 12203 8532 12269 8533
rect 12203 8468 12204 8532
rect 12268 8468 12269 8532
rect 12203 8467 12269 8468
rect 11651 4044 11717 4045
rect 11651 3980 11652 4044
rect 11716 3980 11717 4044
rect 11651 3979 11717 3980
rect 12206 3773 12266 8467
rect 9627 3772 9693 3773
rect 9627 3708 9628 3772
rect 9692 3708 9693 3772
rect 9627 3707 9693 3708
rect 12203 3772 12269 3773
rect 12203 3708 12204 3772
rect 12268 3708 12269 3772
rect 12203 3707 12269 3708
rect 9208 2688 9216 2752
rect 9280 2688 9296 2752
rect 9360 2688 9376 2752
rect 9440 2688 9456 2752
rect 9520 2688 9528 2752
rect 9208 2128 9528 2688
rect 13126 2685 13186 12547
rect 13494 3773 13554 13091
rect 14208 13088 14528 14112
rect 19208 66944 19528 67504
rect 19208 66880 19216 66944
rect 19280 66880 19296 66944
rect 19360 66880 19376 66944
rect 19440 66880 19456 66944
rect 19520 66880 19528 66944
rect 19208 65856 19528 66880
rect 19208 65792 19216 65856
rect 19280 65792 19296 65856
rect 19360 65792 19376 65856
rect 19440 65792 19456 65856
rect 19520 65792 19528 65856
rect 19208 64768 19528 65792
rect 19208 64704 19216 64768
rect 19280 64704 19296 64768
rect 19360 64704 19376 64768
rect 19440 64704 19456 64768
rect 19520 64704 19528 64768
rect 19208 63680 19528 64704
rect 19208 63616 19216 63680
rect 19280 63616 19296 63680
rect 19360 63616 19376 63680
rect 19440 63616 19456 63680
rect 19520 63616 19528 63680
rect 19208 62592 19528 63616
rect 19208 62528 19216 62592
rect 19280 62528 19296 62592
rect 19360 62528 19376 62592
rect 19440 62528 19456 62592
rect 19520 62528 19528 62592
rect 19208 61504 19528 62528
rect 19208 61440 19216 61504
rect 19280 61440 19296 61504
rect 19360 61440 19376 61504
rect 19440 61440 19456 61504
rect 19520 61440 19528 61504
rect 19208 60416 19528 61440
rect 19208 60352 19216 60416
rect 19280 60352 19296 60416
rect 19360 60352 19376 60416
rect 19440 60352 19456 60416
rect 19520 60352 19528 60416
rect 19208 59328 19528 60352
rect 19208 59264 19216 59328
rect 19280 59264 19296 59328
rect 19360 59264 19376 59328
rect 19440 59264 19456 59328
rect 19520 59264 19528 59328
rect 19208 58240 19528 59264
rect 19208 58176 19216 58240
rect 19280 58176 19296 58240
rect 19360 58176 19376 58240
rect 19440 58176 19456 58240
rect 19520 58176 19528 58240
rect 19208 57152 19528 58176
rect 19208 57088 19216 57152
rect 19280 57088 19296 57152
rect 19360 57088 19376 57152
rect 19440 57088 19456 57152
rect 19520 57088 19528 57152
rect 19208 56064 19528 57088
rect 19208 56000 19216 56064
rect 19280 56000 19296 56064
rect 19360 56000 19376 56064
rect 19440 56000 19456 56064
rect 19520 56000 19528 56064
rect 19208 54976 19528 56000
rect 19208 54912 19216 54976
rect 19280 54912 19296 54976
rect 19360 54912 19376 54976
rect 19440 54912 19456 54976
rect 19520 54912 19528 54976
rect 19208 53888 19528 54912
rect 19208 53824 19216 53888
rect 19280 53824 19296 53888
rect 19360 53824 19376 53888
rect 19440 53824 19456 53888
rect 19520 53824 19528 53888
rect 19208 52800 19528 53824
rect 19208 52736 19216 52800
rect 19280 52736 19296 52800
rect 19360 52736 19376 52800
rect 19440 52736 19456 52800
rect 19520 52736 19528 52800
rect 19208 51712 19528 52736
rect 19208 51648 19216 51712
rect 19280 51648 19296 51712
rect 19360 51648 19376 51712
rect 19440 51648 19456 51712
rect 19520 51648 19528 51712
rect 19208 50624 19528 51648
rect 19208 50560 19216 50624
rect 19280 50560 19296 50624
rect 19360 50560 19376 50624
rect 19440 50560 19456 50624
rect 19520 50560 19528 50624
rect 19208 49536 19528 50560
rect 19208 49472 19216 49536
rect 19280 49472 19296 49536
rect 19360 49472 19376 49536
rect 19440 49472 19456 49536
rect 19520 49472 19528 49536
rect 19208 48448 19528 49472
rect 19208 48384 19216 48448
rect 19280 48384 19296 48448
rect 19360 48384 19376 48448
rect 19440 48384 19456 48448
rect 19520 48384 19528 48448
rect 19208 47360 19528 48384
rect 19208 47296 19216 47360
rect 19280 47296 19296 47360
rect 19360 47296 19376 47360
rect 19440 47296 19456 47360
rect 19520 47296 19528 47360
rect 19208 46272 19528 47296
rect 19208 46208 19216 46272
rect 19280 46208 19296 46272
rect 19360 46208 19376 46272
rect 19440 46208 19456 46272
rect 19520 46208 19528 46272
rect 19208 45184 19528 46208
rect 19208 45120 19216 45184
rect 19280 45120 19296 45184
rect 19360 45120 19376 45184
rect 19440 45120 19456 45184
rect 19520 45120 19528 45184
rect 19208 44096 19528 45120
rect 19208 44032 19216 44096
rect 19280 44032 19296 44096
rect 19360 44032 19376 44096
rect 19440 44032 19456 44096
rect 19520 44032 19528 44096
rect 19208 43008 19528 44032
rect 19208 42944 19216 43008
rect 19280 42944 19296 43008
rect 19360 42944 19376 43008
rect 19440 42944 19456 43008
rect 19520 42944 19528 43008
rect 19208 41920 19528 42944
rect 19208 41856 19216 41920
rect 19280 41856 19296 41920
rect 19360 41856 19376 41920
rect 19440 41856 19456 41920
rect 19520 41856 19528 41920
rect 19208 40832 19528 41856
rect 19208 40768 19216 40832
rect 19280 40768 19296 40832
rect 19360 40768 19376 40832
rect 19440 40768 19456 40832
rect 19520 40768 19528 40832
rect 19208 39744 19528 40768
rect 19208 39680 19216 39744
rect 19280 39680 19296 39744
rect 19360 39680 19376 39744
rect 19440 39680 19456 39744
rect 19520 39680 19528 39744
rect 19208 38656 19528 39680
rect 19208 38592 19216 38656
rect 19280 38592 19296 38656
rect 19360 38592 19376 38656
rect 19440 38592 19456 38656
rect 19520 38592 19528 38656
rect 19208 37568 19528 38592
rect 19208 37504 19216 37568
rect 19280 37504 19296 37568
rect 19360 37504 19376 37568
rect 19440 37504 19456 37568
rect 19520 37504 19528 37568
rect 19208 36480 19528 37504
rect 19208 36416 19216 36480
rect 19280 36416 19296 36480
rect 19360 36416 19376 36480
rect 19440 36416 19456 36480
rect 19520 36416 19528 36480
rect 19208 35392 19528 36416
rect 19208 35328 19216 35392
rect 19280 35328 19296 35392
rect 19360 35328 19376 35392
rect 19440 35328 19456 35392
rect 19520 35328 19528 35392
rect 19208 34304 19528 35328
rect 19208 34240 19216 34304
rect 19280 34240 19296 34304
rect 19360 34240 19376 34304
rect 19440 34240 19456 34304
rect 19520 34240 19528 34304
rect 19208 33216 19528 34240
rect 19208 33152 19216 33216
rect 19280 33152 19296 33216
rect 19360 33152 19376 33216
rect 19440 33152 19456 33216
rect 19520 33152 19528 33216
rect 19208 32128 19528 33152
rect 19208 32064 19216 32128
rect 19280 32064 19296 32128
rect 19360 32064 19376 32128
rect 19440 32064 19456 32128
rect 19520 32064 19528 32128
rect 19208 31040 19528 32064
rect 19208 30976 19216 31040
rect 19280 30976 19296 31040
rect 19360 30976 19376 31040
rect 19440 30976 19456 31040
rect 19520 30976 19528 31040
rect 19208 29952 19528 30976
rect 19208 29888 19216 29952
rect 19280 29888 19296 29952
rect 19360 29888 19376 29952
rect 19440 29888 19456 29952
rect 19520 29888 19528 29952
rect 19208 28864 19528 29888
rect 19208 28800 19216 28864
rect 19280 28800 19296 28864
rect 19360 28800 19376 28864
rect 19440 28800 19456 28864
rect 19520 28800 19528 28864
rect 19208 27776 19528 28800
rect 19208 27712 19216 27776
rect 19280 27712 19296 27776
rect 19360 27712 19376 27776
rect 19440 27712 19456 27776
rect 19520 27712 19528 27776
rect 19208 26688 19528 27712
rect 19208 26624 19216 26688
rect 19280 26624 19296 26688
rect 19360 26624 19376 26688
rect 19440 26624 19456 26688
rect 19520 26624 19528 26688
rect 19208 25600 19528 26624
rect 19208 25536 19216 25600
rect 19280 25536 19296 25600
rect 19360 25536 19376 25600
rect 19440 25536 19456 25600
rect 19520 25536 19528 25600
rect 19208 24512 19528 25536
rect 19208 24448 19216 24512
rect 19280 24448 19296 24512
rect 19360 24448 19376 24512
rect 19440 24448 19456 24512
rect 19520 24448 19528 24512
rect 19208 23424 19528 24448
rect 19208 23360 19216 23424
rect 19280 23360 19296 23424
rect 19360 23360 19376 23424
rect 19440 23360 19456 23424
rect 19520 23360 19528 23424
rect 19208 22336 19528 23360
rect 19208 22272 19216 22336
rect 19280 22272 19296 22336
rect 19360 22272 19376 22336
rect 19440 22272 19456 22336
rect 19520 22272 19528 22336
rect 19208 21248 19528 22272
rect 19208 21184 19216 21248
rect 19280 21184 19296 21248
rect 19360 21184 19376 21248
rect 19440 21184 19456 21248
rect 19520 21184 19528 21248
rect 19208 20160 19528 21184
rect 19208 20096 19216 20160
rect 19280 20096 19296 20160
rect 19360 20096 19376 20160
rect 19440 20096 19456 20160
rect 19520 20096 19528 20160
rect 15699 13836 15765 13837
rect 15699 13772 15700 13836
rect 15764 13772 15765 13836
rect 15699 13771 15765 13772
rect 16251 13836 16317 13837
rect 16251 13772 16252 13836
rect 16316 13772 16317 13836
rect 16251 13771 16317 13772
rect 14208 13024 14216 13088
rect 14280 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14528 13088
rect 14208 12000 14528 13024
rect 14208 11936 14216 12000
rect 14280 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14528 12000
rect 13859 11388 13925 11389
rect 13859 11324 13860 11388
rect 13924 11324 13925 11388
rect 13859 11323 13925 11324
rect 13675 7716 13741 7717
rect 13675 7652 13676 7716
rect 13740 7652 13741 7716
rect 13675 7651 13741 7652
rect 13678 4045 13738 7651
rect 13675 4044 13741 4045
rect 13675 3980 13676 4044
rect 13740 3980 13741 4044
rect 13675 3979 13741 3980
rect 13491 3772 13557 3773
rect 13491 3708 13492 3772
rect 13556 3708 13557 3772
rect 13491 3707 13557 3708
rect 13862 2685 13922 11323
rect 14208 10912 14528 11936
rect 14779 11660 14845 11661
rect 14779 11596 14780 11660
rect 14844 11596 14845 11660
rect 14779 11595 14845 11596
rect 14208 10848 14216 10912
rect 14280 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14528 10912
rect 14208 9824 14528 10848
rect 14782 10573 14842 11595
rect 14779 10572 14845 10573
rect 14779 10508 14780 10572
rect 14844 10508 14845 10572
rect 14779 10507 14845 10508
rect 14208 9760 14216 9824
rect 14280 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14528 9824
rect 14043 9076 14109 9077
rect 14043 9012 14044 9076
rect 14108 9012 14109 9076
rect 14043 9011 14109 9012
rect 14046 3909 14106 9011
rect 14208 8736 14528 9760
rect 14782 9349 14842 10507
rect 14779 9348 14845 9349
rect 14779 9284 14780 9348
rect 14844 9284 14845 9348
rect 14779 9283 14845 9284
rect 14595 8940 14661 8941
rect 14595 8876 14596 8940
rect 14660 8876 14661 8940
rect 14595 8875 14661 8876
rect 14208 8672 14216 8736
rect 14280 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14528 8736
rect 14208 7648 14528 8672
rect 14208 7584 14216 7648
rect 14280 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14528 7648
rect 14208 6560 14528 7584
rect 14208 6496 14216 6560
rect 14280 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14528 6560
rect 14208 5472 14528 6496
rect 14598 6357 14658 8875
rect 14595 6356 14661 6357
rect 14595 6292 14596 6356
rect 14660 6292 14661 6356
rect 14595 6291 14661 6292
rect 14208 5408 14216 5472
rect 14280 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14528 5472
rect 14208 4384 14528 5408
rect 14208 4320 14216 4384
rect 14280 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14528 4384
rect 14043 3908 14109 3909
rect 14043 3844 14044 3908
rect 14108 3844 14109 3908
rect 14043 3843 14109 3844
rect 14208 3296 14528 4320
rect 14208 3232 14216 3296
rect 14280 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14528 3296
rect 13123 2684 13189 2685
rect 13123 2620 13124 2684
rect 13188 2620 13189 2684
rect 13123 2619 13189 2620
rect 13859 2684 13925 2685
rect 13859 2620 13860 2684
rect 13924 2620 13925 2684
rect 13859 2619 13925 2620
rect 14208 2208 14528 3232
rect 15702 3093 15762 13771
rect 16254 4045 16314 13771
rect 16251 4044 16317 4045
rect 16251 3980 16252 4044
rect 16316 3980 16317 4044
rect 16251 3979 16317 3980
rect 15699 3092 15765 3093
rect 15699 3028 15700 3092
rect 15764 3028 15765 3092
rect 15699 3027 15765 3028
rect 14208 2144 14216 2208
rect 14280 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14528 2208
rect 19208 2176 19528 20096
rect 24208 67488 24528 67504
rect 24208 67424 24216 67488
rect 24280 67424 24296 67488
rect 24360 67424 24376 67488
rect 24440 67424 24456 67488
rect 24520 67424 24528 67488
rect 24208 66400 24528 67424
rect 24208 66336 24216 66400
rect 24280 66336 24296 66400
rect 24360 66336 24376 66400
rect 24440 66336 24456 66400
rect 24520 66336 24528 66400
rect 24208 65312 24528 66336
rect 24208 65248 24216 65312
rect 24280 65248 24296 65312
rect 24360 65248 24376 65312
rect 24440 65248 24456 65312
rect 24520 65248 24528 65312
rect 24208 64224 24528 65248
rect 24208 64160 24216 64224
rect 24280 64160 24296 64224
rect 24360 64160 24376 64224
rect 24440 64160 24456 64224
rect 24520 64160 24528 64224
rect 24208 63136 24528 64160
rect 24208 63072 24216 63136
rect 24280 63072 24296 63136
rect 24360 63072 24376 63136
rect 24440 63072 24456 63136
rect 24520 63072 24528 63136
rect 24208 62048 24528 63072
rect 24208 61984 24216 62048
rect 24280 61984 24296 62048
rect 24360 61984 24376 62048
rect 24440 61984 24456 62048
rect 24520 61984 24528 62048
rect 24208 60960 24528 61984
rect 24208 60896 24216 60960
rect 24280 60896 24296 60960
rect 24360 60896 24376 60960
rect 24440 60896 24456 60960
rect 24520 60896 24528 60960
rect 24208 59872 24528 60896
rect 24208 59808 24216 59872
rect 24280 59808 24296 59872
rect 24360 59808 24376 59872
rect 24440 59808 24456 59872
rect 24520 59808 24528 59872
rect 24208 58784 24528 59808
rect 24208 58720 24216 58784
rect 24280 58720 24296 58784
rect 24360 58720 24376 58784
rect 24440 58720 24456 58784
rect 24520 58720 24528 58784
rect 24208 57696 24528 58720
rect 24208 57632 24216 57696
rect 24280 57632 24296 57696
rect 24360 57632 24376 57696
rect 24440 57632 24456 57696
rect 24520 57632 24528 57696
rect 24208 56608 24528 57632
rect 24208 56544 24216 56608
rect 24280 56544 24296 56608
rect 24360 56544 24376 56608
rect 24440 56544 24456 56608
rect 24520 56544 24528 56608
rect 24208 55520 24528 56544
rect 24208 55456 24216 55520
rect 24280 55456 24296 55520
rect 24360 55456 24376 55520
rect 24440 55456 24456 55520
rect 24520 55456 24528 55520
rect 24208 54432 24528 55456
rect 24208 54368 24216 54432
rect 24280 54368 24296 54432
rect 24360 54368 24376 54432
rect 24440 54368 24456 54432
rect 24520 54368 24528 54432
rect 24208 53344 24528 54368
rect 24208 53280 24216 53344
rect 24280 53280 24296 53344
rect 24360 53280 24376 53344
rect 24440 53280 24456 53344
rect 24520 53280 24528 53344
rect 24208 52256 24528 53280
rect 24208 52192 24216 52256
rect 24280 52192 24296 52256
rect 24360 52192 24376 52256
rect 24440 52192 24456 52256
rect 24520 52192 24528 52256
rect 24208 51168 24528 52192
rect 24208 51104 24216 51168
rect 24280 51104 24296 51168
rect 24360 51104 24376 51168
rect 24440 51104 24456 51168
rect 24520 51104 24528 51168
rect 24208 50080 24528 51104
rect 24208 50016 24216 50080
rect 24280 50016 24296 50080
rect 24360 50016 24376 50080
rect 24440 50016 24456 50080
rect 24520 50016 24528 50080
rect 24208 48992 24528 50016
rect 24208 48928 24216 48992
rect 24280 48928 24296 48992
rect 24360 48928 24376 48992
rect 24440 48928 24456 48992
rect 24520 48928 24528 48992
rect 24208 47904 24528 48928
rect 24208 47840 24216 47904
rect 24280 47840 24296 47904
rect 24360 47840 24376 47904
rect 24440 47840 24456 47904
rect 24520 47840 24528 47904
rect 24208 46816 24528 47840
rect 24208 46752 24216 46816
rect 24280 46752 24296 46816
rect 24360 46752 24376 46816
rect 24440 46752 24456 46816
rect 24520 46752 24528 46816
rect 24208 45728 24528 46752
rect 24208 45664 24216 45728
rect 24280 45664 24296 45728
rect 24360 45664 24376 45728
rect 24440 45664 24456 45728
rect 24520 45664 24528 45728
rect 24208 44640 24528 45664
rect 24208 44576 24216 44640
rect 24280 44576 24296 44640
rect 24360 44576 24376 44640
rect 24440 44576 24456 44640
rect 24520 44576 24528 44640
rect 24208 43552 24528 44576
rect 24208 43488 24216 43552
rect 24280 43488 24296 43552
rect 24360 43488 24376 43552
rect 24440 43488 24456 43552
rect 24520 43488 24528 43552
rect 24208 42464 24528 43488
rect 24208 42400 24216 42464
rect 24280 42400 24296 42464
rect 24360 42400 24376 42464
rect 24440 42400 24456 42464
rect 24520 42400 24528 42464
rect 24208 41376 24528 42400
rect 24208 41312 24216 41376
rect 24280 41312 24296 41376
rect 24360 41312 24376 41376
rect 24440 41312 24456 41376
rect 24520 41312 24528 41376
rect 24208 40288 24528 41312
rect 24208 40224 24216 40288
rect 24280 40224 24296 40288
rect 24360 40224 24376 40288
rect 24440 40224 24456 40288
rect 24520 40224 24528 40288
rect 24208 39200 24528 40224
rect 24208 39136 24216 39200
rect 24280 39136 24296 39200
rect 24360 39136 24376 39200
rect 24440 39136 24456 39200
rect 24520 39136 24528 39200
rect 24208 38112 24528 39136
rect 24208 38048 24216 38112
rect 24280 38048 24296 38112
rect 24360 38048 24376 38112
rect 24440 38048 24456 38112
rect 24520 38048 24528 38112
rect 24208 37024 24528 38048
rect 24208 36960 24216 37024
rect 24280 36960 24296 37024
rect 24360 36960 24376 37024
rect 24440 36960 24456 37024
rect 24520 36960 24528 37024
rect 24208 35936 24528 36960
rect 24208 35872 24216 35936
rect 24280 35872 24296 35936
rect 24360 35872 24376 35936
rect 24440 35872 24456 35936
rect 24520 35872 24528 35936
rect 24208 34848 24528 35872
rect 24208 34784 24216 34848
rect 24280 34784 24296 34848
rect 24360 34784 24376 34848
rect 24440 34784 24456 34848
rect 24520 34784 24528 34848
rect 24208 33760 24528 34784
rect 24208 33696 24216 33760
rect 24280 33696 24296 33760
rect 24360 33696 24376 33760
rect 24440 33696 24456 33760
rect 24520 33696 24528 33760
rect 24208 32672 24528 33696
rect 24208 32608 24216 32672
rect 24280 32608 24296 32672
rect 24360 32608 24376 32672
rect 24440 32608 24456 32672
rect 24520 32608 24528 32672
rect 24208 31584 24528 32608
rect 24208 31520 24216 31584
rect 24280 31520 24296 31584
rect 24360 31520 24376 31584
rect 24440 31520 24456 31584
rect 24520 31520 24528 31584
rect 24208 30496 24528 31520
rect 24208 30432 24216 30496
rect 24280 30432 24296 30496
rect 24360 30432 24376 30496
rect 24440 30432 24456 30496
rect 24520 30432 24528 30496
rect 24208 29408 24528 30432
rect 24208 29344 24216 29408
rect 24280 29344 24296 29408
rect 24360 29344 24376 29408
rect 24440 29344 24456 29408
rect 24520 29344 24528 29408
rect 24208 28320 24528 29344
rect 24208 28256 24216 28320
rect 24280 28256 24296 28320
rect 24360 28256 24376 28320
rect 24440 28256 24456 28320
rect 24520 28256 24528 28320
rect 24208 27232 24528 28256
rect 24208 27168 24216 27232
rect 24280 27168 24296 27232
rect 24360 27168 24376 27232
rect 24440 27168 24456 27232
rect 24520 27168 24528 27232
rect 24208 26144 24528 27168
rect 24208 26080 24216 26144
rect 24280 26080 24296 26144
rect 24360 26080 24376 26144
rect 24440 26080 24456 26144
rect 24520 26080 24528 26144
rect 24208 25056 24528 26080
rect 24208 24992 24216 25056
rect 24280 24992 24296 25056
rect 24360 24992 24376 25056
rect 24440 24992 24456 25056
rect 24520 24992 24528 25056
rect 24208 23968 24528 24992
rect 24208 23904 24216 23968
rect 24280 23904 24296 23968
rect 24360 23904 24376 23968
rect 24440 23904 24456 23968
rect 24520 23904 24528 23968
rect 24208 22880 24528 23904
rect 24208 22816 24216 22880
rect 24280 22816 24296 22880
rect 24360 22816 24376 22880
rect 24440 22816 24456 22880
rect 24520 22816 24528 22880
rect 24208 21792 24528 22816
rect 24208 21728 24216 21792
rect 24280 21728 24296 21792
rect 24360 21728 24376 21792
rect 24440 21728 24456 21792
rect 24520 21728 24528 21792
rect 24208 20704 24528 21728
rect 24208 20640 24216 20704
rect 24280 20640 24296 20704
rect 24360 20640 24376 20704
rect 24440 20640 24456 20704
rect 24520 20640 24528 20704
rect 24208 19616 24528 20640
rect 24208 19552 24216 19616
rect 24280 19552 24296 19616
rect 24360 19552 24376 19616
rect 24440 19552 24456 19616
rect 24520 19552 24528 19616
rect 24208 15638 24528 19552
rect 24208 15574 24216 15638
rect 24280 15574 24296 15638
rect 24360 15574 24376 15638
rect 24440 15574 24456 15638
rect 24520 15574 24528 15638
rect 24208 15558 24528 15574
rect 24208 15494 24216 15558
rect 24280 15494 24296 15558
rect 24360 15494 24376 15558
rect 24440 15494 24456 15558
rect 24520 15494 24528 15558
rect 24208 15478 24528 15494
rect 24208 15414 24216 15478
rect 24280 15414 24296 15478
rect 24360 15414 24376 15478
rect 24440 15414 24456 15478
rect 24520 15414 24528 15478
rect 24208 15398 24528 15414
rect 24208 15334 24216 15398
rect 24280 15334 24296 15398
rect 24360 15334 24376 15398
rect 24440 15334 24456 15398
rect 24520 15334 24528 15398
rect 24208 15318 24528 15334
rect 24208 15254 24216 15318
rect 24280 15254 24296 15318
rect 24360 15254 24376 15318
rect 24440 15254 24456 15318
rect 24520 15254 24528 15318
rect 24208 11907 24528 15254
rect 24208 11843 24216 11907
rect 24280 11843 24296 11907
rect 24360 11843 24376 11907
rect 24440 11843 24456 11907
rect 24520 11843 24528 11907
rect 24208 11827 24528 11843
rect 24208 11763 24216 11827
rect 24280 11763 24296 11827
rect 24360 11763 24376 11827
rect 24440 11763 24456 11827
rect 24520 11763 24528 11827
rect 24208 11747 24528 11763
rect 24208 11683 24216 11747
rect 24280 11683 24296 11747
rect 24360 11683 24376 11747
rect 24440 11683 24456 11747
rect 24520 11683 24528 11747
rect 24208 11667 24528 11683
rect 24208 11603 24216 11667
rect 24280 11603 24296 11667
rect 24360 11603 24376 11667
rect 24440 11603 24456 11667
rect 24520 11603 24528 11667
rect 24208 9358 24528 11603
rect 24208 9294 24216 9358
rect 24280 9294 24296 9358
rect 24360 9294 24376 9358
rect 24440 9294 24456 9358
rect 24520 9294 24528 9358
rect 24208 9278 24528 9294
rect 24208 9214 24216 9278
rect 24280 9214 24296 9278
rect 24360 9214 24376 9278
rect 24440 9214 24456 9278
rect 24520 9214 24528 9278
rect 24208 9198 24528 9214
rect 24208 9134 24216 9198
rect 24280 9134 24296 9198
rect 24360 9134 24376 9198
rect 24440 9134 24456 9198
rect 24520 9134 24528 9198
rect 24208 9118 24528 9134
rect 24208 9054 24216 9118
rect 24280 9054 24296 9118
rect 24360 9054 24376 9118
rect 24440 9054 24456 9118
rect 24520 9054 24528 9118
rect 24208 6809 24528 9054
rect 24208 6745 24216 6809
rect 24280 6745 24296 6809
rect 24360 6745 24376 6809
rect 24440 6745 24456 6809
rect 24520 6745 24528 6809
rect 24208 6729 24528 6745
rect 24208 6665 24216 6729
rect 24280 6665 24296 6729
rect 24360 6665 24376 6729
rect 24440 6665 24456 6729
rect 24520 6665 24528 6729
rect 24208 6649 24528 6665
rect 24208 6585 24216 6649
rect 24280 6585 24296 6649
rect 24360 6585 24376 6649
rect 24440 6585 24456 6649
rect 24520 6585 24528 6649
rect 24208 6569 24528 6585
rect 24208 6505 24216 6569
rect 24280 6505 24296 6569
rect 24360 6505 24376 6569
rect 24440 6505 24456 6569
rect 24520 6505 24528 6569
rect 24208 3222 24528 6505
rect 29208 66944 29528 67504
rect 29208 66880 29216 66944
rect 29280 66880 29296 66944
rect 29360 66880 29376 66944
rect 29440 66880 29456 66944
rect 29520 66880 29528 66944
rect 29208 65856 29528 66880
rect 29208 65792 29216 65856
rect 29280 65792 29296 65856
rect 29360 65792 29376 65856
rect 29440 65792 29456 65856
rect 29520 65792 29528 65856
rect 29208 64768 29528 65792
rect 29208 64704 29216 64768
rect 29280 64704 29296 64768
rect 29360 64704 29376 64768
rect 29440 64704 29456 64768
rect 29520 64704 29528 64768
rect 29208 63680 29528 64704
rect 29208 63616 29216 63680
rect 29280 63616 29296 63680
rect 29360 63616 29376 63680
rect 29440 63616 29456 63680
rect 29520 63616 29528 63680
rect 29208 62592 29528 63616
rect 29208 62528 29216 62592
rect 29280 62528 29296 62592
rect 29360 62528 29376 62592
rect 29440 62528 29456 62592
rect 29520 62528 29528 62592
rect 29208 61504 29528 62528
rect 29208 61440 29216 61504
rect 29280 61440 29296 61504
rect 29360 61440 29376 61504
rect 29440 61440 29456 61504
rect 29520 61440 29528 61504
rect 29208 60416 29528 61440
rect 29208 60352 29216 60416
rect 29280 60352 29296 60416
rect 29360 60352 29376 60416
rect 29440 60352 29456 60416
rect 29520 60352 29528 60416
rect 29208 59328 29528 60352
rect 29208 59264 29216 59328
rect 29280 59264 29296 59328
rect 29360 59264 29376 59328
rect 29440 59264 29456 59328
rect 29520 59264 29528 59328
rect 29208 58240 29528 59264
rect 29208 58176 29216 58240
rect 29280 58176 29296 58240
rect 29360 58176 29376 58240
rect 29440 58176 29456 58240
rect 29520 58176 29528 58240
rect 29208 57152 29528 58176
rect 29208 57088 29216 57152
rect 29280 57088 29296 57152
rect 29360 57088 29376 57152
rect 29440 57088 29456 57152
rect 29520 57088 29528 57152
rect 29208 56064 29528 57088
rect 29208 56000 29216 56064
rect 29280 56000 29296 56064
rect 29360 56000 29376 56064
rect 29440 56000 29456 56064
rect 29520 56000 29528 56064
rect 29208 54976 29528 56000
rect 29208 54912 29216 54976
rect 29280 54912 29296 54976
rect 29360 54912 29376 54976
rect 29440 54912 29456 54976
rect 29520 54912 29528 54976
rect 29208 53888 29528 54912
rect 29208 53824 29216 53888
rect 29280 53824 29296 53888
rect 29360 53824 29376 53888
rect 29440 53824 29456 53888
rect 29520 53824 29528 53888
rect 29208 52800 29528 53824
rect 29208 52736 29216 52800
rect 29280 52736 29296 52800
rect 29360 52736 29376 52800
rect 29440 52736 29456 52800
rect 29520 52736 29528 52800
rect 29208 51712 29528 52736
rect 29208 51648 29216 51712
rect 29280 51648 29296 51712
rect 29360 51648 29376 51712
rect 29440 51648 29456 51712
rect 29520 51648 29528 51712
rect 29208 50624 29528 51648
rect 29208 50560 29216 50624
rect 29280 50560 29296 50624
rect 29360 50560 29376 50624
rect 29440 50560 29456 50624
rect 29520 50560 29528 50624
rect 29208 49536 29528 50560
rect 29208 49472 29216 49536
rect 29280 49472 29296 49536
rect 29360 49472 29376 49536
rect 29440 49472 29456 49536
rect 29520 49472 29528 49536
rect 29208 48448 29528 49472
rect 29208 48384 29216 48448
rect 29280 48384 29296 48448
rect 29360 48384 29376 48448
rect 29440 48384 29456 48448
rect 29520 48384 29528 48448
rect 29208 47360 29528 48384
rect 29208 47296 29216 47360
rect 29280 47296 29296 47360
rect 29360 47296 29376 47360
rect 29440 47296 29456 47360
rect 29520 47296 29528 47360
rect 29208 46272 29528 47296
rect 29208 46208 29216 46272
rect 29280 46208 29296 46272
rect 29360 46208 29376 46272
rect 29440 46208 29456 46272
rect 29520 46208 29528 46272
rect 29208 45184 29528 46208
rect 29208 45120 29216 45184
rect 29280 45120 29296 45184
rect 29360 45120 29376 45184
rect 29440 45120 29456 45184
rect 29520 45120 29528 45184
rect 29208 44096 29528 45120
rect 29208 44032 29216 44096
rect 29280 44032 29296 44096
rect 29360 44032 29376 44096
rect 29440 44032 29456 44096
rect 29520 44032 29528 44096
rect 29208 43008 29528 44032
rect 29208 42944 29216 43008
rect 29280 42944 29296 43008
rect 29360 42944 29376 43008
rect 29440 42944 29456 43008
rect 29520 42944 29528 43008
rect 29208 41920 29528 42944
rect 29208 41856 29216 41920
rect 29280 41856 29296 41920
rect 29360 41856 29376 41920
rect 29440 41856 29456 41920
rect 29520 41856 29528 41920
rect 29208 40832 29528 41856
rect 29208 40768 29216 40832
rect 29280 40768 29296 40832
rect 29360 40768 29376 40832
rect 29440 40768 29456 40832
rect 29520 40768 29528 40832
rect 29208 39744 29528 40768
rect 29208 39680 29216 39744
rect 29280 39680 29296 39744
rect 29360 39680 29376 39744
rect 29440 39680 29456 39744
rect 29520 39680 29528 39744
rect 29208 38656 29528 39680
rect 29208 38592 29216 38656
rect 29280 38592 29296 38656
rect 29360 38592 29376 38656
rect 29440 38592 29456 38656
rect 29520 38592 29528 38656
rect 29208 37568 29528 38592
rect 29208 37504 29216 37568
rect 29280 37504 29296 37568
rect 29360 37504 29376 37568
rect 29440 37504 29456 37568
rect 29520 37504 29528 37568
rect 29208 36480 29528 37504
rect 29208 36416 29216 36480
rect 29280 36416 29296 36480
rect 29360 36416 29376 36480
rect 29440 36416 29456 36480
rect 29520 36416 29528 36480
rect 29208 35392 29528 36416
rect 29208 35328 29216 35392
rect 29280 35328 29296 35392
rect 29360 35328 29376 35392
rect 29440 35328 29456 35392
rect 29520 35328 29528 35392
rect 29208 34304 29528 35328
rect 29208 34240 29216 34304
rect 29280 34240 29296 34304
rect 29360 34240 29376 34304
rect 29440 34240 29456 34304
rect 29520 34240 29528 34304
rect 29208 33216 29528 34240
rect 29208 33152 29216 33216
rect 29280 33152 29296 33216
rect 29360 33152 29376 33216
rect 29440 33152 29456 33216
rect 29520 33152 29528 33216
rect 29208 32128 29528 33152
rect 29208 32064 29216 32128
rect 29280 32064 29296 32128
rect 29360 32064 29376 32128
rect 29440 32064 29456 32128
rect 29520 32064 29528 32128
rect 29208 31040 29528 32064
rect 29208 30976 29216 31040
rect 29280 30976 29296 31040
rect 29360 30976 29376 31040
rect 29440 30976 29456 31040
rect 29520 30976 29528 31040
rect 29208 29952 29528 30976
rect 29208 29888 29216 29952
rect 29280 29888 29296 29952
rect 29360 29888 29376 29952
rect 29440 29888 29456 29952
rect 29520 29888 29528 29952
rect 29208 28864 29528 29888
rect 29208 28800 29216 28864
rect 29280 28800 29296 28864
rect 29360 28800 29376 28864
rect 29440 28800 29456 28864
rect 29520 28800 29528 28864
rect 29208 27776 29528 28800
rect 29208 27712 29216 27776
rect 29280 27712 29296 27776
rect 29360 27712 29376 27776
rect 29440 27712 29456 27776
rect 29520 27712 29528 27776
rect 29208 26688 29528 27712
rect 29208 26624 29216 26688
rect 29280 26624 29296 26688
rect 29360 26624 29376 26688
rect 29440 26624 29456 26688
rect 29520 26624 29528 26688
rect 29208 25600 29528 26624
rect 29208 25536 29216 25600
rect 29280 25536 29296 25600
rect 29360 25536 29376 25600
rect 29440 25536 29456 25600
rect 29520 25536 29528 25600
rect 29208 24512 29528 25536
rect 29208 24448 29216 24512
rect 29280 24448 29296 24512
rect 29360 24448 29376 24512
rect 29440 24448 29456 24512
rect 29520 24448 29528 24512
rect 29208 23424 29528 24448
rect 29208 23360 29216 23424
rect 29280 23360 29296 23424
rect 29360 23360 29376 23424
rect 29440 23360 29456 23424
rect 29520 23360 29528 23424
rect 29208 22336 29528 23360
rect 29208 22272 29216 22336
rect 29280 22272 29296 22336
rect 29360 22272 29376 22336
rect 29440 22272 29456 22336
rect 29520 22272 29528 22336
rect 29208 21248 29528 22272
rect 29208 21184 29216 21248
rect 29280 21184 29296 21248
rect 29360 21184 29376 21248
rect 29440 21184 29456 21248
rect 29520 21184 29528 21248
rect 29208 20160 29528 21184
rect 29208 20096 29216 20160
rect 29280 20096 29296 20160
rect 29360 20096 29376 20160
rect 29440 20096 29456 20160
rect 29520 20096 29528 20160
rect 29208 16438 29528 20096
rect 29208 16374 29216 16438
rect 29280 16374 29296 16438
rect 29360 16374 29376 16438
rect 29440 16374 29456 16438
rect 29520 16374 29528 16438
rect 29208 16358 29528 16374
rect 29208 16294 29216 16358
rect 29280 16294 29296 16358
rect 29360 16294 29376 16358
rect 29440 16294 29456 16358
rect 29520 16294 29528 16358
rect 29208 16278 29528 16294
rect 29208 16214 29216 16278
rect 29280 16214 29296 16278
rect 29360 16214 29376 16278
rect 29440 16214 29456 16278
rect 29520 16214 29528 16278
rect 29208 16198 29528 16214
rect 29208 16134 29216 16198
rect 29280 16134 29296 16198
rect 29360 16134 29376 16198
rect 29440 16134 29456 16198
rect 29520 16134 29528 16198
rect 29208 16118 29528 16134
rect 29208 16054 29216 16118
rect 29280 16054 29296 16118
rect 29360 16054 29376 16118
rect 29440 16054 29456 16118
rect 29520 16054 29528 16118
rect 29208 10633 29528 16054
rect 29208 10569 29216 10633
rect 29280 10569 29296 10633
rect 29360 10569 29376 10633
rect 29440 10569 29456 10633
rect 29520 10569 29528 10633
rect 29208 10553 29528 10569
rect 29208 10489 29216 10553
rect 29280 10489 29296 10553
rect 29360 10489 29376 10553
rect 29440 10489 29456 10553
rect 29520 10489 29528 10553
rect 29208 10473 29528 10489
rect 29208 10409 29216 10473
rect 29280 10409 29296 10473
rect 29360 10409 29376 10473
rect 29440 10409 29456 10473
rect 29520 10409 29528 10473
rect 29208 10393 29528 10409
rect 29208 10329 29216 10393
rect 29280 10329 29296 10393
rect 29360 10329 29376 10393
rect 29440 10329 29456 10393
rect 29520 10329 29528 10393
rect 29208 8083 29528 10329
rect 29208 8019 29216 8083
rect 29280 8019 29296 8083
rect 29360 8019 29376 8083
rect 29440 8019 29456 8083
rect 29520 8019 29528 8083
rect 29208 8003 29528 8019
rect 29208 7939 29216 8003
rect 29280 7939 29296 8003
rect 29360 7939 29376 8003
rect 29440 7939 29456 8003
rect 29520 7939 29528 8003
rect 29208 7923 29528 7939
rect 29208 7859 29216 7923
rect 29280 7859 29296 7923
rect 29360 7859 29376 7923
rect 29440 7859 29456 7923
rect 29520 7859 29528 7923
rect 29208 7843 29528 7859
rect 29208 7779 29216 7843
rect 29280 7779 29296 7843
rect 29360 7779 29376 7843
rect 29440 7779 29456 7843
rect 29520 7779 29528 7843
rect 27659 5948 27725 5949
rect 27659 5884 27660 5948
rect 27724 5884 27725 5948
rect 27659 5883 27725 5884
rect 24208 3158 24216 3222
rect 24280 3158 24296 3222
rect 24360 3158 24376 3222
rect 24440 3158 24456 3222
rect 24520 3158 24528 3222
rect 24208 3142 24528 3158
rect 24208 3078 24216 3142
rect 24280 3078 24296 3142
rect 24360 3078 24376 3142
rect 24440 3078 24456 3142
rect 24520 3078 24528 3142
rect 24208 3062 24528 3078
rect 24208 2998 24216 3062
rect 24280 2998 24296 3062
rect 24360 2998 24376 3062
rect 24440 2998 24456 3062
rect 24520 2998 24528 3062
rect 24208 2982 24528 2998
rect 24208 2918 24216 2982
rect 24280 2918 24296 2982
rect 24360 2918 24376 2982
rect 24440 2918 24456 2982
rect 24520 2918 24528 2982
rect 24208 2902 24528 2918
rect 24208 2838 24216 2902
rect 24280 2838 24296 2902
rect 24360 2838 24376 2902
rect 24440 2838 24456 2902
rect 24520 2838 24528 2902
rect 24208 2176 24528 2838
rect 14208 2128 14528 2144
rect 5395 2004 5461 2005
rect 5395 1940 5396 2004
rect 5460 1940 5461 2004
rect 5395 1939 5461 1940
rect 27662 1869 27722 5883
rect 28211 3772 28277 3773
rect 28211 3708 28212 3772
rect 28276 3708 28277 3772
rect 28211 3707 28277 3708
rect 28027 3636 28093 3637
rect 28027 3572 28028 3636
rect 28092 3572 28093 3636
rect 28027 3571 28093 3572
rect 28030 1869 28090 3571
rect 27659 1868 27725 1869
rect 27659 1804 27660 1868
rect 27724 1804 27725 1868
rect 27659 1803 27725 1804
rect 28027 1868 28093 1869
rect 28027 1804 28028 1868
rect 28092 1804 28093 1868
rect 28027 1803 28093 1804
rect 28214 1733 28274 3707
rect 29208 2430 29528 7779
rect 34208 67488 34528 67504
rect 34208 67424 34216 67488
rect 34280 67424 34296 67488
rect 34360 67424 34376 67488
rect 34440 67424 34456 67488
rect 34520 67424 34528 67488
rect 34208 66400 34528 67424
rect 34208 66336 34216 66400
rect 34280 66336 34296 66400
rect 34360 66336 34376 66400
rect 34440 66336 34456 66400
rect 34520 66336 34528 66400
rect 34208 65312 34528 66336
rect 34208 65248 34216 65312
rect 34280 65248 34296 65312
rect 34360 65248 34376 65312
rect 34440 65248 34456 65312
rect 34520 65248 34528 65312
rect 34208 64224 34528 65248
rect 34208 64160 34216 64224
rect 34280 64160 34296 64224
rect 34360 64160 34376 64224
rect 34440 64160 34456 64224
rect 34520 64160 34528 64224
rect 34208 63136 34528 64160
rect 34208 63072 34216 63136
rect 34280 63072 34296 63136
rect 34360 63072 34376 63136
rect 34440 63072 34456 63136
rect 34520 63072 34528 63136
rect 34208 62048 34528 63072
rect 34208 61984 34216 62048
rect 34280 61984 34296 62048
rect 34360 61984 34376 62048
rect 34440 61984 34456 62048
rect 34520 61984 34528 62048
rect 34208 60960 34528 61984
rect 34208 60896 34216 60960
rect 34280 60896 34296 60960
rect 34360 60896 34376 60960
rect 34440 60896 34456 60960
rect 34520 60896 34528 60960
rect 34208 59872 34528 60896
rect 34208 59808 34216 59872
rect 34280 59808 34296 59872
rect 34360 59808 34376 59872
rect 34440 59808 34456 59872
rect 34520 59808 34528 59872
rect 34208 58784 34528 59808
rect 34208 58720 34216 58784
rect 34280 58720 34296 58784
rect 34360 58720 34376 58784
rect 34440 58720 34456 58784
rect 34520 58720 34528 58784
rect 34208 57696 34528 58720
rect 34208 57632 34216 57696
rect 34280 57632 34296 57696
rect 34360 57632 34376 57696
rect 34440 57632 34456 57696
rect 34520 57632 34528 57696
rect 34208 56608 34528 57632
rect 34208 56544 34216 56608
rect 34280 56544 34296 56608
rect 34360 56544 34376 56608
rect 34440 56544 34456 56608
rect 34520 56544 34528 56608
rect 34208 55520 34528 56544
rect 34208 55456 34216 55520
rect 34280 55456 34296 55520
rect 34360 55456 34376 55520
rect 34440 55456 34456 55520
rect 34520 55456 34528 55520
rect 34208 54432 34528 55456
rect 34208 54368 34216 54432
rect 34280 54368 34296 54432
rect 34360 54368 34376 54432
rect 34440 54368 34456 54432
rect 34520 54368 34528 54432
rect 34208 53344 34528 54368
rect 34208 53280 34216 53344
rect 34280 53280 34296 53344
rect 34360 53280 34376 53344
rect 34440 53280 34456 53344
rect 34520 53280 34528 53344
rect 34208 52256 34528 53280
rect 34208 52192 34216 52256
rect 34280 52192 34296 52256
rect 34360 52192 34376 52256
rect 34440 52192 34456 52256
rect 34520 52192 34528 52256
rect 34208 51168 34528 52192
rect 34208 51104 34216 51168
rect 34280 51104 34296 51168
rect 34360 51104 34376 51168
rect 34440 51104 34456 51168
rect 34520 51104 34528 51168
rect 34208 50080 34528 51104
rect 34208 50016 34216 50080
rect 34280 50016 34296 50080
rect 34360 50016 34376 50080
rect 34440 50016 34456 50080
rect 34520 50016 34528 50080
rect 34208 48992 34528 50016
rect 34208 48928 34216 48992
rect 34280 48928 34296 48992
rect 34360 48928 34376 48992
rect 34440 48928 34456 48992
rect 34520 48928 34528 48992
rect 34208 47904 34528 48928
rect 34208 47840 34216 47904
rect 34280 47840 34296 47904
rect 34360 47840 34376 47904
rect 34440 47840 34456 47904
rect 34520 47840 34528 47904
rect 34208 46816 34528 47840
rect 34208 46752 34216 46816
rect 34280 46752 34296 46816
rect 34360 46752 34376 46816
rect 34440 46752 34456 46816
rect 34520 46752 34528 46816
rect 34208 45728 34528 46752
rect 34208 45664 34216 45728
rect 34280 45664 34296 45728
rect 34360 45664 34376 45728
rect 34440 45664 34456 45728
rect 34520 45664 34528 45728
rect 34208 44640 34528 45664
rect 34208 44576 34216 44640
rect 34280 44576 34296 44640
rect 34360 44576 34376 44640
rect 34440 44576 34456 44640
rect 34520 44576 34528 44640
rect 34208 43552 34528 44576
rect 34208 43488 34216 43552
rect 34280 43488 34296 43552
rect 34360 43488 34376 43552
rect 34440 43488 34456 43552
rect 34520 43488 34528 43552
rect 34208 42464 34528 43488
rect 34208 42400 34216 42464
rect 34280 42400 34296 42464
rect 34360 42400 34376 42464
rect 34440 42400 34456 42464
rect 34520 42400 34528 42464
rect 34208 41376 34528 42400
rect 34208 41312 34216 41376
rect 34280 41312 34296 41376
rect 34360 41312 34376 41376
rect 34440 41312 34456 41376
rect 34520 41312 34528 41376
rect 34208 40288 34528 41312
rect 34208 40224 34216 40288
rect 34280 40224 34296 40288
rect 34360 40224 34376 40288
rect 34440 40224 34456 40288
rect 34520 40224 34528 40288
rect 34208 39200 34528 40224
rect 34208 39136 34216 39200
rect 34280 39136 34296 39200
rect 34360 39136 34376 39200
rect 34440 39136 34456 39200
rect 34520 39136 34528 39200
rect 34208 38112 34528 39136
rect 34208 38048 34216 38112
rect 34280 38048 34296 38112
rect 34360 38048 34376 38112
rect 34440 38048 34456 38112
rect 34520 38048 34528 38112
rect 34208 37024 34528 38048
rect 34208 36960 34216 37024
rect 34280 36960 34296 37024
rect 34360 36960 34376 37024
rect 34440 36960 34456 37024
rect 34520 36960 34528 37024
rect 34208 35936 34528 36960
rect 34208 35872 34216 35936
rect 34280 35872 34296 35936
rect 34360 35872 34376 35936
rect 34440 35872 34456 35936
rect 34520 35872 34528 35936
rect 34208 34848 34528 35872
rect 34208 34784 34216 34848
rect 34280 34784 34296 34848
rect 34360 34784 34376 34848
rect 34440 34784 34456 34848
rect 34520 34784 34528 34848
rect 34208 33760 34528 34784
rect 34208 33696 34216 33760
rect 34280 33696 34296 33760
rect 34360 33696 34376 33760
rect 34440 33696 34456 33760
rect 34520 33696 34528 33760
rect 34208 32672 34528 33696
rect 34208 32608 34216 32672
rect 34280 32608 34296 32672
rect 34360 32608 34376 32672
rect 34440 32608 34456 32672
rect 34520 32608 34528 32672
rect 34208 31584 34528 32608
rect 39208 66944 39528 67504
rect 39208 66880 39216 66944
rect 39280 66880 39296 66944
rect 39360 66880 39376 66944
rect 39440 66880 39456 66944
rect 39520 66880 39528 66944
rect 39208 65856 39528 66880
rect 39208 65792 39216 65856
rect 39280 65792 39296 65856
rect 39360 65792 39376 65856
rect 39440 65792 39456 65856
rect 39520 65792 39528 65856
rect 39208 64768 39528 65792
rect 39208 64704 39216 64768
rect 39280 64704 39296 64768
rect 39360 64704 39376 64768
rect 39440 64704 39456 64768
rect 39520 64704 39528 64768
rect 39208 63680 39528 64704
rect 39208 63616 39216 63680
rect 39280 63616 39296 63680
rect 39360 63616 39376 63680
rect 39440 63616 39456 63680
rect 39520 63616 39528 63680
rect 39208 62592 39528 63616
rect 39208 62528 39216 62592
rect 39280 62528 39296 62592
rect 39360 62528 39376 62592
rect 39440 62528 39456 62592
rect 39520 62528 39528 62592
rect 39208 61504 39528 62528
rect 39208 61440 39216 61504
rect 39280 61440 39296 61504
rect 39360 61440 39376 61504
rect 39440 61440 39456 61504
rect 39520 61440 39528 61504
rect 39208 60416 39528 61440
rect 39208 60352 39216 60416
rect 39280 60352 39296 60416
rect 39360 60352 39376 60416
rect 39440 60352 39456 60416
rect 39520 60352 39528 60416
rect 39208 59328 39528 60352
rect 39208 59264 39216 59328
rect 39280 59264 39296 59328
rect 39360 59264 39376 59328
rect 39440 59264 39456 59328
rect 39520 59264 39528 59328
rect 39208 58240 39528 59264
rect 39208 58176 39216 58240
rect 39280 58176 39296 58240
rect 39360 58176 39376 58240
rect 39440 58176 39456 58240
rect 39520 58176 39528 58240
rect 39208 57152 39528 58176
rect 39208 57088 39216 57152
rect 39280 57088 39296 57152
rect 39360 57088 39376 57152
rect 39440 57088 39456 57152
rect 39520 57088 39528 57152
rect 39208 56064 39528 57088
rect 39208 56000 39216 56064
rect 39280 56000 39296 56064
rect 39360 56000 39376 56064
rect 39440 56000 39456 56064
rect 39520 56000 39528 56064
rect 39208 54976 39528 56000
rect 39208 54912 39216 54976
rect 39280 54912 39296 54976
rect 39360 54912 39376 54976
rect 39440 54912 39456 54976
rect 39520 54912 39528 54976
rect 39208 53888 39528 54912
rect 39208 53824 39216 53888
rect 39280 53824 39296 53888
rect 39360 53824 39376 53888
rect 39440 53824 39456 53888
rect 39520 53824 39528 53888
rect 39208 52800 39528 53824
rect 39208 52736 39216 52800
rect 39280 52736 39296 52800
rect 39360 52736 39376 52800
rect 39440 52736 39456 52800
rect 39520 52736 39528 52800
rect 39208 51712 39528 52736
rect 39208 51648 39216 51712
rect 39280 51648 39296 51712
rect 39360 51648 39376 51712
rect 39440 51648 39456 51712
rect 39520 51648 39528 51712
rect 39208 50624 39528 51648
rect 39208 50560 39216 50624
rect 39280 50560 39296 50624
rect 39360 50560 39376 50624
rect 39440 50560 39456 50624
rect 39520 50560 39528 50624
rect 39208 49536 39528 50560
rect 39208 49472 39216 49536
rect 39280 49472 39296 49536
rect 39360 49472 39376 49536
rect 39440 49472 39456 49536
rect 39520 49472 39528 49536
rect 39208 48448 39528 49472
rect 39208 48384 39216 48448
rect 39280 48384 39296 48448
rect 39360 48384 39376 48448
rect 39440 48384 39456 48448
rect 39520 48384 39528 48448
rect 39208 47360 39528 48384
rect 39208 47296 39216 47360
rect 39280 47296 39296 47360
rect 39360 47296 39376 47360
rect 39440 47296 39456 47360
rect 39520 47296 39528 47360
rect 39208 46272 39528 47296
rect 39208 46208 39216 46272
rect 39280 46208 39296 46272
rect 39360 46208 39376 46272
rect 39440 46208 39456 46272
rect 39520 46208 39528 46272
rect 39208 45184 39528 46208
rect 39208 45120 39216 45184
rect 39280 45120 39296 45184
rect 39360 45120 39376 45184
rect 39440 45120 39456 45184
rect 39520 45120 39528 45184
rect 39208 44096 39528 45120
rect 39208 44032 39216 44096
rect 39280 44032 39296 44096
rect 39360 44032 39376 44096
rect 39440 44032 39456 44096
rect 39520 44032 39528 44096
rect 39208 43008 39528 44032
rect 39208 42944 39216 43008
rect 39280 42944 39296 43008
rect 39360 42944 39376 43008
rect 39440 42944 39456 43008
rect 39520 42944 39528 43008
rect 39208 41920 39528 42944
rect 39208 41856 39216 41920
rect 39280 41856 39296 41920
rect 39360 41856 39376 41920
rect 39440 41856 39456 41920
rect 39520 41856 39528 41920
rect 39208 40832 39528 41856
rect 39208 40768 39216 40832
rect 39280 40768 39296 40832
rect 39360 40768 39376 40832
rect 39440 40768 39456 40832
rect 39520 40768 39528 40832
rect 39208 39744 39528 40768
rect 39208 39680 39216 39744
rect 39280 39680 39296 39744
rect 39360 39680 39376 39744
rect 39440 39680 39456 39744
rect 39520 39680 39528 39744
rect 39208 38656 39528 39680
rect 39208 38592 39216 38656
rect 39280 38592 39296 38656
rect 39360 38592 39376 38656
rect 39440 38592 39456 38656
rect 39520 38592 39528 38656
rect 39208 37568 39528 38592
rect 39208 37504 39216 37568
rect 39280 37504 39296 37568
rect 39360 37504 39376 37568
rect 39440 37504 39456 37568
rect 39520 37504 39528 37568
rect 39208 36480 39528 37504
rect 39208 36416 39216 36480
rect 39280 36416 39296 36480
rect 39360 36416 39376 36480
rect 39440 36416 39456 36480
rect 39520 36416 39528 36480
rect 39208 35392 39528 36416
rect 39208 35328 39216 35392
rect 39280 35328 39296 35392
rect 39360 35328 39376 35392
rect 39440 35328 39456 35392
rect 39520 35328 39528 35392
rect 39208 34304 39528 35328
rect 39208 34240 39216 34304
rect 39280 34240 39296 34304
rect 39360 34240 39376 34304
rect 39440 34240 39456 34304
rect 39520 34240 39528 34304
rect 39208 33216 39528 34240
rect 39208 33152 39216 33216
rect 39280 33152 39296 33216
rect 39360 33152 39376 33216
rect 39440 33152 39456 33216
rect 39520 33152 39528 33216
rect 38699 32468 38765 32469
rect 38699 32404 38700 32468
rect 38764 32404 38765 32468
rect 38699 32403 38765 32404
rect 34208 31520 34216 31584
rect 34280 31520 34296 31584
rect 34360 31520 34376 31584
rect 34440 31520 34456 31584
rect 34520 31520 34528 31584
rect 34208 30496 34528 31520
rect 34208 30432 34216 30496
rect 34280 30432 34296 30496
rect 34360 30432 34376 30496
rect 34440 30432 34456 30496
rect 34520 30432 34528 30496
rect 34208 29408 34528 30432
rect 34208 29344 34216 29408
rect 34280 29344 34296 29408
rect 34360 29344 34376 29408
rect 34440 29344 34456 29408
rect 34520 29344 34528 29408
rect 34208 28320 34528 29344
rect 34208 28256 34216 28320
rect 34280 28256 34296 28320
rect 34360 28256 34376 28320
rect 34440 28256 34456 28320
rect 34520 28256 34528 28320
rect 34208 27232 34528 28256
rect 34208 27168 34216 27232
rect 34280 27168 34296 27232
rect 34360 27168 34376 27232
rect 34440 27168 34456 27232
rect 34520 27168 34528 27232
rect 34208 26144 34528 27168
rect 34208 26080 34216 26144
rect 34280 26080 34296 26144
rect 34360 26080 34376 26144
rect 34440 26080 34456 26144
rect 34520 26080 34528 26144
rect 34208 25056 34528 26080
rect 34208 24992 34216 25056
rect 34280 24992 34296 25056
rect 34360 24992 34376 25056
rect 34440 24992 34456 25056
rect 34520 24992 34528 25056
rect 34208 23968 34528 24992
rect 34208 23904 34216 23968
rect 34280 23904 34296 23968
rect 34360 23904 34376 23968
rect 34440 23904 34456 23968
rect 34520 23904 34528 23968
rect 34208 22880 34528 23904
rect 34208 22816 34216 22880
rect 34280 22816 34296 22880
rect 34360 22816 34376 22880
rect 34440 22816 34456 22880
rect 34520 22816 34528 22880
rect 34208 21792 34528 22816
rect 34208 21728 34216 21792
rect 34280 21728 34296 21792
rect 34360 21728 34376 21792
rect 34440 21728 34456 21792
rect 34520 21728 34528 21792
rect 34208 20704 34528 21728
rect 34208 20640 34216 20704
rect 34280 20640 34296 20704
rect 34360 20640 34376 20704
rect 34440 20640 34456 20704
rect 34520 20640 34528 20704
rect 34208 19616 34528 20640
rect 34208 19552 34216 19616
rect 34280 19552 34296 19616
rect 34360 19552 34376 19616
rect 34440 19552 34456 19616
rect 34520 19552 34528 19616
rect 34208 11907 34528 19552
rect 38702 12205 38762 32403
rect 39208 32128 39528 33152
rect 39208 32064 39216 32128
rect 39280 32064 39296 32128
rect 39360 32064 39376 32128
rect 39440 32064 39456 32128
rect 39520 32064 39528 32128
rect 39208 31040 39528 32064
rect 39208 30976 39216 31040
rect 39280 30976 39296 31040
rect 39360 30976 39376 31040
rect 39440 30976 39456 31040
rect 39520 30976 39528 31040
rect 39208 29952 39528 30976
rect 39208 29888 39216 29952
rect 39280 29888 39296 29952
rect 39360 29888 39376 29952
rect 39440 29888 39456 29952
rect 39520 29888 39528 29952
rect 39208 28864 39528 29888
rect 39208 28800 39216 28864
rect 39280 28800 39296 28864
rect 39360 28800 39376 28864
rect 39440 28800 39456 28864
rect 39520 28800 39528 28864
rect 39208 27776 39528 28800
rect 39208 27712 39216 27776
rect 39280 27712 39296 27776
rect 39360 27712 39376 27776
rect 39440 27712 39456 27776
rect 39520 27712 39528 27776
rect 39208 26688 39528 27712
rect 39208 26624 39216 26688
rect 39280 26624 39296 26688
rect 39360 26624 39376 26688
rect 39440 26624 39456 26688
rect 39520 26624 39528 26688
rect 39208 25600 39528 26624
rect 39208 25536 39216 25600
rect 39280 25536 39296 25600
rect 39360 25536 39376 25600
rect 39440 25536 39456 25600
rect 39520 25536 39528 25600
rect 39208 24512 39528 25536
rect 39208 24448 39216 24512
rect 39280 24448 39296 24512
rect 39360 24448 39376 24512
rect 39440 24448 39456 24512
rect 39520 24448 39528 24512
rect 39208 23424 39528 24448
rect 39208 23360 39216 23424
rect 39280 23360 39296 23424
rect 39360 23360 39376 23424
rect 39440 23360 39456 23424
rect 39520 23360 39528 23424
rect 39208 22336 39528 23360
rect 39208 22272 39216 22336
rect 39280 22272 39296 22336
rect 39360 22272 39376 22336
rect 39440 22272 39456 22336
rect 39520 22272 39528 22336
rect 39067 21452 39133 21453
rect 39067 21388 39068 21452
rect 39132 21388 39133 21452
rect 39067 21387 39133 21388
rect 39070 13157 39130 21387
rect 39208 21248 39528 22272
rect 39208 21184 39216 21248
rect 39280 21184 39296 21248
rect 39360 21184 39376 21248
rect 39440 21184 39456 21248
rect 39520 21184 39528 21248
rect 39208 20160 39528 21184
rect 39208 20096 39216 20160
rect 39280 20096 39296 20160
rect 39360 20096 39376 20160
rect 39440 20096 39456 20160
rect 39520 20096 39528 20160
rect 39208 19072 39528 20096
rect 39208 19008 39216 19072
rect 39280 19008 39296 19072
rect 39360 19008 39376 19072
rect 39440 19008 39456 19072
rect 39520 19008 39528 19072
rect 39208 17984 39528 19008
rect 39208 17920 39216 17984
rect 39280 17920 39296 17984
rect 39360 17920 39376 17984
rect 39440 17920 39456 17984
rect 39520 17920 39528 17984
rect 39208 16896 39528 17920
rect 44208 67488 44528 67504
rect 44208 67424 44216 67488
rect 44280 67424 44296 67488
rect 44360 67424 44376 67488
rect 44440 67424 44456 67488
rect 44520 67424 44528 67488
rect 44208 66400 44528 67424
rect 44208 66336 44216 66400
rect 44280 66336 44296 66400
rect 44360 66336 44376 66400
rect 44440 66336 44456 66400
rect 44520 66336 44528 66400
rect 44208 65312 44528 66336
rect 44208 65248 44216 65312
rect 44280 65248 44296 65312
rect 44360 65248 44376 65312
rect 44440 65248 44456 65312
rect 44520 65248 44528 65312
rect 44208 64224 44528 65248
rect 44208 64160 44216 64224
rect 44280 64160 44296 64224
rect 44360 64160 44376 64224
rect 44440 64160 44456 64224
rect 44520 64160 44528 64224
rect 44208 63136 44528 64160
rect 44208 63072 44216 63136
rect 44280 63072 44296 63136
rect 44360 63072 44376 63136
rect 44440 63072 44456 63136
rect 44520 63072 44528 63136
rect 44208 62048 44528 63072
rect 44208 61984 44216 62048
rect 44280 61984 44296 62048
rect 44360 61984 44376 62048
rect 44440 61984 44456 62048
rect 44520 61984 44528 62048
rect 44208 60960 44528 61984
rect 44208 60896 44216 60960
rect 44280 60896 44296 60960
rect 44360 60896 44376 60960
rect 44440 60896 44456 60960
rect 44520 60896 44528 60960
rect 44208 59872 44528 60896
rect 44208 59808 44216 59872
rect 44280 59808 44296 59872
rect 44360 59808 44376 59872
rect 44440 59808 44456 59872
rect 44520 59808 44528 59872
rect 44208 58784 44528 59808
rect 44208 58720 44216 58784
rect 44280 58720 44296 58784
rect 44360 58720 44376 58784
rect 44440 58720 44456 58784
rect 44520 58720 44528 58784
rect 44208 57696 44528 58720
rect 44208 57632 44216 57696
rect 44280 57632 44296 57696
rect 44360 57632 44376 57696
rect 44440 57632 44456 57696
rect 44520 57632 44528 57696
rect 44208 56608 44528 57632
rect 44208 56544 44216 56608
rect 44280 56544 44296 56608
rect 44360 56544 44376 56608
rect 44440 56544 44456 56608
rect 44520 56544 44528 56608
rect 44208 55520 44528 56544
rect 44208 55456 44216 55520
rect 44280 55456 44296 55520
rect 44360 55456 44376 55520
rect 44440 55456 44456 55520
rect 44520 55456 44528 55520
rect 44208 54432 44528 55456
rect 44208 54368 44216 54432
rect 44280 54368 44296 54432
rect 44360 54368 44376 54432
rect 44440 54368 44456 54432
rect 44520 54368 44528 54432
rect 44208 53344 44528 54368
rect 44208 53280 44216 53344
rect 44280 53280 44296 53344
rect 44360 53280 44376 53344
rect 44440 53280 44456 53344
rect 44520 53280 44528 53344
rect 44208 52256 44528 53280
rect 44208 52192 44216 52256
rect 44280 52192 44296 52256
rect 44360 52192 44376 52256
rect 44440 52192 44456 52256
rect 44520 52192 44528 52256
rect 44208 51168 44528 52192
rect 44208 51104 44216 51168
rect 44280 51104 44296 51168
rect 44360 51104 44376 51168
rect 44440 51104 44456 51168
rect 44520 51104 44528 51168
rect 44208 50080 44528 51104
rect 44208 50016 44216 50080
rect 44280 50016 44296 50080
rect 44360 50016 44376 50080
rect 44440 50016 44456 50080
rect 44520 50016 44528 50080
rect 44208 48992 44528 50016
rect 44208 48928 44216 48992
rect 44280 48928 44296 48992
rect 44360 48928 44376 48992
rect 44440 48928 44456 48992
rect 44520 48928 44528 48992
rect 44208 47904 44528 48928
rect 44208 47840 44216 47904
rect 44280 47840 44296 47904
rect 44360 47840 44376 47904
rect 44440 47840 44456 47904
rect 44520 47840 44528 47904
rect 44208 46816 44528 47840
rect 44208 46752 44216 46816
rect 44280 46752 44296 46816
rect 44360 46752 44376 46816
rect 44440 46752 44456 46816
rect 44520 46752 44528 46816
rect 44208 45728 44528 46752
rect 44208 45664 44216 45728
rect 44280 45664 44296 45728
rect 44360 45664 44376 45728
rect 44440 45664 44456 45728
rect 44520 45664 44528 45728
rect 44208 44640 44528 45664
rect 44208 44576 44216 44640
rect 44280 44576 44296 44640
rect 44360 44576 44376 44640
rect 44440 44576 44456 44640
rect 44520 44576 44528 44640
rect 44208 43552 44528 44576
rect 44208 43488 44216 43552
rect 44280 43488 44296 43552
rect 44360 43488 44376 43552
rect 44440 43488 44456 43552
rect 44520 43488 44528 43552
rect 44208 42464 44528 43488
rect 44208 42400 44216 42464
rect 44280 42400 44296 42464
rect 44360 42400 44376 42464
rect 44440 42400 44456 42464
rect 44520 42400 44528 42464
rect 44208 41376 44528 42400
rect 44208 41312 44216 41376
rect 44280 41312 44296 41376
rect 44360 41312 44376 41376
rect 44440 41312 44456 41376
rect 44520 41312 44528 41376
rect 44208 40288 44528 41312
rect 44208 40224 44216 40288
rect 44280 40224 44296 40288
rect 44360 40224 44376 40288
rect 44440 40224 44456 40288
rect 44520 40224 44528 40288
rect 44208 39200 44528 40224
rect 44208 39136 44216 39200
rect 44280 39136 44296 39200
rect 44360 39136 44376 39200
rect 44440 39136 44456 39200
rect 44520 39136 44528 39200
rect 44208 38112 44528 39136
rect 44208 38048 44216 38112
rect 44280 38048 44296 38112
rect 44360 38048 44376 38112
rect 44440 38048 44456 38112
rect 44520 38048 44528 38112
rect 44208 37024 44528 38048
rect 44208 36960 44216 37024
rect 44280 36960 44296 37024
rect 44360 36960 44376 37024
rect 44440 36960 44456 37024
rect 44520 36960 44528 37024
rect 44208 35936 44528 36960
rect 44208 35872 44216 35936
rect 44280 35872 44296 35936
rect 44360 35872 44376 35936
rect 44440 35872 44456 35936
rect 44520 35872 44528 35936
rect 44208 34848 44528 35872
rect 44208 34784 44216 34848
rect 44280 34784 44296 34848
rect 44360 34784 44376 34848
rect 44440 34784 44456 34848
rect 44520 34784 44528 34848
rect 44208 33760 44528 34784
rect 44208 33696 44216 33760
rect 44280 33696 44296 33760
rect 44360 33696 44376 33760
rect 44440 33696 44456 33760
rect 44520 33696 44528 33760
rect 44208 32672 44528 33696
rect 44208 32608 44216 32672
rect 44280 32608 44296 32672
rect 44360 32608 44376 32672
rect 44440 32608 44456 32672
rect 44520 32608 44528 32672
rect 44208 31584 44528 32608
rect 44208 31520 44216 31584
rect 44280 31520 44296 31584
rect 44360 31520 44376 31584
rect 44440 31520 44456 31584
rect 44520 31520 44528 31584
rect 44208 30496 44528 31520
rect 44208 30432 44216 30496
rect 44280 30432 44296 30496
rect 44360 30432 44376 30496
rect 44440 30432 44456 30496
rect 44520 30432 44528 30496
rect 44208 29408 44528 30432
rect 44208 29344 44216 29408
rect 44280 29344 44296 29408
rect 44360 29344 44376 29408
rect 44440 29344 44456 29408
rect 44520 29344 44528 29408
rect 44208 28320 44528 29344
rect 44208 28256 44216 28320
rect 44280 28256 44296 28320
rect 44360 28256 44376 28320
rect 44440 28256 44456 28320
rect 44520 28256 44528 28320
rect 44208 27232 44528 28256
rect 44208 27168 44216 27232
rect 44280 27168 44296 27232
rect 44360 27168 44376 27232
rect 44440 27168 44456 27232
rect 44520 27168 44528 27232
rect 44208 26144 44528 27168
rect 44208 26080 44216 26144
rect 44280 26080 44296 26144
rect 44360 26080 44376 26144
rect 44440 26080 44456 26144
rect 44520 26080 44528 26144
rect 44208 25056 44528 26080
rect 44208 24992 44216 25056
rect 44280 24992 44296 25056
rect 44360 24992 44376 25056
rect 44440 24992 44456 25056
rect 44520 24992 44528 25056
rect 44208 23968 44528 24992
rect 44208 23904 44216 23968
rect 44280 23904 44296 23968
rect 44360 23904 44376 23968
rect 44440 23904 44456 23968
rect 44520 23904 44528 23968
rect 44208 22880 44528 23904
rect 44208 22816 44216 22880
rect 44280 22816 44296 22880
rect 44360 22816 44376 22880
rect 44440 22816 44456 22880
rect 44520 22816 44528 22880
rect 44208 21792 44528 22816
rect 44208 21728 44216 21792
rect 44280 21728 44296 21792
rect 44360 21728 44376 21792
rect 44440 21728 44456 21792
rect 44520 21728 44528 21792
rect 44208 20704 44528 21728
rect 44208 20640 44216 20704
rect 44280 20640 44296 20704
rect 44360 20640 44376 20704
rect 44440 20640 44456 20704
rect 44520 20640 44528 20704
rect 44208 19616 44528 20640
rect 44208 19552 44216 19616
rect 44280 19552 44296 19616
rect 44360 19552 44376 19616
rect 44440 19552 44456 19616
rect 44520 19552 44528 19616
rect 44208 18528 44528 19552
rect 44208 18464 44216 18528
rect 44280 18464 44296 18528
rect 44360 18464 44376 18528
rect 44440 18464 44456 18528
rect 44520 18464 44528 18528
rect 44208 17440 44528 18464
rect 44208 17376 44216 17440
rect 44280 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44528 17440
rect 39803 17236 39869 17237
rect 39803 17172 39804 17236
rect 39868 17172 39869 17236
rect 39803 17171 39869 17172
rect 39208 16832 39216 16896
rect 39280 16832 39296 16896
rect 39360 16832 39376 16896
rect 39440 16832 39456 16896
rect 39520 16832 39528 16896
rect 39208 15808 39528 16832
rect 39208 15744 39216 15808
rect 39280 15744 39296 15808
rect 39360 15744 39376 15808
rect 39440 15744 39456 15808
rect 39520 15744 39528 15808
rect 39208 14720 39528 15744
rect 39208 14656 39216 14720
rect 39280 14656 39296 14720
rect 39360 14656 39376 14720
rect 39440 14656 39456 14720
rect 39520 14656 39528 14720
rect 39208 13632 39528 14656
rect 39208 13568 39216 13632
rect 39280 13568 39296 13632
rect 39360 13568 39376 13632
rect 39440 13568 39456 13632
rect 39520 13568 39528 13632
rect 39067 13156 39133 13157
rect 39067 13092 39068 13156
rect 39132 13092 39133 13156
rect 39067 13091 39133 13092
rect 38699 12204 38765 12205
rect 38699 12140 38700 12204
rect 38764 12140 38765 12204
rect 38699 12139 38765 12140
rect 34208 11843 34216 11907
rect 34280 11843 34296 11907
rect 34360 11843 34376 11907
rect 34440 11843 34456 11907
rect 34520 11843 34528 11907
rect 34208 11827 34528 11843
rect 34208 11763 34216 11827
rect 34280 11763 34296 11827
rect 34360 11763 34376 11827
rect 34440 11763 34456 11827
rect 34520 11763 34528 11827
rect 34208 11747 34528 11763
rect 34208 11683 34216 11747
rect 34280 11683 34296 11747
rect 34360 11683 34376 11747
rect 34440 11683 34456 11747
rect 34520 11683 34528 11747
rect 34208 11667 34528 11683
rect 34208 11603 34216 11667
rect 34280 11603 34296 11667
rect 34360 11603 34376 11667
rect 34440 11603 34456 11667
rect 34520 11603 34528 11667
rect 34208 9358 34528 11603
rect 38883 9484 38949 9485
rect 38883 9420 38884 9484
rect 38948 9420 38949 9484
rect 38883 9419 38949 9420
rect 34208 9294 34216 9358
rect 34280 9294 34296 9358
rect 34360 9294 34376 9358
rect 34440 9294 34456 9358
rect 34520 9294 34528 9358
rect 34208 9278 34528 9294
rect 34208 9214 34216 9278
rect 34280 9214 34296 9278
rect 34360 9214 34376 9278
rect 34440 9214 34456 9278
rect 34520 9214 34528 9278
rect 34208 9198 34528 9214
rect 34208 9134 34216 9198
rect 34280 9134 34296 9198
rect 34360 9134 34376 9198
rect 34440 9134 34456 9198
rect 34520 9134 34528 9198
rect 34208 9118 34528 9134
rect 34208 9054 34216 9118
rect 34280 9054 34296 9118
rect 34360 9054 34376 9118
rect 34440 9054 34456 9118
rect 34520 9054 34528 9118
rect 34208 6809 34528 9054
rect 38886 7445 38946 9419
rect 38883 7444 38949 7445
rect 38883 7380 38884 7444
rect 38948 7380 38949 7444
rect 38883 7379 38949 7380
rect 34208 6745 34216 6809
rect 34280 6745 34296 6809
rect 34360 6745 34376 6809
rect 34440 6745 34456 6809
rect 34520 6745 34528 6809
rect 34208 6729 34528 6745
rect 34208 6665 34216 6729
rect 34280 6665 34296 6729
rect 34360 6665 34376 6729
rect 34440 6665 34456 6729
rect 34520 6665 34528 6729
rect 34208 6649 34528 6665
rect 34208 6585 34216 6649
rect 34280 6585 34296 6649
rect 34360 6585 34376 6649
rect 34440 6585 34456 6649
rect 34520 6585 34528 6649
rect 34208 6569 34528 6585
rect 34208 6505 34216 6569
rect 34280 6505 34296 6569
rect 34360 6505 34376 6569
rect 34440 6505 34456 6569
rect 34520 6505 34528 6569
rect 30419 6084 30485 6085
rect 30419 6020 30420 6084
rect 30484 6020 30485 6084
rect 30419 6019 30485 6020
rect 30051 5268 30117 5269
rect 30051 5204 30052 5268
rect 30116 5204 30117 5268
rect 30051 5203 30117 5204
rect 29208 2366 29216 2430
rect 29280 2366 29296 2430
rect 29360 2366 29376 2430
rect 29440 2366 29456 2430
rect 29520 2366 29528 2430
rect 29208 2350 29528 2366
rect 29208 2286 29216 2350
rect 29280 2286 29296 2350
rect 29360 2286 29376 2350
rect 29440 2286 29456 2350
rect 29520 2286 29528 2350
rect 29208 2270 29528 2286
rect 29208 2206 29216 2270
rect 29280 2206 29296 2270
rect 29360 2206 29376 2270
rect 29440 2206 29456 2270
rect 29520 2206 29528 2270
rect 29208 2176 29528 2206
rect 30054 1869 30114 5203
rect 30422 1869 30482 6019
rect 30603 5540 30669 5541
rect 30603 5476 30604 5540
rect 30668 5476 30669 5540
rect 30603 5475 30669 5476
rect 30051 1868 30117 1869
rect 30051 1804 30052 1868
rect 30116 1804 30117 1868
rect 30051 1803 30117 1804
rect 30419 1868 30485 1869
rect 30419 1804 30420 1868
rect 30484 1804 30485 1868
rect 30419 1803 30485 1804
rect 30606 1733 30666 5475
rect 31891 5404 31957 5405
rect 31891 5340 31892 5404
rect 31956 5340 31957 5404
rect 31891 5339 31957 5340
rect 31155 4724 31221 4725
rect 31155 4660 31156 4724
rect 31220 4660 31221 4724
rect 31155 4659 31221 4660
rect 31158 1869 31218 4659
rect 31155 1868 31221 1869
rect 31155 1804 31156 1868
rect 31220 1804 31221 1868
rect 31155 1803 31221 1804
rect 28211 1732 28277 1733
rect 28211 1668 28212 1732
rect 28276 1668 28277 1732
rect 28211 1667 28277 1668
rect 30603 1732 30669 1733
rect 30603 1668 30604 1732
rect 30668 1668 30669 1732
rect 30603 1667 30669 1668
rect 31894 1189 31954 5339
rect 33731 3772 33797 3773
rect 33731 3708 33732 3772
rect 33796 3770 33797 3772
rect 33796 3710 33978 3770
rect 33796 3708 33797 3710
rect 33731 3707 33797 3708
rect 33918 2957 33978 3710
rect 33915 2956 33981 2957
rect 33915 2892 33916 2956
rect 33980 2892 33981 2956
rect 33915 2891 33981 2892
rect 34208 2176 34528 6505
rect 38883 4452 38949 4453
rect 38883 4388 38884 4452
rect 38948 4388 38949 4452
rect 38883 4387 38949 4388
rect 38886 3909 38946 4387
rect 38883 3908 38949 3909
rect 38883 3844 38884 3908
rect 38948 3844 38949 3908
rect 38883 3843 38949 3844
rect 39070 3365 39130 13091
rect 39208 12544 39528 13568
rect 39806 13021 39866 17171
rect 44208 16352 44528 17376
rect 44208 16288 44216 16352
rect 44280 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44528 16352
rect 44208 15264 44528 16288
rect 44208 15200 44216 15264
rect 44280 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44528 15264
rect 40171 14516 40237 14517
rect 40171 14452 40172 14516
rect 40236 14452 40237 14516
rect 40171 14451 40237 14452
rect 39803 13020 39869 13021
rect 39803 12956 39804 13020
rect 39868 12956 39869 13020
rect 39803 12955 39869 12956
rect 39208 12480 39216 12544
rect 39280 12480 39296 12544
rect 39360 12480 39376 12544
rect 39440 12480 39456 12544
rect 39520 12480 39528 12544
rect 39208 11456 39528 12480
rect 39619 12476 39685 12477
rect 39619 12412 39620 12476
rect 39684 12412 39685 12476
rect 39619 12411 39685 12412
rect 39208 11392 39216 11456
rect 39280 11392 39296 11456
rect 39360 11392 39376 11456
rect 39440 11392 39456 11456
rect 39520 11392 39528 11456
rect 39208 10368 39528 11392
rect 39208 10304 39216 10368
rect 39280 10304 39296 10368
rect 39360 10304 39376 10368
rect 39440 10304 39456 10368
rect 39520 10304 39528 10368
rect 39208 9280 39528 10304
rect 39208 9216 39216 9280
rect 39280 9216 39296 9280
rect 39360 9216 39376 9280
rect 39440 9216 39456 9280
rect 39520 9216 39528 9280
rect 39208 8192 39528 9216
rect 39208 8128 39216 8192
rect 39280 8128 39296 8192
rect 39360 8128 39376 8192
rect 39440 8128 39456 8192
rect 39520 8128 39528 8192
rect 39208 7104 39528 8128
rect 39208 7040 39216 7104
rect 39280 7040 39296 7104
rect 39360 7040 39376 7104
rect 39440 7040 39456 7104
rect 39520 7040 39528 7104
rect 39208 6016 39528 7040
rect 39622 7037 39682 12411
rect 39803 12204 39869 12205
rect 39803 12140 39804 12204
rect 39868 12140 39869 12204
rect 39803 12139 39869 12140
rect 39619 7036 39685 7037
rect 39619 6972 39620 7036
rect 39684 6972 39685 7036
rect 39619 6971 39685 6972
rect 39208 5952 39216 6016
rect 39280 5952 39296 6016
rect 39360 5952 39376 6016
rect 39440 5952 39456 6016
rect 39520 5952 39528 6016
rect 39208 4928 39528 5952
rect 39208 4864 39216 4928
rect 39280 4864 39296 4928
rect 39360 4864 39376 4928
rect 39440 4864 39456 4928
rect 39520 4864 39528 4928
rect 39208 3840 39528 4864
rect 39208 3776 39216 3840
rect 39280 3776 39296 3840
rect 39360 3776 39376 3840
rect 39440 3776 39456 3840
rect 39520 3776 39528 3840
rect 39067 3364 39133 3365
rect 39067 3300 39068 3364
rect 39132 3300 39133 3364
rect 39067 3299 39133 3300
rect 39208 2752 39528 3776
rect 39806 3365 39866 12139
rect 40174 9077 40234 14451
rect 44208 14176 44528 15200
rect 44208 14112 44216 14176
rect 44280 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44528 14176
rect 44208 13088 44528 14112
rect 44208 13024 44216 13088
rect 44280 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44528 13088
rect 40723 12612 40789 12613
rect 40723 12548 40724 12612
rect 40788 12548 40789 12612
rect 40723 12547 40789 12548
rect 40355 10572 40421 10573
rect 40355 10508 40356 10572
rect 40420 10508 40421 10572
rect 40355 10507 40421 10508
rect 40171 9076 40237 9077
rect 40171 9012 40172 9076
rect 40236 9012 40237 9076
rect 40171 9011 40237 9012
rect 39987 8940 40053 8941
rect 39987 8876 39988 8940
rect 40052 8876 40053 8940
rect 39987 8875 40053 8876
rect 39990 4589 40050 8875
rect 40358 8533 40418 10507
rect 40355 8532 40421 8533
rect 40355 8468 40356 8532
rect 40420 8468 40421 8532
rect 40355 8467 40421 8468
rect 39987 4588 40053 4589
rect 39987 4524 39988 4588
rect 40052 4524 40053 4588
rect 39987 4523 40053 4524
rect 39803 3364 39869 3365
rect 39803 3300 39804 3364
rect 39868 3300 39869 3364
rect 39803 3299 39869 3300
rect 40726 3093 40786 12547
rect 44208 12000 44528 13024
rect 44208 11936 44216 12000
rect 44280 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44528 12000
rect 42563 11116 42629 11117
rect 42563 11052 42564 11116
rect 42628 11052 42629 11116
rect 42563 11051 42629 11052
rect 40907 9212 40973 9213
rect 40907 9148 40908 9212
rect 40972 9148 40973 9212
rect 40907 9147 40973 9148
rect 40910 4725 40970 9147
rect 41459 9076 41525 9077
rect 41459 9012 41460 9076
rect 41524 9012 41525 9076
rect 41459 9011 41525 9012
rect 41275 8260 41341 8261
rect 41275 8196 41276 8260
rect 41340 8196 41341 8260
rect 41275 8195 41341 8196
rect 40907 4724 40973 4725
rect 40907 4660 40908 4724
rect 40972 4660 40973 4724
rect 40907 4659 40973 4660
rect 40723 3092 40789 3093
rect 40723 3028 40724 3092
rect 40788 3028 40789 3092
rect 40723 3027 40789 3028
rect 39208 2688 39216 2752
rect 39280 2688 39296 2752
rect 39360 2688 39376 2752
rect 39440 2688 39456 2752
rect 39520 2688 39528 2752
rect 39208 2128 39528 2688
rect 41278 1325 41338 8195
rect 41462 3093 41522 9011
rect 42379 8940 42445 8941
rect 42379 8876 42380 8940
rect 42444 8876 42445 8940
rect 42379 8875 42445 8876
rect 42011 6084 42077 6085
rect 42011 6020 42012 6084
rect 42076 6020 42077 6084
rect 42011 6019 42077 6020
rect 41459 3092 41525 3093
rect 41459 3028 41460 3092
rect 41524 3028 41525 3092
rect 41459 3027 41525 3028
rect 42014 2277 42074 6019
rect 42382 3093 42442 8875
rect 42379 3092 42445 3093
rect 42379 3028 42380 3092
rect 42444 3028 42445 3092
rect 42379 3027 42445 3028
rect 42566 2685 42626 11051
rect 44208 10912 44528 11936
rect 44208 10848 44216 10912
rect 44280 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44528 10912
rect 44208 9824 44528 10848
rect 44208 9760 44216 9824
rect 44280 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44528 9824
rect 43851 9484 43917 9485
rect 43851 9420 43852 9484
rect 43916 9420 43917 9484
rect 43851 9419 43917 9420
rect 43854 3093 43914 9419
rect 44035 8940 44101 8941
rect 44035 8876 44036 8940
rect 44100 8876 44101 8940
rect 44035 8875 44101 8876
rect 44038 3773 44098 8875
rect 44208 8736 44528 9760
rect 44208 8672 44216 8736
rect 44280 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44528 8736
rect 44208 7648 44528 8672
rect 49208 66944 49528 67504
rect 49208 66880 49216 66944
rect 49280 66880 49296 66944
rect 49360 66880 49376 66944
rect 49440 66880 49456 66944
rect 49520 66880 49528 66944
rect 49208 65856 49528 66880
rect 49208 65792 49216 65856
rect 49280 65792 49296 65856
rect 49360 65792 49376 65856
rect 49440 65792 49456 65856
rect 49520 65792 49528 65856
rect 49208 64768 49528 65792
rect 49208 64704 49216 64768
rect 49280 64704 49296 64768
rect 49360 64704 49376 64768
rect 49440 64704 49456 64768
rect 49520 64704 49528 64768
rect 49208 63680 49528 64704
rect 49208 63616 49216 63680
rect 49280 63616 49296 63680
rect 49360 63616 49376 63680
rect 49440 63616 49456 63680
rect 49520 63616 49528 63680
rect 49208 62592 49528 63616
rect 49208 62528 49216 62592
rect 49280 62528 49296 62592
rect 49360 62528 49376 62592
rect 49440 62528 49456 62592
rect 49520 62528 49528 62592
rect 49208 61504 49528 62528
rect 49208 61440 49216 61504
rect 49280 61440 49296 61504
rect 49360 61440 49376 61504
rect 49440 61440 49456 61504
rect 49520 61440 49528 61504
rect 49208 60416 49528 61440
rect 49208 60352 49216 60416
rect 49280 60352 49296 60416
rect 49360 60352 49376 60416
rect 49440 60352 49456 60416
rect 49520 60352 49528 60416
rect 49208 59328 49528 60352
rect 49208 59264 49216 59328
rect 49280 59264 49296 59328
rect 49360 59264 49376 59328
rect 49440 59264 49456 59328
rect 49520 59264 49528 59328
rect 49208 58240 49528 59264
rect 49208 58176 49216 58240
rect 49280 58176 49296 58240
rect 49360 58176 49376 58240
rect 49440 58176 49456 58240
rect 49520 58176 49528 58240
rect 49208 57152 49528 58176
rect 49208 57088 49216 57152
rect 49280 57088 49296 57152
rect 49360 57088 49376 57152
rect 49440 57088 49456 57152
rect 49520 57088 49528 57152
rect 49208 56064 49528 57088
rect 49208 56000 49216 56064
rect 49280 56000 49296 56064
rect 49360 56000 49376 56064
rect 49440 56000 49456 56064
rect 49520 56000 49528 56064
rect 49208 54976 49528 56000
rect 49208 54912 49216 54976
rect 49280 54912 49296 54976
rect 49360 54912 49376 54976
rect 49440 54912 49456 54976
rect 49520 54912 49528 54976
rect 49208 53888 49528 54912
rect 49208 53824 49216 53888
rect 49280 53824 49296 53888
rect 49360 53824 49376 53888
rect 49440 53824 49456 53888
rect 49520 53824 49528 53888
rect 49208 52800 49528 53824
rect 49208 52736 49216 52800
rect 49280 52736 49296 52800
rect 49360 52736 49376 52800
rect 49440 52736 49456 52800
rect 49520 52736 49528 52800
rect 49208 51712 49528 52736
rect 49208 51648 49216 51712
rect 49280 51648 49296 51712
rect 49360 51648 49376 51712
rect 49440 51648 49456 51712
rect 49520 51648 49528 51712
rect 49208 50624 49528 51648
rect 49208 50560 49216 50624
rect 49280 50560 49296 50624
rect 49360 50560 49376 50624
rect 49440 50560 49456 50624
rect 49520 50560 49528 50624
rect 49208 49536 49528 50560
rect 49208 49472 49216 49536
rect 49280 49472 49296 49536
rect 49360 49472 49376 49536
rect 49440 49472 49456 49536
rect 49520 49472 49528 49536
rect 49208 48448 49528 49472
rect 49208 48384 49216 48448
rect 49280 48384 49296 48448
rect 49360 48384 49376 48448
rect 49440 48384 49456 48448
rect 49520 48384 49528 48448
rect 49208 47360 49528 48384
rect 49208 47296 49216 47360
rect 49280 47296 49296 47360
rect 49360 47296 49376 47360
rect 49440 47296 49456 47360
rect 49520 47296 49528 47360
rect 49208 46272 49528 47296
rect 49208 46208 49216 46272
rect 49280 46208 49296 46272
rect 49360 46208 49376 46272
rect 49440 46208 49456 46272
rect 49520 46208 49528 46272
rect 49208 45184 49528 46208
rect 49208 45120 49216 45184
rect 49280 45120 49296 45184
rect 49360 45120 49376 45184
rect 49440 45120 49456 45184
rect 49520 45120 49528 45184
rect 49208 44096 49528 45120
rect 49208 44032 49216 44096
rect 49280 44032 49296 44096
rect 49360 44032 49376 44096
rect 49440 44032 49456 44096
rect 49520 44032 49528 44096
rect 49208 43008 49528 44032
rect 49208 42944 49216 43008
rect 49280 42944 49296 43008
rect 49360 42944 49376 43008
rect 49440 42944 49456 43008
rect 49520 42944 49528 43008
rect 49208 41920 49528 42944
rect 49208 41856 49216 41920
rect 49280 41856 49296 41920
rect 49360 41856 49376 41920
rect 49440 41856 49456 41920
rect 49520 41856 49528 41920
rect 49208 40832 49528 41856
rect 49208 40768 49216 40832
rect 49280 40768 49296 40832
rect 49360 40768 49376 40832
rect 49440 40768 49456 40832
rect 49520 40768 49528 40832
rect 49208 39744 49528 40768
rect 49208 39680 49216 39744
rect 49280 39680 49296 39744
rect 49360 39680 49376 39744
rect 49440 39680 49456 39744
rect 49520 39680 49528 39744
rect 49208 38656 49528 39680
rect 49208 38592 49216 38656
rect 49280 38592 49296 38656
rect 49360 38592 49376 38656
rect 49440 38592 49456 38656
rect 49520 38592 49528 38656
rect 49208 37568 49528 38592
rect 49208 37504 49216 37568
rect 49280 37504 49296 37568
rect 49360 37504 49376 37568
rect 49440 37504 49456 37568
rect 49520 37504 49528 37568
rect 49208 36480 49528 37504
rect 49208 36416 49216 36480
rect 49280 36416 49296 36480
rect 49360 36416 49376 36480
rect 49440 36416 49456 36480
rect 49520 36416 49528 36480
rect 49208 35392 49528 36416
rect 49208 35328 49216 35392
rect 49280 35328 49296 35392
rect 49360 35328 49376 35392
rect 49440 35328 49456 35392
rect 49520 35328 49528 35392
rect 49208 34304 49528 35328
rect 49208 34240 49216 34304
rect 49280 34240 49296 34304
rect 49360 34240 49376 34304
rect 49440 34240 49456 34304
rect 49520 34240 49528 34304
rect 49208 33216 49528 34240
rect 49208 33152 49216 33216
rect 49280 33152 49296 33216
rect 49360 33152 49376 33216
rect 49440 33152 49456 33216
rect 49520 33152 49528 33216
rect 49208 32128 49528 33152
rect 49208 32064 49216 32128
rect 49280 32064 49296 32128
rect 49360 32064 49376 32128
rect 49440 32064 49456 32128
rect 49520 32064 49528 32128
rect 49208 31040 49528 32064
rect 49208 30976 49216 31040
rect 49280 30976 49296 31040
rect 49360 30976 49376 31040
rect 49440 30976 49456 31040
rect 49520 30976 49528 31040
rect 49208 29952 49528 30976
rect 49208 29888 49216 29952
rect 49280 29888 49296 29952
rect 49360 29888 49376 29952
rect 49440 29888 49456 29952
rect 49520 29888 49528 29952
rect 49208 28864 49528 29888
rect 49208 28800 49216 28864
rect 49280 28800 49296 28864
rect 49360 28800 49376 28864
rect 49440 28800 49456 28864
rect 49520 28800 49528 28864
rect 49208 27776 49528 28800
rect 49208 27712 49216 27776
rect 49280 27712 49296 27776
rect 49360 27712 49376 27776
rect 49440 27712 49456 27776
rect 49520 27712 49528 27776
rect 49208 26688 49528 27712
rect 49208 26624 49216 26688
rect 49280 26624 49296 26688
rect 49360 26624 49376 26688
rect 49440 26624 49456 26688
rect 49520 26624 49528 26688
rect 49208 25600 49528 26624
rect 49208 25536 49216 25600
rect 49280 25536 49296 25600
rect 49360 25536 49376 25600
rect 49440 25536 49456 25600
rect 49520 25536 49528 25600
rect 49208 24512 49528 25536
rect 49208 24448 49216 24512
rect 49280 24448 49296 24512
rect 49360 24448 49376 24512
rect 49440 24448 49456 24512
rect 49520 24448 49528 24512
rect 49208 23424 49528 24448
rect 49208 23360 49216 23424
rect 49280 23360 49296 23424
rect 49360 23360 49376 23424
rect 49440 23360 49456 23424
rect 49520 23360 49528 23424
rect 49208 22336 49528 23360
rect 49208 22272 49216 22336
rect 49280 22272 49296 22336
rect 49360 22272 49376 22336
rect 49440 22272 49456 22336
rect 49520 22272 49528 22336
rect 49208 21248 49528 22272
rect 49208 21184 49216 21248
rect 49280 21184 49296 21248
rect 49360 21184 49376 21248
rect 49440 21184 49456 21248
rect 49520 21184 49528 21248
rect 49208 20160 49528 21184
rect 49208 20096 49216 20160
rect 49280 20096 49296 20160
rect 49360 20096 49376 20160
rect 49440 20096 49456 20160
rect 49520 20096 49528 20160
rect 49208 19072 49528 20096
rect 49208 19008 49216 19072
rect 49280 19008 49296 19072
rect 49360 19008 49376 19072
rect 49440 19008 49456 19072
rect 49520 19008 49528 19072
rect 49208 17984 49528 19008
rect 49208 17920 49216 17984
rect 49280 17920 49296 17984
rect 49360 17920 49376 17984
rect 49440 17920 49456 17984
rect 49520 17920 49528 17984
rect 49208 16896 49528 17920
rect 49208 16832 49216 16896
rect 49280 16832 49296 16896
rect 49360 16832 49376 16896
rect 49440 16832 49456 16896
rect 49520 16832 49528 16896
rect 49208 15808 49528 16832
rect 49208 15744 49216 15808
rect 49280 15744 49296 15808
rect 49360 15744 49376 15808
rect 49440 15744 49456 15808
rect 49520 15744 49528 15808
rect 49208 14720 49528 15744
rect 49208 14656 49216 14720
rect 49280 14656 49296 14720
rect 49360 14656 49376 14720
rect 49440 14656 49456 14720
rect 49520 14656 49528 14720
rect 49208 13632 49528 14656
rect 49208 13568 49216 13632
rect 49280 13568 49296 13632
rect 49360 13568 49376 13632
rect 49440 13568 49456 13632
rect 49520 13568 49528 13632
rect 49208 12544 49528 13568
rect 49208 12480 49216 12544
rect 49280 12480 49296 12544
rect 49360 12480 49376 12544
rect 49440 12480 49456 12544
rect 49520 12480 49528 12544
rect 49208 11456 49528 12480
rect 49208 11392 49216 11456
rect 49280 11392 49296 11456
rect 49360 11392 49376 11456
rect 49440 11392 49456 11456
rect 49520 11392 49528 11456
rect 49208 10368 49528 11392
rect 49208 10304 49216 10368
rect 49280 10304 49296 10368
rect 49360 10304 49376 10368
rect 49440 10304 49456 10368
rect 49520 10304 49528 10368
rect 49208 9280 49528 10304
rect 49208 9216 49216 9280
rect 49280 9216 49296 9280
rect 49360 9216 49376 9280
rect 49440 9216 49456 9280
rect 49520 9216 49528 9280
rect 44955 8532 45021 8533
rect 44955 8468 44956 8532
rect 45020 8468 45021 8532
rect 44955 8467 45021 8468
rect 44208 7584 44216 7648
rect 44280 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44528 7648
rect 44208 6560 44528 7584
rect 44208 6496 44216 6560
rect 44280 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44528 6560
rect 44208 5472 44528 6496
rect 44208 5408 44216 5472
rect 44280 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44528 5472
rect 44208 4384 44528 5408
rect 44208 4320 44216 4384
rect 44280 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44528 4384
rect 44035 3772 44101 3773
rect 44035 3708 44036 3772
rect 44100 3708 44101 3772
rect 44035 3707 44101 3708
rect 44208 3296 44528 4320
rect 44208 3232 44216 3296
rect 44280 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44528 3296
rect 43851 3092 43917 3093
rect 43851 3028 43852 3092
rect 43916 3028 43917 3092
rect 43851 3027 43917 3028
rect 42563 2684 42629 2685
rect 42563 2620 42564 2684
rect 42628 2620 42629 2684
rect 42563 2619 42629 2620
rect 42011 2276 42077 2277
rect 42011 2212 42012 2276
rect 42076 2212 42077 2276
rect 42011 2211 42077 2212
rect 44208 2208 44528 3232
rect 44958 2821 45018 8467
rect 49208 8192 49528 9216
rect 49208 8128 49216 8192
rect 49280 8128 49296 8192
rect 49360 8128 49376 8192
rect 49440 8128 49456 8192
rect 49520 8128 49528 8192
rect 46795 7852 46861 7853
rect 46795 7788 46796 7852
rect 46860 7788 46861 7852
rect 46795 7787 46861 7788
rect 46611 5812 46677 5813
rect 46611 5748 46612 5812
rect 46676 5748 46677 5812
rect 46611 5747 46677 5748
rect 44955 2820 45021 2821
rect 44955 2756 44956 2820
rect 45020 2756 45021 2820
rect 44955 2755 45021 2756
rect 44208 2144 44216 2208
rect 44280 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44528 2208
rect 44208 2128 44528 2144
rect 46614 2005 46674 5747
rect 46798 3365 46858 7787
rect 49208 7104 49528 8128
rect 49208 7040 49216 7104
rect 49280 7040 49296 7104
rect 49360 7040 49376 7104
rect 49440 7040 49456 7104
rect 49520 7040 49528 7104
rect 49208 6016 49528 7040
rect 49208 5952 49216 6016
rect 49280 5952 49296 6016
rect 49360 5952 49376 6016
rect 49440 5952 49456 6016
rect 49520 5952 49528 6016
rect 49208 4928 49528 5952
rect 54208 67488 54528 67504
rect 54208 67424 54216 67488
rect 54280 67424 54296 67488
rect 54360 67424 54376 67488
rect 54440 67424 54456 67488
rect 54520 67424 54528 67488
rect 54208 66400 54528 67424
rect 54208 66336 54216 66400
rect 54280 66336 54296 66400
rect 54360 66336 54376 66400
rect 54440 66336 54456 66400
rect 54520 66336 54528 66400
rect 54208 65312 54528 66336
rect 54208 65248 54216 65312
rect 54280 65248 54296 65312
rect 54360 65248 54376 65312
rect 54440 65248 54456 65312
rect 54520 65248 54528 65312
rect 54208 64224 54528 65248
rect 54208 64160 54216 64224
rect 54280 64160 54296 64224
rect 54360 64160 54376 64224
rect 54440 64160 54456 64224
rect 54520 64160 54528 64224
rect 54208 63136 54528 64160
rect 54208 63072 54216 63136
rect 54280 63072 54296 63136
rect 54360 63072 54376 63136
rect 54440 63072 54456 63136
rect 54520 63072 54528 63136
rect 54208 62048 54528 63072
rect 54208 61984 54216 62048
rect 54280 61984 54296 62048
rect 54360 61984 54376 62048
rect 54440 61984 54456 62048
rect 54520 61984 54528 62048
rect 54208 60960 54528 61984
rect 54208 60896 54216 60960
rect 54280 60896 54296 60960
rect 54360 60896 54376 60960
rect 54440 60896 54456 60960
rect 54520 60896 54528 60960
rect 54208 59872 54528 60896
rect 54208 59808 54216 59872
rect 54280 59808 54296 59872
rect 54360 59808 54376 59872
rect 54440 59808 54456 59872
rect 54520 59808 54528 59872
rect 54208 58784 54528 59808
rect 54208 58720 54216 58784
rect 54280 58720 54296 58784
rect 54360 58720 54376 58784
rect 54440 58720 54456 58784
rect 54520 58720 54528 58784
rect 54208 57696 54528 58720
rect 54208 57632 54216 57696
rect 54280 57632 54296 57696
rect 54360 57632 54376 57696
rect 54440 57632 54456 57696
rect 54520 57632 54528 57696
rect 54208 56608 54528 57632
rect 54208 56544 54216 56608
rect 54280 56544 54296 56608
rect 54360 56544 54376 56608
rect 54440 56544 54456 56608
rect 54520 56544 54528 56608
rect 54208 55520 54528 56544
rect 54208 55456 54216 55520
rect 54280 55456 54296 55520
rect 54360 55456 54376 55520
rect 54440 55456 54456 55520
rect 54520 55456 54528 55520
rect 54208 54432 54528 55456
rect 54208 54368 54216 54432
rect 54280 54368 54296 54432
rect 54360 54368 54376 54432
rect 54440 54368 54456 54432
rect 54520 54368 54528 54432
rect 54208 53344 54528 54368
rect 54208 53280 54216 53344
rect 54280 53280 54296 53344
rect 54360 53280 54376 53344
rect 54440 53280 54456 53344
rect 54520 53280 54528 53344
rect 54208 52256 54528 53280
rect 54208 52192 54216 52256
rect 54280 52192 54296 52256
rect 54360 52192 54376 52256
rect 54440 52192 54456 52256
rect 54520 52192 54528 52256
rect 54208 51168 54528 52192
rect 54208 51104 54216 51168
rect 54280 51104 54296 51168
rect 54360 51104 54376 51168
rect 54440 51104 54456 51168
rect 54520 51104 54528 51168
rect 54208 50080 54528 51104
rect 54208 50016 54216 50080
rect 54280 50016 54296 50080
rect 54360 50016 54376 50080
rect 54440 50016 54456 50080
rect 54520 50016 54528 50080
rect 54208 48992 54528 50016
rect 54208 48928 54216 48992
rect 54280 48928 54296 48992
rect 54360 48928 54376 48992
rect 54440 48928 54456 48992
rect 54520 48928 54528 48992
rect 54208 47904 54528 48928
rect 54208 47840 54216 47904
rect 54280 47840 54296 47904
rect 54360 47840 54376 47904
rect 54440 47840 54456 47904
rect 54520 47840 54528 47904
rect 54208 46816 54528 47840
rect 54208 46752 54216 46816
rect 54280 46752 54296 46816
rect 54360 46752 54376 46816
rect 54440 46752 54456 46816
rect 54520 46752 54528 46816
rect 54208 45728 54528 46752
rect 54208 45664 54216 45728
rect 54280 45664 54296 45728
rect 54360 45664 54376 45728
rect 54440 45664 54456 45728
rect 54520 45664 54528 45728
rect 54208 44640 54528 45664
rect 54208 44576 54216 44640
rect 54280 44576 54296 44640
rect 54360 44576 54376 44640
rect 54440 44576 54456 44640
rect 54520 44576 54528 44640
rect 54208 43552 54528 44576
rect 54208 43488 54216 43552
rect 54280 43488 54296 43552
rect 54360 43488 54376 43552
rect 54440 43488 54456 43552
rect 54520 43488 54528 43552
rect 54208 42464 54528 43488
rect 54208 42400 54216 42464
rect 54280 42400 54296 42464
rect 54360 42400 54376 42464
rect 54440 42400 54456 42464
rect 54520 42400 54528 42464
rect 54208 41376 54528 42400
rect 54208 41312 54216 41376
rect 54280 41312 54296 41376
rect 54360 41312 54376 41376
rect 54440 41312 54456 41376
rect 54520 41312 54528 41376
rect 54208 40288 54528 41312
rect 54208 40224 54216 40288
rect 54280 40224 54296 40288
rect 54360 40224 54376 40288
rect 54440 40224 54456 40288
rect 54520 40224 54528 40288
rect 54208 39200 54528 40224
rect 54208 39136 54216 39200
rect 54280 39136 54296 39200
rect 54360 39136 54376 39200
rect 54440 39136 54456 39200
rect 54520 39136 54528 39200
rect 54208 38112 54528 39136
rect 54208 38048 54216 38112
rect 54280 38048 54296 38112
rect 54360 38048 54376 38112
rect 54440 38048 54456 38112
rect 54520 38048 54528 38112
rect 54208 37024 54528 38048
rect 54208 36960 54216 37024
rect 54280 36960 54296 37024
rect 54360 36960 54376 37024
rect 54440 36960 54456 37024
rect 54520 36960 54528 37024
rect 54208 35936 54528 36960
rect 54208 35872 54216 35936
rect 54280 35872 54296 35936
rect 54360 35872 54376 35936
rect 54440 35872 54456 35936
rect 54520 35872 54528 35936
rect 54208 34848 54528 35872
rect 54208 34784 54216 34848
rect 54280 34784 54296 34848
rect 54360 34784 54376 34848
rect 54440 34784 54456 34848
rect 54520 34784 54528 34848
rect 54208 33760 54528 34784
rect 54208 33696 54216 33760
rect 54280 33696 54296 33760
rect 54360 33696 54376 33760
rect 54440 33696 54456 33760
rect 54520 33696 54528 33760
rect 54208 32672 54528 33696
rect 54208 32608 54216 32672
rect 54280 32608 54296 32672
rect 54360 32608 54376 32672
rect 54440 32608 54456 32672
rect 54520 32608 54528 32672
rect 54208 31584 54528 32608
rect 54208 31520 54216 31584
rect 54280 31520 54296 31584
rect 54360 31520 54376 31584
rect 54440 31520 54456 31584
rect 54520 31520 54528 31584
rect 54208 30496 54528 31520
rect 54208 30432 54216 30496
rect 54280 30432 54296 30496
rect 54360 30432 54376 30496
rect 54440 30432 54456 30496
rect 54520 30432 54528 30496
rect 54208 29408 54528 30432
rect 54208 29344 54216 29408
rect 54280 29344 54296 29408
rect 54360 29344 54376 29408
rect 54440 29344 54456 29408
rect 54520 29344 54528 29408
rect 54208 28320 54528 29344
rect 54208 28256 54216 28320
rect 54280 28256 54296 28320
rect 54360 28256 54376 28320
rect 54440 28256 54456 28320
rect 54520 28256 54528 28320
rect 54208 27232 54528 28256
rect 54208 27168 54216 27232
rect 54280 27168 54296 27232
rect 54360 27168 54376 27232
rect 54440 27168 54456 27232
rect 54520 27168 54528 27232
rect 54208 26144 54528 27168
rect 54208 26080 54216 26144
rect 54280 26080 54296 26144
rect 54360 26080 54376 26144
rect 54440 26080 54456 26144
rect 54520 26080 54528 26144
rect 54208 25056 54528 26080
rect 54208 24992 54216 25056
rect 54280 24992 54296 25056
rect 54360 24992 54376 25056
rect 54440 24992 54456 25056
rect 54520 24992 54528 25056
rect 54208 23968 54528 24992
rect 54208 23904 54216 23968
rect 54280 23904 54296 23968
rect 54360 23904 54376 23968
rect 54440 23904 54456 23968
rect 54520 23904 54528 23968
rect 54208 22880 54528 23904
rect 54208 22816 54216 22880
rect 54280 22816 54296 22880
rect 54360 22816 54376 22880
rect 54440 22816 54456 22880
rect 54520 22816 54528 22880
rect 54208 21792 54528 22816
rect 54208 21728 54216 21792
rect 54280 21728 54296 21792
rect 54360 21728 54376 21792
rect 54440 21728 54456 21792
rect 54520 21728 54528 21792
rect 54208 20704 54528 21728
rect 54208 20640 54216 20704
rect 54280 20640 54296 20704
rect 54360 20640 54376 20704
rect 54440 20640 54456 20704
rect 54520 20640 54528 20704
rect 54208 19616 54528 20640
rect 54208 19552 54216 19616
rect 54280 19552 54296 19616
rect 54360 19552 54376 19616
rect 54440 19552 54456 19616
rect 54520 19552 54528 19616
rect 54208 18528 54528 19552
rect 54208 18464 54216 18528
rect 54280 18464 54296 18528
rect 54360 18464 54376 18528
rect 54440 18464 54456 18528
rect 54520 18464 54528 18528
rect 54208 17440 54528 18464
rect 54208 17376 54216 17440
rect 54280 17376 54296 17440
rect 54360 17376 54376 17440
rect 54440 17376 54456 17440
rect 54520 17376 54528 17440
rect 54208 16352 54528 17376
rect 54208 16288 54216 16352
rect 54280 16288 54296 16352
rect 54360 16288 54376 16352
rect 54440 16288 54456 16352
rect 54520 16288 54528 16352
rect 54208 15264 54528 16288
rect 54208 15200 54216 15264
rect 54280 15200 54296 15264
rect 54360 15200 54376 15264
rect 54440 15200 54456 15264
rect 54520 15200 54528 15264
rect 54208 14176 54528 15200
rect 54208 14112 54216 14176
rect 54280 14112 54296 14176
rect 54360 14112 54376 14176
rect 54440 14112 54456 14176
rect 54520 14112 54528 14176
rect 54208 13088 54528 14112
rect 54208 13024 54216 13088
rect 54280 13024 54296 13088
rect 54360 13024 54376 13088
rect 54440 13024 54456 13088
rect 54520 13024 54528 13088
rect 54208 12000 54528 13024
rect 54208 11936 54216 12000
rect 54280 11936 54296 12000
rect 54360 11936 54376 12000
rect 54440 11936 54456 12000
rect 54520 11936 54528 12000
rect 54208 10912 54528 11936
rect 54208 10848 54216 10912
rect 54280 10848 54296 10912
rect 54360 10848 54376 10912
rect 54440 10848 54456 10912
rect 54520 10848 54528 10912
rect 54208 9824 54528 10848
rect 54208 9760 54216 9824
rect 54280 9760 54296 9824
rect 54360 9760 54376 9824
rect 54440 9760 54456 9824
rect 54520 9760 54528 9824
rect 54208 8736 54528 9760
rect 54208 8672 54216 8736
rect 54280 8672 54296 8736
rect 54360 8672 54376 8736
rect 54440 8672 54456 8736
rect 54520 8672 54528 8736
rect 54208 7648 54528 8672
rect 54208 7584 54216 7648
rect 54280 7584 54296 7648
rect 54360 7584 54376 7648
rect 54440 7584 54456 7648
rect 54520 7584 54528 7648
rect 54208 6560 54528 7584
rect 54208 6496 54216 6560
rect 54280 6496 54296 6560
rect 54360 6496 54376 6560
rect 54440 6496 54456 6560
rect 54520 6496 54528 6560
rect 54208 5472 54528 6496
rect 54208 5408 54216 5472
rect 54280 5408 54296 5472
rect 54360 5408 54376 5472
rect 54440 5408 54456 5472
rect 54520 5408 54528 5472
rect 53603 4996 53669 4997
rect 53603 4932 53604 4996
rect 53668 4932 53669 4996
rect 53603 4931 53669 4932
rect 49208 4864 49216 4928
rect 49280 4864 49296 4928
rect 49360 4864 49376 4928
rect 49440 4864 49456 4928
rect 49520 4864 49528 4928
rect 49208 3840 49528 4864
rect 49739 4044 49805 4045
rect 49739 3980 49740 4044
rect 49804 3980 49805 4044
rect 49739 3979 49805 3980
rect 49208 3776 49216 3840
rect 49280 3776 49296 3840
rect 49360 3776 49376 3840
rect 49440 3776 49456 3840
rect 49520 3776 49528 3840
rect 46795 3364 46861 3365
rect 46795 3300 46796 3364
rect 46860 3300 46861 3364
rect 46795 3299 46861 3300
rect 49208 2752 49528 3776
rect 49208 2688 49216 2752
rect 49280 2688 49296 2752
rect 49360 2688 49376 2752
rect 49440 2688 49456 2752
rect 49520 2688 49528 2752
rect 49208 2128 49528 2688
rect 49742 2277 49802 3979
rect 53606 2549 53666 4931
rect 54208 4384 54528 5408
rect 59208 66944 59528 67504
rect 59208 66880 59216 66944
rect 59280 66880 59296 66944
rect 59360 66880 59376 66944
rect 59440 66880 59456 66944
rect 59520 66880 59528 66944
rect 59208 65856 59528 66880
rect 59208 65792 59216 65856
rect 59280 65792 59296 65856
rect 59360 65792 59376 65856
rect 59440 65792 59456 65856
rect 59520 65792 59528 65856
rect 59208 64768 59528 65792
rect 59208 64704 59216 64768
rect 59280 64704 59296 64768
rect 59360 64704 59376 64768
rect 59440 64704 59456 64768
rect 59520 64704 59528 64768
rect 59208 63680 59528 64704
rect 59208 63616 59216 63680
rect 59280 63616 59296 63680
rect 59360 63616 59376 63680
rect 59440 63616 59456 63680
rect 59520 63616 59528 63680
rect 59208 62592 59528 63616
rect 59208 62528 59216 62592
rect 59280 62528 59296 62592
rect 59360 62528 59376 62592
rect 59440 62528 59456 62592
rect 59520 62528 59528 62592
rect 59208 61504 59528 62528
rect 59208 61440 59216 61504
rect 59280 61440 59296 61504
rect 59360 61440 59376 61504
rect 59440 61440 59456 61504
rect 59520 61440 59528 61504
rect 59208 60416 59528 61440
rect 59208 60352 59216 60416
rect 59280 60352 59296 60416
rect 59360 60352 59376 60416
rect 59440 60352 59456 60416
rect 59520 60352 59528 60416
rect 59208 59328 59528 60352
rect 59208 59264 59216 59328
rect 59280 59264 59296 59328
rect 59360 59264 59376 59328
rect 59440 59264 59456 59328
rect 59520 59264 59528 59328
rect 59208 58240 59528 59264
rect 59208 58176 59216 58240
rect 59280 58176 59296 58240
rect 59360 58176 59376 58240
rect 59440 58176 59456 58240
rect 59520 58176 59528 58240
rect 59208 57152 59528 58176
rect 59208 57088 59216 57152
rect 59280 57088 59296 57152
rect 59360 57088 59376 57152
rect 59440 57088 59456 57152
rect 59520 57088 59528 57152
rect 59208 56064 59528 57088
rect 59208 56000 59216 56064
rect 59280 56000 59296 56064
rect 59360 56000 59376 56064
rect 59440 56000 59456 56064
rect 59520 56000 59528 56064
rect 59208 54976 59528 56000
rect 59208 54912 59216 54976
rect 59280 54912 59296 54976
rect 59360 54912 59376 54976
rect 59440 54912 59456 54976
rect 59520 54912 59528 54976
rect 59208 53888 59528 54912
rect 59208 53824 59216 53888
rect 59280 53824 59296 53888
rect 59360 53824 59376 53888
rect 59440 53824 59456 53888
rect 59520 53824 59528 53888
rect 59208 52800 59528 53824
rect 59208 52736 59216 52800
rect 59280 52736 59296 52800
rect 59360 52736 59376 52800
rect 59440 52736 59456 52800
rect 59520 52736 59528 52800
rect 59208 51712 59528 52736
rect 59208 51648 59216 51712
rect 59280 51648 59296 51712
rect 59360 51648 59376 51712
rect 59440 51648 59456 51712
rect 59520 51648 59528 51712
rect 59208 50624 59528 51648
rect 59208 50560 59216 50624
rect 59280 50560 59296 50624
rect 59360 50560 59376 50624
rect 59440 50560 59456 50624
rect 59520 50560 59528 50624
rect 59208 49536 59528 50560
rect 59208 49472 59216 49536
rect 59280 49472 59296 49536
rect 59360 49472 59376 49536
rect 59440 49472 59456 49536
rect 59520 49472 59528 49536
rect 59208 48448 59528 49472
rect 59208 48384 59216 48448
rect 59280 48384 59296 48448
rect 59360 48384 59376 48448
rect 59440 48384 59456 48448
rect 59520 48384 59528 48448
rect 59208 47360 59528 48384
rect 59208 47296 59216 47360
rect 59280 47296 59296 47360
rect 59360 47296 59376 47360
rect 59440 47296 59456 47360
rect 59520 47296 59528 47360
rect 59208 46272 59528 47296
rect 59208 46208 59216 46272
rect 59280 46208 59296 46272
rect 59360 46208 59376 46272
rect 59440 46208 59456 46272
rect 59520 46208 59528 46272
rect 59208 45184 59528 46208
rect 59208 45120 59216 45184
rect 59280 45120 59296 45184
rect 59360 45120 59376 45184
rect 59440 45120 59456 45184
rect 59520 45120 59528 45184
rect 59208 44096 59528 45120
rect 59208 44032 59216 44096
rect 59280 44032 59296 44096
rect 59360 44032 59376 44096
rect 59440 44032 59456 44096
rect 59520 44032 59528 44096
rect 59208 43008 59528 44032
rect 59208 42944 59216 43008
rect 59280 42944 59296 43008
rect 59360 42944 59376 43008
rect 59440 42944 59456 43008
rect 59520 42944 59528 43008
rect 59208 41920 59528 42944
rect 59208 41856 59216 41920
rect 59280 41856 59296 41920
rect 59360 41856 59376 41920
rect 59440 41856 59456 41920
rect 59520 41856 59528 41920
rect 59208 40832 59528 41856
rect 59208 40768 59216 40832
rect 59280 40768 59296 40832
rect 59360 40768 59376 40832
rect 59440 40768 59456 40832
rect 59520 40768 59528 40832
rect 59208 39744 59528 40768
rect 59208 39680 59216 39744
rect 59280 39680 59296 39744
rect 59360 39680 59376 39744
rect 59440 39680 59456 39744
rect 59520 39680 59528 39744
rect 59208 38656 59528 39680
rect 59208 38592 59216 38656
rect 59280 38592 59296 38656
rect 59360 38592 59376 38656
rect 59440 38592 59456 38656
rect 59520 38592 59528 38656
rect 59208 37568 59528 38592
rect 59208 37504 59216 37568
rect 59280 37504 59296 37568
rect 59360 37504 59376 37568
rect 59440 37504 59456 37568
rect 59520 37504 59528 37568
rect 59208 36480 59528 37504
rect 59208 36416 59216 36480
rect 59280 36416 59296 36480
rect 59360 36416 59376 36480
rect 59440 36416 59456 36480
rect 59520 36416 59528 36480
rect 59208 35392 59528 36416
rect 59208 35328 59216 35392
rect 59280 35328 59296 35392
rect 59360 35328 59376 35392
rect 59440 35328 59456 35392
rect 59520 35328 59528 35392
rect 59208 34304 59528 35328
rect 59208 34240 59216 34304
rect 59280 34240 59296 34304
rect 59360 34240 59376 34304
rect 59440 34240 59456 34304
rect 59520 34240 59528 34304
rect 59208 33216 59528 34240
rect 59208 33152 59216 33216
rect 59280 33152 59296 33216
rect 59360 33152 59376 33216
rect 59440 33152 59456 33216
rect 59520 33152 59528 33216
rect 59208 32128 59528 33152
rect 59208 32064 59216 32128
rect 59280 32064 59296 32128
rect 59360 32064 59376 32128
rect 59440 32064 59456 32128
rect 59520 32064 59528 32128
rect 59208 31040 59528 32064
rect 59208 30976 59216 31040
rect 59280 30976 59296 31040
rect 59360 30976 59376 31040
rect 59440 30976 59456 31040
rect 59520 30976 59528 31040
rect 59208 29952 59528 30976
rect 59208 29888 59216 29952
rect 59280 29888 59296 29952
rect 59360 29888 59376 29952
rect 59440 29888 59456 29952
rect 59520 29888 59528 29952
rect 59208 28864 59528 29888
rect 59208 28800 59216 28864
rect 59280 28800 59296 28864
rect 59360 28800 59376 28864
rect 59440 28800 59456 28864
rect 59520 28800 59528 28864
rect 59208 27776 59528 28800
rect 59208 27712 59216 27776
rect 59280 27712 59296 27776
rect 59360 27712 59376 27776
rect 59440 27712 59456 27776
rect 59520 27712 59528 27776
rect 59208 26688 59528 27712
rect 59208 26624 59216 26688
rect 59280 26624 59296 26688
rect 59360 26624 59376 26688
rect 59440 26624 59456 26688
rect 59520 26624 59528 26688
rect 59208 25600 59528 26624
rect 59208 25536 59216 25600
rect 59280 25536 59296 25600
rect 59360 25536 59376 25600
rect 59440 25536 59456 25600
rect 59520 25536 59528 25600
rect 59208 24512 59528 25536
rect 59208 24448 59216 24512
rect 59280 24448 59296 24512
rect 59360 24448 59376 24512
rect 59440 24448 59456 24512
rect 59520 24448 59528 24512
rect 59208 23424 59528 24448
rect 59208 23360 59216 23424
rect 59280 23360 59296 23424
rect 59360 23360 59376 23424
rect 59440 23360 59456 23424
rect 59520 23360 59528 23424
rect 59208 22336 59528 23360
rect 59208 22272 59216 22336
rect 59280 22272 59296 22336
rect 59360 22272 59376 22336
rect 59440 22272 59456 22336
rect 59520 22272 59528 22336
rect 59208 21248 59528 22272
rect 59208 21184 59216 21248
rect 59280 21184 59296 21248
rect 59360 21184 59376 21248
rect 59440 21184 59456 21248
rect 59520 21184 59528 21248
rect 59208 20160 59528 21184
rect 59208 20096 59216 20160
rect 59280 20096 59296 20160
rect 59360 20096 59376 20160
rect 59440 20096 59456 20160
rect 59520 20096 59528 20160
rect 59208 19072 59528 20096
rect 59208 19008 59216 19072
rect 59280 19008 59296 19072
rect 59360 19008 59376 19072
rect 59440 19008 59456 19072
rect 59520 19008 59528 19072
rect 59208 17984 59528 19008
rect 59208 17920 59216 17984
rect 59280 17920 59296 17984
rect 59360 17920 59376 17984
rect 59440 17920 59456 17984
rect 59520 17920 59528 17984
rect 59208 16896 59528 17920
rect 59208 16832 59216 16896
rect 59280 16832 59296 16896
rect 59360 16832 59376 16896
rect 59440 16832 59456 16896
rect 59520 16832 59528 16896
rect 59208 15808 59528 16832
rect 59208 15744 59216 15808
rect 59280 15744 59296 15808
rect 59360 15744 59376 15808
rect 59440 15744 59456 15808
rect 59520 15744 59528 15808
rect 59208 14720 59528 15744
rect 59208 14656 59216 14720
rect 59280 14656 59296 14720
rect 59360 14656 59376 14720
rect 59440 14656 59456 14720
rect 59520 14656 59528 14720
rect 59208 13632 59528 14656
rect 59208 13568 59216 13632
rect 59280 13568 59296 13632
rect 59360 13568 59376 13632
rect 59440 13568 59456 13632
rect 59520 13568 59528 13632
rect 59208 12544 59528 13568
rect 59208 12480 59216 12544
rect 59280 12480 59296 12544
rect 59360 12480 59376 12544
rect 59440 12480 59456 12544
rect 59520 12480 59528 12544
rect 59208 11456 59528 12480
rect 59208 11392 59216 11456
rect 59280 11392 59296 11456
rect 59360 11392 59376 11456
rect 59440 11392 59456 11456
rect 59520 11392 59528 11456
rect 59208 10368 59528 11392
rect 59208 10304 59216 10368
rect 59280 10304 59296 10368
rect 59360 10304 59376 10368
rect 59440 10304 59456 10368
rect 59520 10304 59528 10368
rect 59208 9280 59528 10304
rect 59208 9216 59216 9280
rect 59280 9216 59296 9280
rect 59360 9216 59376 9280
rect 59440 9216 59456 9280
rect 59520 9216 59528 9280
rect 59208 8192 59528 9216
rect 59208 8128 59216 8192
rect 59280 8128 59296 8192
rect 59360 8128 59376 8192
rect 59440 8128 59456 8192
rect 59520 8128 59528 8192
rect 59208 7104 59528 8128
rect 59208 7040 59216 7104
rect 59280 7040 59296 7104
rect 59360 7040 59376 7104
rect 59440 7040 59456 7104
rect 59520 7040 59528 7104
rect 59208 6016 59528 7040
rect 59208 5952 59216 6016
rect 59280 5952 59296 6016
rect 59360 5952 59376 6016
rect 59440 5952 59456 6016
rect 59520 5952 59528 6016
rect 55995 5268 56061 5269
rect 55995 5204 55996 5268
rect 56060 5204 56061 5268
rect 55995 5203 56061 5204
rect 54891 4996 54957 4997
rect 54891 4932 54892 4996
rect 54956 4932 54957 4996
rect 54891 4931 54957 4932
rect 54208 4320 54216 4384
rect 54280 4320 54296 4384
rect 54360 4320 54376 4384
rect 54440 4320 54456 4384
rect 54520 4320 54528 4384
rect 54208 3296 54528 4320
rect 54208 3232 54216 3296
rect 54280 3232 54296 3296
rect 54360 3232 54376 3296
rect 54440 3232 54456 3296
rect 54520 3232 54528 3296
rect 53603 2548 53669 2549
rect 53603 2484 53604 2548
rect 53668 2484 53669 2548
rect 53603 2483 53669 2484
rect 49739 2276 49805 2277
rect 49739 2212 49740 2276
rect 49804 2212 49805 2276
rect 49739 2211 49805 2212
rect 54208 2208 54528 3232
rect 54208 2144 54216 2208
rect 54280 2144 54296 2208
rect 54360 2144 54376 2208
rect 54440 2144 54456 2208
rect 54520 2144 54528 2208
rect 54208 2128 54528 2144
rect 54894 2005 54954 4931
rect 55998 3773 56058 5203
rect 59208 4928 59528 5952
rect 59208 4864 59216 4928
rect 59280 4864 59296 4928
rect 59360 4864 59376 4928
rect 59440 4864 59456 4928
rect 59520 4864 59528 4928
rect 59208 3840 59528 4864
rect 59208 3776 59216 3840
rect 59280 3776 59296 3840
rect 59360 3776 59376 3840
rect 59440 3776 59456 3840
rect 59520 3776 59528 3840
rect 55995 3772 56061 3773
rect 55995 3708 55996 3772
rect 56060 3708 56061 3772
rect 55995 3707 56061 3708
rect 59208 2752 59528 3776
rect 59208 2688 59216 2752
rect 59280 2688 59296 2752
rect 59360 2688 59376 2752
rect 59440 2688 59456 2752
rect 59520 2688 59528 2752
rect 59208 2128 59528 2688
rect 64208 67488 64528 67504
rect 64208 67424 64216 67488
rect 64280 67424 64296 67488
rect 64360 67424 64376 67488
rect 64440 67424 64456 67488
rect 64520 67424 64528 67488
rect 64208 66400 64528 67424
rect 64208 66336 64216 66400
rect 64280 66336 64296 66400
rect 64360 66336 64376 66400
rect 64440 66336 64456 66400
rect 64520 66336 64528 66400
rect 64208 65312 64528 66336
rect 64208 65248 64216 65312
rect 64280 65248 64296 65312
rect 64360 65248 64376 65312
rect 64440 65248 64456 65312
rect 64520 65248 64528 65312
rect 64208 64224 64528 65248
rect 64208 64160 64216 64224
rect 64280 64160 64296 64224
rect 64360 64160 64376 64224
rect 64440 64160 64456 64224
rect 64520 64160 64528 64224
rect 64208 63136 64528 64160
rect 64208 63072 64216 63136
rect 64280 63072 64296 63136
rect 64360 63072 64376 63136
rect 64440 63072 64456 63136
rect 64520 63072 64528 63136
rect 64208 62048 64528 63072
rect 64208 61984 64216 62048
rect 64280 61984 64296 62048
rect 64360 61984 64376 62048
rect 64440 61984 64456 62048
rect 64520 61984 64528 62048
rect 64208 60960 64528 61984
rect 64208 60896 64216 60960
rect 64280 60896 64296 60960
rect 64360 60896 64376 60960
rect 64440 60896 64456 60960
rect 64520 60896 64528 60960
rect 64208 59872 64528 60896
rect 64208 59808 64216 59872
rect 64280 59808 64296 59872
rect 64360 59808 64376 59872
rect 64440 59808 64456 59872
rect 64520 59808 64528 59872
rect 64208 58784 64528 59808
rect 64208 58720 64216 58784
rect 64280 58720 64296 58784
rect 64360 58720 64376 58784
rect 64440 58720 64456 58784
rect 64520 58720 64528 58784
rect 64208 57696 64528 58720
rect 64208 57632 64216 57696
rect 64280 57632 64296 57696
rect 64360 57632 64376 57696
rect 64440 57632 64456 57696
rect 64520 57632 64528 57696
rect 64208 56608 64528 57632
rect 64208 56544 64216 56608
rect 64280 56544 64296 56608
rect 64360 56544 64376 56608
rect 64440 56544 64456 56608
rect 64520 56544 64528 56608
rect 64208 55520 64528 56544
rect 64208 55456 64216 55520
rect 64280 55456 64296 55520
rect 64360 55456 64376 55520
rect 64440 55456 64456 55520
rect 64520 55456 64528 55520
rect 64208 54432 64528 55456
rect 64208 54368 64216 54432
rect 64280 54368 64296 54432
rect 64360 54368 64376 54432
rect 64440 54368 64456 54432
rect 64520 54368 64528 54432
rect 64208 53344 64528 54368
rect 64208 53280 64216 53344
rect 64280 53280 64296 53344
rect 64360 53280 64376 53344
rect 64440 53280 64456 53344
rect 64520 53280 64528 53344
rect 64208 52256 64528 53280
rect 64208 52192 64216 52256
rect 64280 52192 64296 52256
rect 64360 52192 64376 52256
rect 64440 52192 64456 52256
rect 64520 52192 64528 52256
rect 64208 51168 64528 52192
rect 64208 51104 64216 51168
rect 64280 51104 64296 51168
rect 64360 51104 64376 51168
rect 64440 51104 64456 51168
rect 64520 51104 64528 51168
rect 64208 50080 64528 51104
rect 64208 50016 64216 50080
rect 64280 50016 64296 50080
rect 64360 50016 64376 50080
rect 64440 50016 64456 50080
rect 64520 50016 64528 50080
rect 64208 48992 64528 50016
rect 64208 48928 64216 48992
rect 64280 48928 64296 48992
rect 64360 48928 64376 48992
rect 64440 48928 64456 48992
rect 64520 48928 64528 48992
rect 64208 47904 64528 48928
rect 64208 47840 64216 47904
rect 64280 47840 64296 47904
rect 64360 47840 64376 47904
rect 64440 47840 64456 47904
rect 64520 47840 64528 47904
rect 64208 46816 64528 47840
rect 64208 46752 64216 46816
rect 64280 46752 64296 46816
rect 64360 46752 64376 46816
rect 64440 46752 64456 46816
rect 64520 46752 64528 46816
rect 64208 45728 64528 46752
rect 64208 45664 64216 45728
rect 64280 45664 64296 45728
rect 64360 45664 64376 45728
rect 64440 45664 64456 45728
rect 64520 45664 64528 45728
rect 64208 44640 64528 45664
rect 64208 44576 64216 44640
rect 64280 44576 64296 44640
rect 64360 44576 64376 44640
rect 64440 44576 64456 44640
rect 64520 44576 64528 44640
rect 64208 43552 64528 44576
rect 64208 43488 64216 43552
rect 64280 43488 64296 43552
rect 64360 43488 64376 43552
rect 64440 43488 64456 43552
rect 64520 43488 64528 43552
rect 64208 42464 64528 43488
rect 64208 42400 64216 42464
rect 64280 42400 64296 42464
rect 64360 42400 64376 42464
rect 64440 42400 64456 42464
rect 64520 42400 64528 42464
rect 64208 41376 64528 42400
rect 64208 41312 64216 41376
rect 64280 41312 64296 41376
rect 64360 41312 64376 41376
rect 64440 41312 64456 41376
rect 64520 41312 64528 41376
rect 64208 40288 64528 41312
rect 64208 40224 64216 40288
rect 64280 40224 64296 40288
rect 64360 40224 64376 40288
rect 64440 40224 64456 40288
rect 64520 40224 64528 40288
rect 64208 39200 64528 40224
rect 64208 39136 64216 39200
rect 64280 39136 64296 39200
rect 64360 39136 64376 39200
rect 64440 39136 64456 39200
rect 64520 39136 64528 39200
rect 64208 38112 64528 39136
rect 64208 38048 64216 38112
rect 64280 38048 64296 38112
rect 64360 38048 64376 38112
rect 64440 38048 64456 38112
rect 64520 38048 64528 38112
rect 64208 37024 64528 38048
rect 64208 36960 64216 37024
rect 64280 36960 64296 37024
rect 64360 36960 64376 37024
rect 64440 36960 64456 37024
rect 64520 36960 64528 37024
rect 64208 35936 64528 36960
rect 64208 35872 64216 35936
rect 64280 35872 64296 35936
rect 64360 35872 64376 35936
rect 64440 35872 64456 35936
rect 64520 35872 64528 35936
rect 64208 34848 64528 35872
rect 64208 34784 64216 34848
rect 64280 34784 64296 34848
rect 64360 34784 64376 34848
rect 64440 34784 64456 34848
rect 64520 34784 64528 34848
rect 64208 33760 64528 34784
rect 64208 33696 64216 33760
rect 64280 33696 64296 33760
rect 64360 33696 64376 33760
rect 64440 33696 64456 33760
rect 64520 33696 64528 33760
rect 64208 32672 64528 33696
rect 64208 32608 64216 32672
rect 64280 32608 64296 32672
rect 64360 32608 64376 32672
rect 64440 32608 64456 32672
rect 64520 32608 64528 32672
rect 64208 31584 64528 32608
rect 64208 31520 64216 31584
rect 64280 31520 64296 31584
rect 64360 31520 64376 31584
rect 64440 31520 64456 31584
rect 64520 31520 64528 31584
rect 64208 30496 64528 31520
rect 64208 30432 64216 30496
rect 64280 30432 64296 30496
rect 64360 30432 64376 30496
rect 64440 30432 64456 30496
rect 64520 30432 64528 30496
rect 64208 29408 64528 30432
rect 64208 29344 64216 29408
rect 64280 29344 64296 29408
rect 64360 29344 64376 29408
rect 64440 29344 64456 29408
rect 64520 29344 64528 29408
rect 64208 28320 64528 29344
rect 64208 28256 64216 28320
rect 64280 28256 64296 28320
rect 64360 28256 64376 28320
rect 64440 28256 64456 28320
rect 64520 28256 64528 28320
rect 64208 27232 64528 28256
rect 64208 27168 64216 27232
rect 64280 27168 64296 27232
rect 64360 27168 64376 27232
rect 64440 27168 64456 27232
rect 64520 27168 64528 27232
rect 64208 26144 64528 27168
rect 64208 26080 64216 26144
rect 64280 26080 64296 26144
rect 64360 26080 64376 26144
rect 64440 26080 64456 26144
rect 64520 26080 64528 26144
rect 64208 25056 64528 26080
rect 64208 24992 64216 25056
rect 64280 24992 64296 25056
rect 64360 24992 64376 25056
rect 64440 24992 64456 25056
rect 64520 24992 64528 25056
rect 64208 23968 64528 24992
rect 64208 23904 64216 23968
rect 64280 23904 64296 23968
rect 64360 23904 64376 23968
rect 64440 23904 64456 23968
rect 64520 23904 64528 23968
rect 64208 22880 64528 23904
rect 64208 22816 64216 22880
rect 64280 22816 64296 22880
rect 64360 22816 64376 22880
rect 64440 22816 64456 22880
rect 64520 22816 64528 22880
rect 64208 21792 64528 22816
rect 64208 21728 64216 21792
rect 64280 21728 64296 21792
rect 64360 21728 64376 21792
rect 64440 21728 64456 21792
rect 64520 21728 64528 21792
rect 64208 20704 64528 21728
rect 64208 20640 64216 20704
rect 64280 20640 64296 20704
rect 64360 20640 64376 20704
rect 64440 20640 64456 20704
rect 64520 20640 64528 20704
rect 64208 19616 64528 20640
rect 64208 19552 64216 19616
rect 64280 19552 64296 19616
rect 64360 19552 64376 19616
rect 64440 19552 64456 19616
rect 64520 19552 64528 19616
rect 64208 18528 64528 19552
rect 64208 18464 64216 18528
rect 64280 18464 64296 18528
rect 64360 18464 64376 18528
rect 64440 18464 64456 18528
rect 64520 18464 64528 18528
rect 64208 17440 64528 18464
rect 64208 17376 64216 17440
rect 64280 17376 64296 17440
rect 64360 17376 64376 17440
rect 64440 17376 64456 17440
rect 64520 17376 64528 17440
rect 64208 16352 64528 17376
rect 64208 16288 64216 16352
rect 64280 16288 64296 16352
rect 64360 16288 64376 16352
rect 64440 16288 64456 16352
rect 64520 16288 64528 16352
rect 64208 15264 64528 16288
rect 64208 15200 64216 15264
rect 64280 15200 64296 15264
rect 64360 15200 64376 15264
rect 64440 15200 64456 15264
rect 64520 15200 64528 15264
rect 64208 14176 64528 15200
rect 64208 14112 64216 14176
rect 64280 14112 64296 14176
rect 64360 14112 64376 14176
rect 64440 14112 64456 14176
rect 64520 14112 64528 14176
rect 64208 13088 64528 14112
rect 64208 13024 64216 13088
rect 64280 13024 64296 13088
rect 64360 13024 64376 13088
rect 64440 13024 64456 13088
rect 64520 13024 64528 13088
rect 64208 12000 64528 13024
rect 64208 11936 64216 12000
rect 64280 11936 64296 12000
rect 64360 11936 64376 12000
rect 64440 11936 64456 12000
rect 64520 11936 64528 12000
rect 64208 10912 64528 11936
rect 64208 10848 64216 10912
rect 64280 10848 64296 10912
rect 64360 10848 64376 10912
rect 64440 10848 64456 10912
rect 64520 10848 64528 10912
rect 64208 9824 64528 10848
rect 64208 9760 64216 9824
rect 64280 9760 64296 9824
rect 64360 9760 64376 9824
rect 64440 9760 64456 9824
rect 64520 9760 64528 9824
rect 64208 8736 64528 9760
rect 64208 8672 64216 8736
rect 64280 8672 64296 8736
rect 64360 8672 64376 8736
rect 64440 8672 64456 8736
rect 64520 8672 64528 8736
rect 64208 7648 64528 8672
rect 64208 7584 64216 7648
rect 64280 7584 64296 7648
rect 64360 7584 64376 7648
rect 64440 7584 64456 7648
rect 64520 7584 64528 7648
rect 64208 6560 64528 7584
rect 64208 6496 64216 6560
rect 64280 6496 64296 6560
rect 64360 6496 64376 6560
rect 64440 6496 64456 6560
rect 64520 6496 64528 6560
rect 64208 5472 64528 6496
rect 64208 5408 64216 5472
rect 64280 5408 64296 5472
rect 64360 5408 64376 5472
rect 64440 5408 64456 5472
rect 64520 5408 64528 5472
rect 64208 4384 64528 5408
rect 64643 4588 64709 4589
rect 64643 4524 64644 4588
rect 64708 4524 64709 4588
rect 64643 4523 64709 4524
rect 64208 4320 64216 4384
rect 64280 4320 64296 4384
rect 64360 4320 64376 4384
rect 64440 4320 64456 4384
rect 64520 4320 64528 4384
rect 64208 3296 64528 4320
rect 64208 3232 64216 3296
rect 64280 3232 64296 3296
rect 64360 3232 64376 3296
rect 64440 3232 64456 3296
rect 64520 3232 64528 3296
rect 64208 2208 64528 3232
rect 64208 2144 64216 2208
rect 64280 2144 64296 2208
rect 64360 2144 64376 2208
rect 64440 2144 64456 2208
rect 64520 2144 64528 2208
rect 64208 2128 64528 2144
rect 64646 2005 64706 4523
rect 46611 2004 46677 2005
rect 46611 1940 46612 2004
rect 46676 1940 46677 2004
rect 46611 1939 46677 1940
rect 54891 2004 54957 2005
rect 54891 1940 54892 2004
rect 54956 1940 54957 2004
rect 54891 1939 54957 1940
rect 64643 2004 64709 2005
rect 64643 1940 64644 2004
rect 64708 1940 64709 2004
rect 64643 1939 64709 1940
rect 41275 1324 41341 1325
rect 41275 1260 41276 1324
rect 41340 1260 41341 1324
rect 41275 1259 41341 1260
rect 31891 1188 31957 1189
rect 31891 1124 31892 1188
rect 31956 1124 31957 1188
rect 31891 1123 31957 1124
use sky130_fd_sc_hd__decap_4  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2576 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  input296 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_238 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1624635492
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1624635492
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output575 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1522 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1624635492
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1624635492
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output577
timestamp 1624635492
transform -1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output576
timestamp 1624635492
transform -1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1523
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1624635492
transform 1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1624635492
transform 1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output580
timestamp 1624635492
transform -1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output579
timestamp 1624635492
transform -1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output578
timestamp 1624635492
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1624635492
transform 1 0 9936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1624635492
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output581
timestamp 1624635492
transform -1 0 9936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1524
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1624635492
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1624635492
transform 1 0 10672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output582
timestamp 1624635492
transform -1 0 10672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output527
timestamp 1624635492
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1525
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133
timestamp 1624635492
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1624635492
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output482
timestamp 1624635492
transform 1 0 12236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output479
timestamp 1624635492
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output436
timestamp 1624635492
transform -1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_6
timestamp 1624635492
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input308
timestamp 1624635492
transform -1 0 2300 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1624635492
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1624635492
transform 1 0 2300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input319
timestamp 1624635492
transform -1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output398
timestamp 1624635492
transform -1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output587
timestamp 1624635492
transform -1 0 3680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1624635492
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1624635492
transform 1 0 3680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2944 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_28
timestamp 1624635492
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output598
timestamp 1624635492
transform -1 0 4416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output603
timestamp 1624635492
transform -1 0 4600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1624635492
transform 1 0 4416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_38
timestamp 1624635492
transform 1 0 4600 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output601
timestamp 1624635492
transform -1 0 5152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1624635492
transform 1 0 5152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output602
timestamp 1624635492
transform -1 0 5888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output604
timestamp 1624635492
transform -1 0 5796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1624635492
transform 1 0 5336 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1624635492
transform 1 0 5888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1624635492
transform 1 0 5796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output606
timestamp 1624635492
transform -1 0 6532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56
timestamp 1624635492
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1624635492
transform 1 0 6532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input298
timestamp 1624635492
transform 1 0 6900 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output607
timestamp 1624635492
transform -1 0 7176 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7176 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1624635492
transform 1 0 7176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input217
timestamp 1624635492
transform -1 0 8096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input299
timestamp 1624635492
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_72
timestamp 1624635492
transform 1 0 7728 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1624635492
transform 1 0 7820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input301
timestamp 1624635492
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1624635492
transform 1 0 8096 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output583
timestamp 1624635492
transform -1 0 8832 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp 1624635492
transform 1 0 8832 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_80
timestamp 1624635492
transform 1 0 8464 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output584
timestamp 1624635492
transform -1 0 9568 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_92
timestamp 1624635492
transform 1 0 9568 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1624635492
transform 1 0 9384 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output585
timestamp 1624635492
transform -1 0 10304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output586
timestamp 1624635492
transform -1 0 10120 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1624635492
transform 1 0 10120 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1624635492
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_108
timestamp 1624635492
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1624635492
transform 1 0 10304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output589
timestamp 1624635492
transform -1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output588
timestamp 1624635492
transform -1 0 11040 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 12052 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1624635492
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_127
timestamp 1624635492
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_131
timestamp 1624635492
transform 1 0 13156 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1624635492
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output593
timestamp 1624635492
transform -1 0 13524 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output591
timestamp 1624635492
transform -1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output590
timestamp 1624635492
transform -1 0 13156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1624635492
transform 1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_14
timestamp 1624635492
transform 1 0 2392 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_6
timestamp 1624635492
transform 1 0 1656 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input322
timestamp 1624635492
transform -1 0 2760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input297
timestamp 1624635492
transform -1 0 1656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1624635492
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 1624635492
transform 1 0 4048 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1624635492
transform 1 0 3404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input215_A
timestamp 1624635492
transform -1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input324
timestamp 1624635492
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input323
timestamp 1624635492
transform -1 0 3404 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1624635492
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1624635492
transform 1 0 5336 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output605
timestamp 1624635492
transform -1 0 5336 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_78
timestamp 1624635492
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_72
timestamp 1624635492
transform 1 0 7728 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_65
timestamp 1624635492
transform 1 0 7084 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input303
timestamp 1624635492
transform 1 0 8372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input302
timestamp 1624635492
transform 1 0 7452 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input300
timestamp 1624635492
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1624635492
transform 1 0 9936 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1624635492
transform 1 0 9292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_82
timestamp 1624635492
transform 1 0 8648 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input304
timestamp 1624635492
transform 1 0 9016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input215
timestamp 1624635492
transform -1 0 9936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1624635492
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1624635492
transform 1 0 10580 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output592
timestamp 1624635492
transform -1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input209
timestamp 1624635492
transform -1 0 10580 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input201
timestamp 1624635492
transform -1 0 11224 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1624635492
transform 1 0 13156 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1624635492
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output595
timestamp 1624635492
transform -1 0 13892 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output594
timestamp 1624635492
transform -1 0 13156 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1624635492
transform 1 0 2760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1624635492
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output397
timestamp 1624635492
transform -1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input330
timestamp 1624635492
transform -1 0 2760 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1624635492
transform 1 0 4692 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1624635492
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_25
timestamp 1624635492
transform 1 0 3404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input352
timestamp 1624635492
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input325
timestamp 1624635492
transform -1 0 4692 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1624635492
transform 1 0 5980 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_46
timestamp 1624635492
transform 1 0 5336 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input328
timestamp 1624635492
transform 1 0 6348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input327
timestamp 1624635492
transform 1 0 5704 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input326
timestamp 1624635492
transform -1 0 5336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_78
timestamp 1624635492
transform 1 0 8280 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1624635492
transform 1 0 7912 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_67
timestamp 1624635492
transform 1 0 7268 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1624635492
transform 1 0 6624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input332
timestamp 1624635492
transform 1 0 7636 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input331
timestamp 1624635492
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input312
timestamp 1624635492
transform -1 0 8648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_94
timestamp 1624635492
transform 1 0 9752 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1624635492
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input305
timestamp 1624635492
transform -1 0 9752 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1624635492
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_111
timestamp 1624635492
transform 1 0 11316 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1624635492
transform 1 0 10672 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1624635492
transform 1 0 10304 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input228
timestamp 1624635492
transform -1 0 10672 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input206
timestamp 1624635492
transform -1 0 11316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input189
timestamp 1624635492
transform -1 0 11960 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_132
timestamp 1624635492
transform 1 0 13248 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_125
timestamp 1624635492
transform 1 0 12604 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1624635492
transform -1 0 12604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1624635492
transform -1 0 13248 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1624635492
transform -1 0 13892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1624635492
transform 1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1624635492
transform 1 0 1656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input355
timestamp 1624635492
transform -1 0 2944 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input341
timestamp 1624635492
transform 1 0 2024 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input329
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1624635492
transform 1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1624635492
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_20
timestamp 1624635492
transform 1 0 2944 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input358
timestamp 1624635492
transform -1 0 4876 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input357
timestamp 1624635492
transform -1 0 4232 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input356
timestamp 1624635492
transform -1 0 3588 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1624635492
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1624635492
transform 1 0 5520 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_41
timestamp 1624635492
transform 1 0 4876 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input359
timestamp 1624635492
transform -1 0 5520 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1624635492
transform 1 0 7820 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_69
timestamp 1624635492
transform 1 0 7452 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_65
timestamp 1624635492
transform 1 0 7084 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input335
timestamp 1624635492
transform 1 0 8188 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input334
timestamp 1624635492
transform 1 0 7544 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input333
timestamp 1624635492
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1624635492
transform 1 0 9752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_87
timestamp 1624635492
transform 1 0 9108 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_80
timestamp 1624635492
transform 1 0 8464 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input336
timestamp 1624635492
transform -1 0 9108 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input307
timestamp 1624635492
transform 1 0 10120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input306
timestamp 1624635492
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1624635492
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_101
timestamp 1624635492
transform 1 0 10396 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1624635492
transform -1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input250
timestamp 1624635492
transform -1 0 11224 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_134
timestamp 1624635492
transform 1 0 13432 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_127
timestamp 1624635492
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_120
timestamp 1624635492
transform 1 0 12144 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input199
timestamp 1624635492
transform -1 0 12788 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input155
timestamp 1624635492
transform -1 0 13432 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_18
timestamp 1624635492
transform 1 0 2760 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1624635492
transform 1 0 2116 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output435
timestamp 1624635492
transform -1 0 2116 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input363
timestamp 1624635492
transform -1 0 2760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1624635492
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_25
timestamp 1624635492
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input296_A
timestamp 1624635492
transform -1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input364
timestamp 1624635492
transform -1 0 3404 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_57
timestamp 1624635492
transform 1 0 6348 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1624635492
transform 1 0 5796 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp 1624635492
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_40
timestamp 1624635492
transform 1 0 4784 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input300_A
timestamp 1624635492
transform -1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input361
timestamp 1624635492
transform -1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input360
timestamp 1624635492
transform -1 0 5152 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1624635492
transform 1 0 8004 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_69
timestamp 1624635492
transform 1 0 7452 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1624635492
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input250_A
timestamp 1624635492
transform -1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input208_A
timestamp 1624635492
transform -1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input199_A
timestamp 1624635492
transform -1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input337
timestamp 1624635492
transform 1 0 8372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_94
timestamp 1624635492
transform 1 0 9752 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_82
timestamp 1624635492
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input309
timestamp 1624635492
transform 1 0 10120 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _136_
timestamp 1624635492
transform -1 0 9752 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_118
timestamp 1624635492
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_114
timestamp 1624635492
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_108
timestamp 1624635492
transform 1 0 11040 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 1624635492
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input310
timestamp 1624635492
transform 1 0 10764 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input294
timestamp 1624635492
transform -1 0 11960 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_132
timestamp 1624635492
transform 1 0 13248 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_125
timestamp 1624635492
transform 1 0 12604 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input208
timestamp 1624635492
transform -1 0 12604 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input202
timestamp 1624635492
transform -1 0 13248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1624635492
transform -1 0 13892 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1624635492
transform -1 0 1656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input362
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1624635492
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1624635492
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input366
timestamp 1624635492
transform 1 0 2024 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_13
timestamp 1624635492
transform 1 0 2300 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1624635492
transform 1 0 2208 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input308_A
timestamp 1624635492
transform -1 0 2760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_19
timestamp 1624635492
transform 1 0 2852 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1624635492
transform 1 0 2760 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input365
timestamp 1624635492
transform -1 0 3220 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input322_A
timestamp 1624635492
transform -1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1624635492
transform 1 0 3220 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1624635492
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input319_A
timestamp 1624635492
transform -1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_29
timestamp 1624635492
transform 1 0 3772 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1624635492
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input323_A
timestamp 1624635492
transform -1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input324_A
timestamp 1624635492
transform -1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1624635492
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input325_A
timestamp 1624635492
transform -1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input330_A
timestamp 1624635492
transform -1 0 4600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1624635492
transform 1 0 4324 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1624635492
transform 1 0 4600 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input338_A
timestamp 1624635492
transform -1 0 5244 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1624635492
transform 1 0 4876 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_42
timestamp 1624635492
transform 1 0 4968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input326_A
timestamp 1624635492
transform -1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input333_A
timestamp 1624635492
transform -1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1624635492
transform 1 0 5428 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_45
timestamp 1624635492
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input327_A
timestamp 1624635492
transform -1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_53
timestamp 1624635492
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1624635492
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input328_A
timestamp 1624635492
transform -1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1624635492
transform 1 0 6348 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input283_A
timestamp 1624635492
transform -1 0 7452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input298_A
timestamp 1624635492
transform -1 0 6900 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input299_A
timestamp 1624635492
transform -1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input302_A
timestamp 1624635492
transform -1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_63
timestamp 1624635492
transform 1 0 6900 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_61
timestamp 1624635492
transform 1 0 6716 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_64
timestamp 1624635492
transform 1 0 6992 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input209_A
timestamp 1624635492
transform -1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input217_A
timestamp 1624635492
transform -1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1624635492
transform 1 0 7452 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1624635492
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_70
timestamp 1624635492
transform 1 0 7544 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input338
timestamp 1624635492
transform -1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1624635492
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input339
timestamp 1624635492
transform -1 0 9476 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_82
timestamp 1624635492
transform 1 0 8648 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input340
timestamp 1624635492
transform 1 0 9844 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input342
timestamp 1624635492
transform -1 0 10304 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input167_A
timestamp 1624635492
transform -1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_91
timestamp 1624635492
transform 1 0 9476 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1624635492
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_98
timestamp 1624635492
transform 1 0 10120 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_106
timestamp 1624635492
transform 1 0 10856 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_100
timestamp 1624635492
transform 1 0 10304 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_106
timestamp 1624635492
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input311
timestamp 1624635492
transform -1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input318
timestamp 1624635492
transform -1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_110
timestamp 1624635492
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_110
timestamp 1624635492
transform 1 0 11224 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input313
timestamp 1624635492
transform -1 0 11868 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1624635492
transform -1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1624635492
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_117
timestamp 1624635492
transform 1 0 11868 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input283
timestamp 1624635492
transform -1 0 12604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input314
timestamp 1624635492
transform -1 0 12512 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input315
timestamp 1624635492
transform 1 0 12880 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1624635492
transform 1 0 12604 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_124
timestamp 1624635492
transform 1 0 12512 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input214
timestamp 1624635492
transform -1 0 13248 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1624635492
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1624635492
transform 1 0 13156 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input207
timestamp 1624635492
transform -1 0 13892 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input272
timestamp 1624635492
transform -1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1624635492
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1624635492
transform 1 0 2208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1624635492
transform 1 0 1656 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input297_A
timestamp 1624635492
transform -1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input367
timestamp 1624635492
transform -1 0 1656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2576 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1624635492
transform 1 0 4324 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input355_A
timestamp 1624635492
transform -1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1624635492
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_47
timestamp 1624635492
transform 1 0 5428 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1624635492
transform 1 0 4876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input359_A
timestamp 1624635492
transform -1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input358_A
timestamp 1624635492
transform -1 0 5428 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_77
timestamp 1624635492
transform 1 0 8188 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 1624635492
transform 1 0 7452 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input301_A
timestamp 1624635492
transform -1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_2  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6808 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_94
timestamp 1624635492
transform 1 0 9752 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1624635492
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1624635492
transform 1 0 8924 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input261_A
timestamp 1624635492
transform -1 0 9200 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input206_A
timestamp 1624635492
transform -1 0 9752 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input189_A
timestamp 1624635492
transform -1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1624635492
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_107
timestamp 1624635492
transform 1 0 10948 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_100
timestamp 1624635492
transform 1 0 10304 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input345
timestamp 1624635492
transform -1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input343
timestamp 1624635492
transform -1 0 10948 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1624635492
transform 1 0 13156 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_122
timestamp 1624635492
transform 1 0 12328 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input317
timestamp 1624635492
transform 1 0 13524 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input316
timestamp 1624635492
transform -1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_19
timestamp 1624635492
transform 1 0 2852 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_15
timestamp 1624635492
transform 1 0 2484 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_11
timestamp 1624635492
transform 1 0 2116 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_5
timestamp 1624635492
transform 1 0 1564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input341_A
timestamp 1624635492
transform -1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input329_A
timestamp 1624635492
transform -1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _330_
timestamp 1624635492
transform 1 0 2576 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_38
timestamp 1624635492
transform 1 0 4600 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1624635492
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_25
timestamp 1624635492
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input357_A
timestamp 1624635492
transform -1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input356_A
timestamp 1624635492
transform -1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input352_A
timestamp 1624635492
transform -1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_58
timestamp 1624635492
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp 1624635492
transform 1 0 5888 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1624635492
transform 1 0 5336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A1
timestamp 1624635492
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input361_A
timestamp 1624635492
transform -1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input360_A
timestamp 1624635492
transform -1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_79
timestamp 1624635492
transform 1 0 8372 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_71
timestamp 1624635492
transform 1 0 7636 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_68
timestamp 1624635492
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1624635492
transform 1 0 6992 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input332_A
timestamp 1624635492
transform -1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input331_A
timestamp 1624635492
transform -1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input303_A
timestamp 1624635492
transform -1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_99
timestamp 1624635492
transform 1 0 10212 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_95
timestamp 1624635492
transform 1 0 9844 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_89
timestamp 1624635492
transform 1 0 9292 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1624635492
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input305_A
timestamp 1624635492
transform -1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input304_A
timestamp 1624635492
transform -1 0 9292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1624635492
transform 1 0 11960 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_109
timestamp 1624635492
transform 1 0 11132 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1624635492
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input201_A
timestamp 1624635492
transform -1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input346
timestamp 1624635492
transform -1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input344
timestamp 1624635492
transform -1 0 11132 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_132
timestamp 1624635492
transform 1 0 13248 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1624635492
transform 1 0 12604 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input348
timestamp 1624635492
transform 1 0 12972 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input347
timestamp 1624635492
transform -1 0 12604 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input320
timestamp 1624635492
transform -1 0 13892 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1624635492
transform 1 0 2760 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1624635492
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output396
timestamp 1624635492
transform -1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _202_
timestamp 1624635492
transform 1 0 2484 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1624635492
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_34
timestamp 1624635492
transform 1 0 4232 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1624635492
transform 1 0 3864 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1624635492
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__D
timestamp 1624635492
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input364_A
timestamp 1624635492
transform -1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input363_A
timestamp 1624635492
transform -1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_49
timestamp 1624635492
transform 1 0 5612 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1624635492
transform 1 0 5060 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output575_A
timestamp 1624635492
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output398_A
timestamp 1624635492
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1624635492
transform 1 0 8188 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1624635492
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_70
timestamp 1624635492
transform 1 0 7544 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 1624635492
transform 1 0 6992 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B1
timestamp 1624635492
transform -1 0 6992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input335_A
timestamp 1624635492
transform -1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input334_A
timestamp 1624635492
transform -1 0 7544 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_98
timestamp 1624635492
transform 1 0 10120 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_95
timestamp 1624635492
transform 1 0 9844 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1624635492
transform 1 0 9476 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_88
timestamp 1624635492
transform 1 0 9200 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1624635492
transform 1 0 8832 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_81
timestamp 1624635492
transform 1 0 8556 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input312_A
timestamp 1624635492
transform -1 0 8832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input307_A
timestamp 1624635492
transform -1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input306_A
timestamp 1624635492
transform -1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_119
timestamp 1624635492
transform 1 0 12052 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1624635492
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input228_A
timestamp 1624635492
transform -1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input166_A
timestamp 1624635492
transform -1 0 12052 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_132
timestamp 1624635492
transform 1 0 13248 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1624635492
transform 1 0 12604 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1624635492
transform -1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input349
timestamp 1624635492
transform -1 0 13248 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_17
timestamp 1624635492
transform 1 0 2668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1624635492
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_5
timestamp 1624635492
transform 1 0 1564 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input367_A
timestamp 1624635492
transform -1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input366_A
timestamp 1624635492
transform -1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input362_A
timestamp 1624635492
transform -1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_38
timestamp 1624635492
transform 1 0 4600 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1624635492
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_25
timestamp 1624635492
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output436_A
timestamp 1624635492
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output397_A
timestamp 1624635492
transform -1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input365_A
timestamp 1624635492
transform -1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_56
timestamp 1624635492
transform 1 0 6256 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_48
timestamp 1624635492
transform 1 0 5520 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output577_A
timestamp 1624635492
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output576_A
timestamp 1624635492
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_79
timestamp 1624635492
transform 1 0 8372 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_71
timestamp 1624635492
transform 1 0 7636 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1624635492
transform 1 0 7084 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_62
timestamp 1624635492
transform 1 0 6808 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output578_A
timestamp 1624635492
transform -1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A2
timestamp 1624635492
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input337_A
timestamp 1624635492
transform -1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1624635492
transform 1 0 10120 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_95
timestamp 1624635492
transform 1 0 9844 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_89
timestamp 1624635492
transform 1 0 9292 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1624635492
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input336_A
timestamp 1624635492
transform -1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input309_A
timestamp 1624635492
transform -1 0 10120 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1624635492
transform 1 0 11960 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_115
timestamp 1624635492
transform 1 0 11684 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_111
timestamp 1624635492
transform 1 0 11316 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_105
timestamp 1624635492
transform 1 0 10764 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1624635492
transform 1 0 10488 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input311_A
timestamp 1624635492
transform -1 0 11316 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input310_A
timestamp 1624635492
transform -1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input239_A
timestamp 1624635492
transform -1 0 11960 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_130
timestamp 1624635492
transform 1 0 13064 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_124
timestamp 1624635492
transform 1 0 12512 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input207_A
timestamp 1624635492
transform -1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input155_A
timestamp 1624635492
transform -1 0 13064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input350
timestamp 1624635492
transform -1 0 13708 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1624635492
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output434
timestamp 1624635492
transform -1 0 2116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _339_
timestamp 1624635492
transform -1 0 4048 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1624635492
transform 1 0 4600 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_32
timestamp 1624635492
transform 1 0 4048 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__D
timestamp 1624635492
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1624635492
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1624635492
transform 1 0 5704 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_44
timestamp 1624635492
transform 1 0 5152 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output604_A
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output601_A
timestamp 1624635492
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output598_A
timestamp 1624635492
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1624635492
transform 1 0 8004 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1624635492
transform 1 0 7452 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1624635492
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_60
timestamp 1624635492
transform 1 0 6624 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output596_A
timestamp 1624635492
transform -1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output579_A
timestamp 1624635492
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output538_A
timestamp 1624635492
transform -1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1624635492
transform 1 0 9660 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_87
timestamp 1624635492
transform 1 0 9108 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_81
timestamp 1624635492
transform 1 0 8556 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__B
timestamp 1624635492
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input339_A
timestamp 1624635492
transform -1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1624635492
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1624635492
transform 1 0 10672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input318_A
timestamp 1624635492
transform -1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input294_A
timestamp 1624635492
transform -1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _277_
timestamp 1624635492
transform 1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_134
timestamp 1624635492
transform 1 0 13432 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_128
timestamp 1624635492
transform 1 0 12880 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_120
timestamp 1624635492
transform 1 0 12144 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input214_A
timestamp 1624635492
transform -1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input202_A
timestamp 1624635492
transform -1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1624635492
transform 1 0 2852 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1624635492
transform 1 0 2300 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output435_A
timestamp 1624635492
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output434_A
timestamp 1624635492
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1624635492
transform 1 0 4416 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_33
timestamp 1624635492
transform 1 0 4140 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_27
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1624635492
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__CLK
timestamp 1624635492
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output603_A
timestamp 1624635492
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output587_A
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output605_A
timestamp 1624635492
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__CLK
timestamp 1624635492
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_40
timestamp 1624635492
transform 1 0 4784 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_48
timestamp 1624635492
transform 1 0 5520 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output606_A
timestamp 1624635492
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_56
timestamp 1624635492
transform 1 0 6256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_54
timestamp 1624635492
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1624635492
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1624635492
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_76
timestamp 1624635492
transform 1 0 8096 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_68
timestamp 1624635492
transform 1 0 7360 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_65
timestamp 1624635492
transform 1 0 7084 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1624635492
transform 1 0 6716 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output607_A
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output592_A
timestamp 1624635492
transform -1 0 8096 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output580_A
timestamp 1624635492
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output583_A
timestamp 1624635492
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1624635492
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1624635492
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output560_A
timestamp 1624635492
transform -1 0 9292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_89
timestamp 1624635492
transform 1 0 9292 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1624635492
transform 1 0 9016 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input340_A
timestamp 1624635492
transform -1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output584_A
timestamp 1624635492
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_92
timestamp 1624635492
transform 1 0 9568 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output549_A
timestamp 1624635492
transform -1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_95
timestamp 1624635492
transform 1 0 9844 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1624635492
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_99
timestamp 1624635492
transform 1 0 10212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input342_A
timestamp 1624635492
transform -1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input343_A
timestamp 1624635492
transform -1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__D
timestamp 1624635492
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output484_A
timestamp 1624635492
transform -1 0 10672 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1624635492
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_108
timestamp 1624635492
transform 1 0 11040 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_104
timestamp 1624635492
transform 1 0 10672 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input344_A
timestamp 1624635492
transform -1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1624635492
transform 1 0 11776 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1624635492
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input313_A
timestamp 1624635492
transform -1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1624635492
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1624635492
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_133
timestamp 1624635492
transform 1 0 13340 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_123
timestamp 1624635492
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_131
timestamp 1624635492
transform 1 0 13156 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1624635492
transform 1 0 12604 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input345_A
timestamp 1624635492
transform -1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input316_A
timestamp 1624635492
transform -1 0 13340 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input315_A
timestamp 1624635492
transform -1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input314_A
timestamp 1624635492
transform -1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_12
timestamp 1624635492
transform 1 0 2208 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 1624635492
transform 1 0 1656 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1624635492
transform -1 0 1656 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1624635492
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1624635492
transform 1 0 3312 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1624635492
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624635492
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1624635492
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1624635492
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_98
timestamp 1624635492
transform 1 0 10120 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1624635492
transform 1 0 9568 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output585_A
timestamp 1624635492
transform -1 0 9568 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output581_A
timestamp 1624635492
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114
timestamp 1624635492
transform 1 0 11592 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_108
timestamp 1624635492
transform 1 0 11040 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output527_A
timestamp 1624635492
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1624635492
transform -1 0 11592 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input346_A
timestamp 1624635492
transform -1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1624635492
transform 1 0 13524 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_132
timestamp 1624635492
transform 1 0 13248 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_126
timestamp 1624635492
transform 1 0 12696 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1624635492
transform 1 0 12144 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input347_A
timestamp 1624635492
transform -1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input317_A
timestamp 1624635492
transform -1 0 13524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1624635492
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1624635492
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1624635492
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1624635492
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1624635492
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1624635492
transform 1 0 9752 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1624635492
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output586_A
timestamp 1624635492
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1624635492
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_100
timestamp 1624635492
transform 1 0 10304 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output582_A
timestamp 1624635492
transform -1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output482_A
timestamp 1624635492
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1624635492
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_129
timestamp 1624635492
transform 1 0 12972 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_121
timestamp 1624635492
transform 1 0 12236 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input349_A
timestamp 1624635492
transform -1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input348_A
timestamp 1624635492
transform -1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624635492
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1624635492
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1624635492
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1624635492
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1624635492
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_99
timestamp 1624635492
transform 1 0 10212 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_118
timestamp 1624635492
transform 1 0 11960 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_110
timestamp 1624635492
transform 1 0 11224 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1624635492
transform 1 0 10948 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output589_A
timestamp 1624635492
transform -1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output588_A
timestamp 1624635492
transform -1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_133
timestamp 1624635492
transform 1 0 13340 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1624635492
transform 1 0 12788 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1624635492
transform 1 0 12236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output505_A
timestamp 1624635492
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output477_A
timestamp 1624635492
transform -1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_13
timestamp 1624635492
transform 1 0 2300 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output395_A
timestamp 1624635492
transform -1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1624635492
transform 1 0 4508 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1624635492
transform 1 0 3404 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_49
timestamp 1624635492
transform 1 0 5612 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1624635492
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1624635492
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1624635492
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1624635492
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_135
timestamp 1624635492
transform 1 0 13524 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 1624635492
transform 1 0 12972 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1624635492
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output591_A
timestamp 1624635492
transform 1 0 12236 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output590_A
timestamp 1624635492
transform -1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output479_A
timestamp 1624635492
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1624635492
transform 1 0 2760 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_11
timestamp 1624635492
transform 1 0 2116 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output395
timestamp 1624635492
transform -1 0 2116 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _176_
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_26
timestamp 1624635492
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1624635492
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1624635492
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1624635492
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1624635492
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1624635492
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 1624635492
transform 1 0 12052 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_111
timestamp 1624635492
transform 1 0 11316 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1624635492
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__CLK
timestamp 1624635492
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output593_A
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1624635492
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1624635492
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1624635492
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1624635492
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1624635492
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1624635492
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1624635492
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1624635492
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1624635492
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1624635492
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1624635492
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1624635492
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1624635492
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1624635492
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1624635492
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1624635492
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1624635492
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_17
timestamp 1624635492
transform 1 0 2668 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1624635492
transform 1 0 2116 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output433_A
timestamp 1624635492
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output433
timestamp 1624635492
transform -1 0 2116 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_29
timestamp 1624635492
transform 1 0 3772 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1624635492
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_41
timestamp 1624635492
transform 1 0 4876 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1624635492
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_95
timestamp 1624635492
transform 1 0 9844 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1624635492
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_82
timestamp 1624635492
transform 1 0 8648 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _116_
timestamp 1624635492
transform 1 0 9568 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1624635492
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_107
timestamp 1624635492
transform 1 0 10948 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1624635492
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1624635492
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1624635492
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_55
timestamp 1624635492
transform 1 0 6164 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_50
timestamp 1624635492
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_42
timestamp 1624635492
transform 1 0 4968 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _131_
timestamp 1624635492
transform -1 0 6164 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_79
timestamp 1624635492
transform 1 0 8372 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_67
timestamp 1624635492
transform 1 0 7268 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_99
timestamp 1624635492
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1624635492
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_114
timestamp 1624635492
transform 1 0 11592 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_103
timestamp 1624635492
transform 1 0 10580 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1624635492
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_4  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 11592 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_24_126
timestamp 1624635492
transform 1 0 12696 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_12
timestamp 1624635492
transform 1 0 2208 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1624635492
transform 1 0 1656 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 2208 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1624635492
transform -1 0 1656 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_36
timestamp 1624635492
transform 1 0 4416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_24
timestamp 1624635492
transform 1 0 3312 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1624635492
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1624635492
transform 1 0 5520 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_77
timestamp 1624635492
transform 1 0 8188 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_65
timestamp 1624635492
transform 1 0 7084 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _147_
timestamp 1624635492
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_89
timestamp 1624635492
transform 1 0 9292 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1624635492
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_101
timestamp 1624635492
transform 1 0 10396 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1624635492
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1624635492
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1624635492
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1624635492
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1624635492
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1624635492
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1624635492
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1624635492
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1624635492
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1624635492
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1624635492
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1526
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output477
timestamp 1624635492
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1624635492
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output444
timestamp 1624635492
transform -1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1624635492
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1624635492
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output466
timestamp 1624635492
transform 1 0 16376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624635492
transform -1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_162
timestamp 1624635492
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1527
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1624635492
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output455
timestamp 1624635492
transform 1 0 17940 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1624635492
transform 1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1624635492
transform -1 0 18952 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output560
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1624635492
transform -1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1624635492
transform 1 0 14260 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output483
timestamp 1624635492
transform -1 0 15732 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output505
timestamp 1624635492
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output549
timestamp 1624635492
transform 1 0 14996 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1624635492
transform 1 0 14996 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_147
timestamp 1624635492
transform 1 0 14628 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_155
timestamp 1624635492
transform 1 0 15364 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output481
timestamp 1624635492
transform 1 0 16100 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output489
timestamp 1624635492
transform 1 0 15732 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1624635492
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1624635492
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output480
timestamp 1624635492
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output484
timestamp 1624635492
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1624635492
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_171
timestamp 1624635492
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _221_
timestamp 1624635492
transform 1 0 17296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output475
timestamp 1624635492
transform 1 0 17940 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output476
timestamp 1624635492
transform 1 0 17940 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1624635492
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1624635492
transform 1 0 17572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 18952 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 18952 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1624635492
transform 1 0 18308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1624635492
transform 1 0 18308 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output596
timestamp 1624635492
transform -1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1624635492
transform 1 0 13892 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output571
timestamp 1624635492
transform 1 0 15272 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_147
timestamp 1624635492
transform 1 0 14628 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_153
timestamp 1624635492
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output494
timestamp 1624635492
transform -1 0 16376 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_158
timestamp 1624635492
transform 1 0 15640 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_166
timestamp 1624635492
transform 1 0 16376 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_170
timestamp 1624635492
transform 1 0 16744 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1624635492
transform -1 0 17572 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output478
timestamp 1624635492
transform 1 0 17940 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1624635492
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 18952 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1624635492
transform 1 0 18308 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_139
timestamp 1624635492
transform 1 0 13892 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output597
timestamp 1624635492
transform -1 0 15088 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output600
timestamp 1624635492
transform -1 0 15824 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1624635492
transform 1 0 15088 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1624635492
transform -1 0 16468 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1624635492
transform 1 0 15824 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output516
timestamp 1624635492
transform -1 0 17204 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1624635492
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_175
timestamp 1624635492
transform 1 0 17204 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output485
timestamp 1624635492
transform 1 0 17940 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 18952 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1624635492
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1624635492
transform -1 0 14076 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output599
timestamp 1624635492
transform -1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1624635492
transform 1 0 14076 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1624635492
transform -1 0 15456 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1624635492
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_156
timestamp 1624635492
transform 1 0 15456 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1624635492
transform -1 0 16468 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1624635492
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_174
timestamp 1624635492
transform 1 0 17112 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output538
timestamp 1624635492
transform -1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_184
timestamp 1624635492
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 18952 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_190
timestamp 1624635492
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_139
timestamp 1624635492
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 1624635492
transform 1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1624635492
transform -1 0 14996 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_151
timestamp 1624635492
transform 1 0 14996 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1624635492
transform -1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1624635492
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1624635492
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_166
timestamp 1624635492
transform 1 0 16376 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1624635492
transform -1 0 17020 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp 1624635492
transform 1 0 17020 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _325_
timestamp 1624635492
transform -1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1624635492
transform -1 0 17664 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1624635492
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1624635492
transform 1 0 18308 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input200
timestamp 1624635492
transform -1 0 14536 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1624635492
transform 1 0 13892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1624635492
transform 1 0 14536 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139
timestamp 1624635492
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input133
timestamp 1624635492
transform -1 0 15180 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input198
timestamp 1624635492
transform -1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1624635492
transform -1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1624635492
transform 1 0 15180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1624635492
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1624635492
transform 1 0 15456 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1624635492
transform -1 0 16468 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1624635492
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1624635492
transform -1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_160
timestamp 1624635492
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_163
timestamp 1624635492
transform 1 0 16100 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1624635492
transform -1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1624635492
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_169
timestamp 1624635492
transform 1 0 16652 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1624635492
transform 1 0 17020 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1624635492
transform -1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1624635492
transform -1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1624635492
transform -1 0 18308 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1624635492
transform -1 0 17664 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_176
timestamp 1624635492
transform 1 0 17296 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_180
timestamp 1624635492
transform 1 0 17664 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_180
timestamp 1624635492
transform 1 0 17664 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 18952 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 18952 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1624635492
transform 1 0 18308 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_187
timestamp 1624635492
transform 1 0 18308 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input261
timestamp 1624635492
transform -1 0 14536 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1624635492
transform 1 0 13800 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1624635492
transform 1 0 14168 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_146
timestamp 1624635492
transform 1 0 14536 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input212
timestamp 1624635492
transform -1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1624635492
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input178
timestamp 1624635492
transform -1 0 16468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input205
timestamp 1624635492
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1624635492
transform 1 0 15824 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1624635492
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_172
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1624635492
transform -1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1624635492
transform -1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_176
timestamp 1624635492
transform 1 0 17296 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1624635492
transform 1 0 17664 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 18952 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_187
timestamp 1624635492
transform 1 0 18308 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_139
timestamp 1624635492
transform 1 0 13892 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input239
timestamp 1624635492
transform -1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1624635492
transform -1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1624635492
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_156
timestamp 1624635492
transform 1 0 15456 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input210
timestamp 1624635492
transform -1 0 16100 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1624635492
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input122
timestamp 1624635492
transform 1 0 17112 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input204
timestamp 1624635492
transform -1 0 16744 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1624635492
transform 1 0 16744 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1624635492
transform -1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_177
timestamp 1624635492
transform 1 0 17388 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_183
timestamp 1624635492
transform 1 0 17940 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 18952 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1624635492
transform 1 0 18308 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input321
timestamp 1624635492
transform -1 0 14352 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1624635492
transform 1 0 13984 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1624635492
transform 1 0 14352 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14720 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input213
timestamp 1624635492
transform -1 0 16468 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_157
timestamp 1624635492
transform 1 0 15548 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_163
timestamp 1624635492
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_167
timestamp 1624635492
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input144
timestamp 1624635492
transform -1 0 18216 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input203
timestamp 1624635492
transform -1 0 17572 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1624635492
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 18952 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1624635492
transform 1 0 18216 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1624635492
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_137
timestamp 1624635492
transform 1 0 13708 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input353
timestamp 1624635492
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input354
timestamp 1624635492
transform 1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_151
timestamp 1624635492
transform 1 0 14996 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1624635492
transform -1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_158
timestamp 1624635492
transform 1 0 15640 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_164
timestamp 1624635492
transform 1 0 16192 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1624635492
transform -1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1624635492
transform 1 0 16468 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1624635492
transform 1 0 17020 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _209_
timestamp 1624635492
transform 1 0 18032 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input211
timestamp 1624635492
transform -1 0 17664 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1624635492
transform 1 0 17664 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 18952 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1624635492
transform 1 0 18308 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input351
timestamp 1624635492
transform -1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_141
timestamp 1624635492
transform 1 0 14076 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1624635492
transform -1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1624635492
transform -1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1624635492
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1624635492
transform 1 0 15364 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1624635492
transform -1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1624635492
transform -1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_161
timestamp 1624635492
transform 1 0 15916 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_167
timestamp 1624635492
transform 1 0 16468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_172
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _129_
timestamp 1624635492
transform -1 0 18308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _290_
timestamp 1624635492
transform 1 0 17388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_176
timestamp 1624635492
transform 1 0 17296 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_180
timestamp 1624635492
transform 1 0 17664 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1624635492
transform 1 0 18308 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _303_
timestamp 1624635492
transform -1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input198_A
timestamp 1624635492
transform -1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input213_A
timestamp 1624635492
transform -1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_139
timestamp 1624635492
transform 1 0 13892 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1624635492
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_156
timestamp 1624635492
transform 1 0 15456 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1624635492
transform -1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1624635492
transform -1 0 16560 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1624635492
transform -1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1624635492
transform 1 0 16008 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1624635492
transform 1 0 16560 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1624635492
transform 1 0 17112 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _281_
timestamp 1624635492
transform 1 0 18032 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 18952 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1624635492
transform -1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1624635492
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1624635492
transform 1 0 18308 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1624635492
transform -1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input200_A
timestamp 1624635492
transform -1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input272_A
timestamp 1624635492
transform -1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_141
timestamp 1624635492
transform 1 0 14076 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_145
timestamp 1624635492
transform 1 0 14444 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1624635492
transform 1 0 14720 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_152
timestamp 1624635492
transform 1 0 15088 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_155
timestamp 1624635492
transform 1 0 15364 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _254_
timestamp 1624635492
transform 1 0 17296 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1624635492
transform -1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_165
timestamp 1624635492
transform 1 0 16284 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _224_
timestamp 1624635492
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 18952 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1624635492
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_183
timestamp 1624635492
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1624635492
transform 1 0 18308 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input212_A
timestamp 1624635492
transform -1 0 15364 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input320_A
timestamp 1624635492
transform -1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1624635492
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1624635492
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1624635492
transform 1 0 15364 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1624635492
transform -1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input178_A
timestamp 1624635492
transform -1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input205_A
timestamp 1624635492
transform -1 0 16008 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_159
timestamp 1624635492
transform 1 0 15732 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1624635492
transform 1 0 16008 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_166
timestamp 1624635492
transform 1 0 16376 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_169
timestamp 1624635492
transform 1 0 16652 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_173
timestamp 1624635492
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_176
timestamp 1624635492
transform 1 0 17296 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 18952 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1624635492
transform -1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_182
timestamp 1624635492
transform 1 0 17848 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_190
timestamp 1624635492
transform 1 0 18584 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input321_A
timestamp 1624635492
transform -1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input351_A
timestamp 1624635492
transform -1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input354_A
timestamp 1624635492
transform -1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_143
timestamp 1624635492
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1624635492
transform 1 0 14536 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1624635492
transform 1 0 15088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input204_A
timestamp 1624635492
transform -1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input210_A
timestamp 1624635492
transform -1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_158
timestamp 1624635492
transform 1 0 15640 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_162
timestamp 1624635492
transform 1 0 16008 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_165
timestamp 1624635492
transform 1 0 16284 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_174
timestamp 1624635492
transform 1 0 17112 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 18952 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1624635492
transform -1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input203_A
timestamp 1624635492
transform -1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_178
timestamp 1624635492
transform 1 0 17480 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1624635492
transform 1 0 17756 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_187
timestamp 1624635492
transform 1 0 18308 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input350_A
timestamp 1624635492
transform -1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input353_A
timestamp 1624635492
transform -1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__D
timestamp 1624635492
transform 1 0 15088 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1624635492
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1624635492
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_154
timestamp 1624635492
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _337_
timestamp 1624635492
transform -1 0 18308 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A3
timestamp 1624635492
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_164
timestamp 1624635492
transform 1 0 16192 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1624635492
transform 1 0 18308 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_137
timestamp 1624635492
transform 1 0 13708 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1624635492
transform 1 0 14260 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B1
timestamp 1624635492
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_151
timestamp 1624635492
transform 1 0 14996 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1624635492
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A2
timestamp 1624635492
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _193_
timestamp 1624635492
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 15824 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_159
timestamp 1624635492
transform 1 0 15732 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_160
timestamp 1624635492
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output444_A
timestamp 1624635492
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__C
timestamp 1624635492
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_169
timestamp 1624635492
transform 1 0 16652 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1624635492
transform 1 0 16284 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_170
timestamp 1624635492
transform 1 0 16744 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_166
timestamp 1624635492
transform 1 0 16376 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output466_A
timestamp 1624635492
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A1
timestamp 1624635492
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_172
timestamp 1624635492
transform 1 0 16928 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_176
timestamp 1624635492
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__D
timestamp 1624635492
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _261_
timestamp 1624635492
transform 1 0 18032 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 18952 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 18952 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input211_A
timestamp 1624635492
transform -1 0 17848 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output455_A
timestamp 1624635492
transform -1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_182
timestamp 1624635492
transform 1 0 17848 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_190
timestamp 1624635492
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1624635492
transform 1 0 17664 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1624635492
transform 1 0 18308 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output571_A
timestamp 1624635492
transform -1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output595_A
timestamp 1624635492
transform -1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output599_A
timestamp 1624635492
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_141
timestamp 1624635492
transform 1 0 14076 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_145
timestamp 1624635492
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1624635492
transform 1 0 14720 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_154
timestamp 1624635492
transform 1 0 15272 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output478_A
timestamp 1624635492
transform -1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output481_A
timestamp 1624635492
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output483_A
timestamp 1624635492
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_158
timestamp 1624635492
transform 1 0 15640 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_161
timestamp 1624635492
transform 1 0 15916 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_167
timestamp 1624635492
transform 1 0 16468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_174
timestamp 1624635492
transform 1 0 17112 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _302_
timestamp 1624635492
transform -1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 18952 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output475_A
timestamp 1624635492
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1624635492
transform 1 0 17664 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_187
timestamp 1624635492
transform 1 0 18308 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output597_A
timestamp 1624635492
transform 1 0 15088 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_154
timestamp 1624635492
transform 1 0 15272 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output480_A
timestamp 1624635492
transform -1 0 17388 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output489_A
timestamp 1624635492
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output494_A
timestamp 1624635492
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_162
timestamp 1624635492
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_165
timestamp 1624635492
transform 1 0 16284 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1624635492
transform 1 0 16836 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 18952 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output476_A
timestamp 1624635492
transform 1 0 17756 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1624635492
transform 1 0 17388 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_183
timestamp 1624635492
transform 1 0 17940 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1624635492
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1624635492
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output516_A
timestamp 1624635492
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1624635492
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output485_A
timestamp 1624635492
transform -1 0 18308 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_177
timestamp 1624635492
transform 1 0 17388 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1624635492
transform 1 0 18308 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_138
timestamp 1624635492
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1624635492
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1624635492
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_168
timestamp 1624635492
transform 1 0 16560 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_176
timestamp 1624635492
transform 1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 18952 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__CLK
timestamp 1624635492
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_adc.COMP_clk
timestamp 1624635492
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1624635492
transform 1 0 17756 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1624635492
transform 1 0 18308 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1624635492
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1624635492
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1624635492
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1624635492
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1624635492
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _125_
timestamp 1624635492
transform -1 0 18308 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _274_
timestamp 1624635492
transform 1 0 18032 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 18952 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 18952 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1624635492
transform 1 0 18308 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1624635492
transform 1 0 17664 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1624635492
transform 1 0 18308 0 -1 16864
box -38 -48 406 592
use ACMP  adc.COMP
timestamp 1626122236
transform 1 0 22000 0 1 2000
box 0 0 12564 14476
use sky130_fd_sc_hd__decap_4  FILLER_2_400
timestamp 1624635492
transform 1 0 37904 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_400
timestamp 1624635492
transform 1 0 37904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_400
timestamp 1624635492
transform 1 0 37904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1624635492
transform 1 0 37628 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1624635492
transform 1 0 37628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1624635492
transform 1 0 37628 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_408
timestamp 1624635492
transform 1 0 38640 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_408
timestamp 1624635492
transform 1 0 38640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_408
timestamp 1624635492
transform 1 0 38640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output493
timestamp 1624635492
transform -1 0 38640 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output491
timestamp 1624635492
transform -1 0 38640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output486
timestamp 1624635492
transform -1 0 38640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_400
timestamp 1624635492
transform 1 0 37904 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_400
timestamp 1624635492
transform 1 0 37904 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1624635492
transform 1 0 37628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1624635492
transform 1 0 37628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_408
timestamp 1624635492
transform 1 0 38640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_408
timestamp 1624635492
transform 1 0 38640 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output502
timestamp 1624635492
transform -1 0 38640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output498
timestamp 1624635492
transform -1 0 38640 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_400
timestamp 1624635492
transform 1 0 37904 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_400
timestamp 1624635492
transform 1 0 37904 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1624635492
transform 1 0 37628 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1624635492
transform 1 0 37628 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_408
timestamp 1624635492
transform 1 0 38640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_408
timestamp 1624635492
transform 1 0 38640 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output518
timestamp 1624635492
transform -1 0 38640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output509
timestamp 1624635492
transform -1 0 38640 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1624635492
transform -1 0 38180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1624635492
transform -1 0 38180 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1624635492
transform 1 0 37628 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1624635492
transform 1 0 37628 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1624635492
transform 1 0 37628 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _188_
timestamp 1624635492
transform -1 0 38180 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1624635492
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1624635492
transform 1 0 38180 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1624635492
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 1624635492
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1624635492
transform 1 0 38548 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _217_
timestamp 1624635492
transform 1 0 38548 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input109
timestamp 1624635492
transform -1 0 38180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 1624635492
transform -1 0 38180 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1624635492
transform 1 0 37628 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1624635492
transform 1 0 37628 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1624635492
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1624635492
transform 1 0 38180 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input216
timestamp 1624635492
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1624635492
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input230
timestamp 1624635492
transform 1 0 37904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input218
timestamp 1624635492
transform -1 0 38180 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1624635492
transform 1 0 37628 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1624635492
transform 1 0 37628 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1624635492
transform 1 0 37628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _319_
timestamp 1624635492
transform -1 0 38180 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1624635492
transform 1 0 38180 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1624635492
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_403
timestamp 1624635492
transform 1 0 38180 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input238
timestamp 1624635492
transform 1 0 38548 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input226
timestamp 1624635492
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _157_
timestamp 1624635492
transform 1 0 38732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input242
timestamp 1624635492
transform 1 0 37904 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1624635492
transform 1 0 37628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1624635492
transform 1 0 37628 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _327_
timestamp 1624635492
transform -1 0 38180 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_409
timestamp 1624635492
transform 1 0 38732 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1624635492
transform 1 0 38180 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_409
timestamp 1624635492
transform 1 0 38732 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1624635492
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1624635492
transform -1 0 38732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1624635492
transform -1 0 38732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input230_A
timestamp 1624635492
transform -1 0 38088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_278
timestamp 1624635492
transform 1 0 37628 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1624635492
transform 1 0 37628 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1624635492
transform 1 0 37628 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _257_
timestamp 1624635492
transform 1 0 37904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 38180 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_408
timestamp 1624635492
transform 1 0 38640 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_402
timestamp 1624635492
transform 1 0 38088 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_409
timestamp 1624635492
transform 1 0 38732 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1624635492
transform 1 0 38180 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_409
timestamp 1624635492
transform 1 0 38732 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1624635492
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input238_A
timestamp 1624635492
transform -1 0 38640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input218_A
timestamp 1624635492
transform -1 0 38732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1624635492
transform -1 0 38732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input242_A
timestamp 1624635492
transform -1 0 38088 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_282
timestamp 1624635492
transform 1 0 37628 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_280
timestamp 1624635492
transform 1 0 37628 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _236_
timestamp 1624635492
transform 1 0 37904 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_409
timestamp 1624635492
transform 1 0 38732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1624635492
transform 1 0 38180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_402
timestamp 1624635492
transform 1 0 38088 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output493_A
timestamp 1624635492
transform -1 0 38732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output491_A
timestamp 1624635492
transform 1 0 38640 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_400
timestamp 1624635492
transform 1 0 37904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_400
timestamp 1624635492
transform 1 0 37904 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_286
timestamp 1624635492
transform 1 0 37628 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_284
timestamp 1624635492
transform 1 0 37628 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_404
timestamp 1624635492
transform 1 0 38272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output518_A
timestamp 1624635492
transform 1 0 38088 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_400
timestamp 1624635492
transform 1 0 37904 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_400
timestamp 1624635492
transform 1 0 37904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_400
timestamp 1624635492
transform 1 0 37904 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_292
timestamp 1624635492
transform 1 0 37628 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_290
timestamp 1624635492
transform 1 0 37628 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_288
timestamp 1624635492
transform 1 0 37628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_422
timestamp 1624635492
transform 1 0 39928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1624635492
transform 1 0 39376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output486_A
timestamp 1624635492
transform -1 0 39928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output487
timestamp 1624635492
transform -1 0 39376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_435
timestamp 1624635492
transform 1 0 41124 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_427
timestamp 1624635492
transform 1 0 40388 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output490
timestamp 1624635492
transform -1 0 41124 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1528
timestamp 1624635492
transform 1 0 40296 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1624635492
transform 1 0 41860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output496
timestamp 1624635492
transform -1 0 42596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output492
timestamp 1624635492
transform -1 0 41860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_456
timestamp 1624635492
transform 1 0 43056 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_451
timestamp 1624635492
transform 1 0 42596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output500
timestamp 1624635492
transform -1 0 43792 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1529
timestamp 1624635492
transform 1 0 42964 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1624635492
transform 1 0 44528 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_464
timestamp 1624635492
transform 1 0 43792 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output507
timestamp 1624635492
transform -1 0 44528 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_485
timestamp 1624635492
transform 1 0 45724 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1624635492
transform 1 0 45264 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output511
timestamp 1624635492
transform -1 0 45264 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1530
timestamp 1624635492
transform 1 0 45632 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_493
timestamp 1624635492
transform 1 0 46460 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output529
timestamp 1624635492
transform -1 0 47196 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output522
timestamp 1624635492
transform -1 0 46460 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_509
timestamp 1624635492
transform 1 0 47932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_501
timestamp 1624635492
transform 1 0 47196 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output532
timestamp 1624635492
transform -1 0 47932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_522
timestamp 1624635492
transform 1 0 49128 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_514
timestamp 1624635492
transform 1 0 48392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output537
timestamp 1624635492
transform -1 0 49128 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1531
timestamp 1624635492
transform 1 0 48300 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_538
timestamp 1624635492
transform 1 0 50600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_530
timestamp 1624635492
transform 1 0 49864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output541
timestamp 1624635492
transform -1 0 50600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output540
timestamp 1624635492
transform -1 0 49864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1624635492
transform 1 0 51060 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1532
timestamp 1624635492
transform 1 0 50968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_422
timestamp 1624635492
transform 1 0 39928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1624635492
transform 1 0 39376 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_416
timestamp 1624635492
transform 1 0 39376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1624635492
transform -1 0 39928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output497
timestamp 1624635492
transform -1 0 39376 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output495
timestamp 1624635492
transform -1 0 39376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output488
timestamp 1624635492
transform -1 0 40112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_435
timestamp 1624635492
transform 1 0 41124 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_427
timestamp 1624635492
transform 1 0 40388 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_432
timestamp 1624635492
transform 1 0 40848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1624635492
transform 1 0 40112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output514
timestamp 1624635492
transform -1 0 41124 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output499
timestamp 1624635492
transform -1 0 40848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1544
timestamp 1624635492
transform 1 0 40296 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_448
timestamp 1624635492
transform 1 0 42320 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_443
timestamp 1624635492
transform 1 0 41860 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_448
timestamp 1624635492
transform 1 0 42320 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_440
timestamp 1624635492
transform 1 0 41584 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output517
timestamp 1624635492
transform -1 0 42320 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output508
timestamp 1624635492
transform -1 0 42320 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output504
timestamp 1624635492
transform -1 0 41584 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_456
timestamp 1624635492
transform 1 0 43056 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_455
timestamp 1624635492
transform 1 0 42964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output528
timestamp 1624635492
transform -1 0 43700 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output525
timestamp 1624635492
transform -1 0 43792 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output521
timestamp 1624635492
transform -1 0 43056 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1539
timestamp 1624635492
transform 1 0 42872 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1624635492
transform 1 0 44528 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_464
timestamp 1624635492
transform 1 0 43792 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_471
timestamp 1624635492
transform 1 0 44436 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_463
timestamp 1624635492
transform 1 0 43700 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output533
timestamp 1624635492
transform -1 0 44528 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output531
timestamp 1624635492
transform -1 0 44436 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_486
timestamp 1624635492
transform 1 0 45816 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_482
timestamp 1624635492
transform 1 0 45448 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_478
timestamp 1624635492
transform 1 0 45080 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_479
timestamp 1624635492
transform 1 0 45172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1624635492
transform -1 0 45816 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1624635492
transform -1 0 45080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output536
timestamp 1624635492
transform -1 0 45908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output534
timestamp 1624635492
transform -1 0 45172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1545
timestamp 1624635492
transform 1 0 45540 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_498
timestamp 1624635492
transform 1 0 46920 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_495
timestamp 1624635492
transform 1 0 46644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1624635492
transform 1 0 45908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output543
timestamp 1624635492
transform -1 0 46920 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output542
timestamp 1624635492
transform -1 0 47380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output539
timestamp 1624635492
transform -1 0 46644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_508
timestamp 1624635492
transform 1 0 47840 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1624635492
transform 1 0 48208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_503
timestamp 1624635492
transform 1 0 47380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output545
timestamp 1624635492
transform -1 0 47840 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1624635492
transform 1 0 48208 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1540
timestamp 1624635492
transform 1 0 48116 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_522
timestamp 1624635492
transform 1 0 49128 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_515
timestamp 1624635492
transform 1 0 48484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_520
timestamp 1624635492
transform 1 0 48944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output548
timestamp 1624635492
transform -1 0 49680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output546
timestamp 1624635492
transform -1 0 48944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input140
timestamp 1624635492
transform 1 0 48852 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_536
timestamp 1624635492
transform 1 0 50416 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_529
timestamp 1624635492
transform 1 0 49772 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1624635492
transform 1 0 50416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_528
timestamp 1624635492
transform 1 0 49680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output551
timestamp 1624635492
transform -1 0 50416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input145
timestamp 1624635492
transform -1 0 50416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1624635492
transform -1 0 49772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_541
timestamp 1624635492
transform 1 0 50876 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_544
timestamp 1624635492
transform 1 0 51152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output552
timestamp 1624635492
transform -1 0 51152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1624635492
transform -1 0 51520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1546
timestamp 1624635492
transform 1 0 50784 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_416
timestamp 1624635492
transform 1 0 39376 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output503
timestamp 1624635492
transform -1 0 40112 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output501
timestamp 1624635492
transform -1 0 39376 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_432
timestamp 1624635492
transform 1 0 40848 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_424
timestamp 1624635492
transform 1 0 40112 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output506
timestamp 1624635492
transform -1 0 40848 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_448
timestamp 1624635492
transform 1 0 42320 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_440
timestamp 1624635492
transform 1 0 41584 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output519
timestamp 1624635492
transform -1 0 42320 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output512
timestamp 1624635492
transform -1 0 41584 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_455
timestamp 1624635492
transform 1 0 42964 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output530
timestamp 1624635492
transform -1 0 43700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1550
timestamp 1624635492
transform 1 0 42872 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_463
timestamp 1624635492
transform 1 0 43700 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output535
timestamp 1624635492
transform -1 0 44804 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_482
timestamp 1624635492
transform 1 0 45448 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_475
timestamp 1624635492
transform 1 0 44804 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input124
timestamp 1624635492
transform -1 0 46092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1624635492
transform -1 0 45448 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_496
timestamp 1624635492
transform 1 0 46736 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1624635492
transform 1 0 46092 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input128
timestamp 1624635492
transform -1 0 46736 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1624635492
transform 1 0 48208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_503
timestamp 1624635492
transform 1 0 47380 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input131
timestamp 1624635492
transform -1 0 47380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1551
timestamp 1624635492
transform 1 0 48116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_519
timestamp 1624635492
transform 1 0 48852 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1624635492
transform 1 0 49220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1624635492
transform -1 0 48852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_533
timestamp 1624635492
transform 1 0 50140 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_526
timestamp 1624635492
transform 1 0 49496 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1624635492
transform -1 0 50784 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input146
timestamp 1624635492
transform 1 0 49864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_540
timestamp 1624635492
transform 1 0 50784 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input149
timestamp 1624635492
transform -1 0 51428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_422
timestamp 1624635492
transform 1 0 39928 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1624635492
transform 1 0 39376 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_adc.COMP_INP
timestamp 1624635492
transform -1 0 39928 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output510
timestamp 1624635492
transform -1 0 39376 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_435
timestamp 1624635492
transform 1 0 41124 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_427
timestamp 1624635492
transform 1 0 40388 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output526
timestamp 1624635492
transform -1 0 41124 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1555
timestamp 1624635492
transform 1 0 40296 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_448
timestamp 1624635492
transform 1 0 42320 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_443
timestamp 1624635492
transform 1 0 41860 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output523
timestamp 1624635492
transform -1 0 42320 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_461
timestamp 1624635492
transform 1 0 43516 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_455
timestamp 1624635492
transform 1 0 42964 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1624635492
transform -1 0 43516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 1624635492
transform -1 0 42964 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_468
timestamp 1624635492
transform 1 0 44160 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 1624635492
transform -1 0 44804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _269_
timestamp 1624635492
transform 1 0 43884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_484
timestamp 1624635492
transform 1 0 45632 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_475
timestamp 1624635492
transform 1 0 44804 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1556
timestamp 1624635492
transform 1 0 45540 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_497
timestamp 1624635492
transform 1 0 46828 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_491
timestamp 1624635492
transform 1 0 46276 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1624635492
transform -1 0 46828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input130
timestamp 1624635492
transform -1 0 46276 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_511
timestamp 1624635492
transform 1 0 48116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_504
timestamp 1624635492
transform 1 0 47472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input139
timestamp 1624635492
transform -1 0 48116 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input136
timestamp 1624635492
transform -1 0 47472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_525
timestamp 1624635492
transform 1 0 49404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_518
timestamp 1624635492
transform 1 0 48760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input262
timestamp 1624635492
transform 1 0 49128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input253
timestamp 1624635492
transform 1 0 48484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_532
timestamp 1624635492
transform 1 0 50048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input266
timestamp 1624635492
transform -1 0 50048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_541
timestamp 1624635492
transform 1 0 50876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input274
timestamp 1624635492
transform -1 0 51520 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1557
timestamp 1624635492
transform 1 0 50784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_416
timestamp 1624635492
transform 1 0 39376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output515
timestamp 1624635492
transform -1 0 40112 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output513
timestamp 1624635492
transform -1 0 39376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_432
timestamp 1624635492
transform 1 0 40848 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_424
timestamp 1624635492
transform 1 0 40112 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output520
timestamp 1624635492
transform -1 0 40848 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_447
timestamp 1624635492
transform 1 0 42228 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_440
timestamp 1624635492
transform 1 0 41584 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output524
timestamp 1624635492
transform -1 0 41584 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1624635492
transform -1 0 42228 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_455
timestamp 1624635492
transform 1 0 42964 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_453
timestamp 1624635492
transform 1 0 42780 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1624635492
transform -1 0 43608 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1561
timestamp 1624635492
transform 1 0 42872 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_469
timestamp 1624635492
transform 1 0 44252 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_462
timestamp 1624635492
transform 1 0 43608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input121
timestamp 1624635492
transform 1 0 44620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1624635492
transform -1 0 44252 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_483
timestamp 1624635492
transform 1 0 45540 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_476
timestamp 1624635492
transform 1 0 44896 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input129
timestamp 1624635492
transform -1 0 45540 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_497
timestamp 1624635492
transform 1 0 46828 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_490
timestamp 1624635492
transform 1 0 46184 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input135
timestamp 1624635492
transform -1 0 46828 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input134
timestamp 1624635492
transform -1 0 46184 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1624635492
transform 1 0 48208 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_510
timestamp 1624635492
transform 1 0 48024 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_504
timestamp 1624635492
transform 1 0 47472 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1624635492
transform -1 0 47472 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1562
timestamp 1624635492
transform 1 0 48116 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_519
timestamp 1624635492
transform 1 0 48852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input267
timestamp 1624635492
transform -1 0 48852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _231_
timestamp 1624635492
transform -1 0 49680 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_535
timestamp 1624635492
transform 1 0 50324 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_528
timestamp 1624635492
transform 1 0 49680 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input268
timestamp 1624635492
transform 1 0 50048 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_543
timestamp 1624635492
transform 1 0 51060 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_2  _077_
timestamp 1624635492
transform 1 0 51152 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_422
timestamp 1624635492
transform 1 0 39928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_415
timestamp 1624635492
transform 1 0 39284 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1624635492
transform -1 0 39928 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _294_
timestamp 1624635492
transform 1 0 39008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_435
timestamp 1624635492
transform 1 0 41124 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_431
timestamp 1624635492
transform 1 0 40756 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_427
timestamp 1624635492
transform 1 0 40388 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1624635492
transform -1 0 41124 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1566
timestamp 1624635492
transform 1 0 40296 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_442
timestamp 1624635492
transform 1 0 41768 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1624635492
transform -1 0 42412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1624635492
transform -1 0 41768 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_456
timestamp 1624635492
transform 1 0 43056 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_449
timestamp 1624635492
transform 1 0 42412 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1624635492
transform -1 0 43700 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 1624635492
transform 1 0 42780 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_470
timestamp 1624635492
transform 1 0 44344 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_463
timestamp 1624635492
transform 1 0 43700 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input125
timestamp 1624635492
transform -1 0 44344 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_486
timestamp 1624635492
transform 1 0 45816 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_477
timestamp 1624635492
transform 1 0 44988 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1624635492
transform -1 0 45816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input127
timestamp 1624635492
transform -1 0 44988 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1567
timestamp 1624635492
transform 1 0 45540 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_497
timestamp 1624635492
transform 1 0 46828 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input245
timestamp 1624635492
transform -1 0 46828 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_511
timestamp 1624635492
transform 1 0 48116 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_504
timestamp 1624635492
transform 1 0 47472 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input260
timestamp 1624635492
transform -1 0 48116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input254
timestamp 1624635492
transform 1 0 47196 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_525
timestamp 1624635492
transform 1 0 49404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_518
timestamp 1624635492
transform 1 0 48760 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input269
timestamp 1624635492
transform -1 0 49404 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input265
timestamp 1624635492
transform -1 0 48760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_532
timestamp 1624635492
transform 1 0 50048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input270
timestamp 1624635492
transform -1 0 50048 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_541
timestamp 1624635492
transform 1 0 50876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input276
timestamp 1624635492
transform -1 0 51520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1568
timestamp 1624635492
transform 1 0 50784 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_417
timestamp 1624635492
transform 1 0 39468 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_410
timestamp 1624635492
transform 1 0 38824 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_419
timestamp 1624635492
transform 1 0 39652 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_410
timestamp 1624635492
transform 1 0 38824 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1624635492
transform -1 0 39468 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _108_
timestamp 1624635492
transform 1 0 39376 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_429
timestamp 1624635492
transform 1 0 40572 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_425
timestamp 1624635492
transform 1 0 40204 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_433
timestamp 1624635492
transform 1 0 40940 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_426
timestamp 1624635492
transform 1 0 40296 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1624635492
transform -1 0 40572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 1624635492
transform 1 0 40664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1577
timestamp 1624635492
transform 1 0 40296 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _121_
timestamp 1624635492
transform -1 0 40296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_447
timestamp 1624635492
transform 1 0 42228 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_440
timestamp 1624635492
transform 1 0 41584 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_448
timestamp 1624635492
transform 1 0 42320 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_441
timestamp 1624635492
transform 1 0 41676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_437
timestamp 1624635492
transform 1 0 41308 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1624635492
transform -1 0 42228 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 1624635492
transform 1 0 41308 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1624635492
transform 1 0 42044 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 1624635492
transform 1 0 41400 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_458
timestamp 1624635492
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_454
timestamp 1624635492
transform 1 0 42872 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_455
timestamp 1624635492
transform 1 0 42964 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input224
timestamp 1624635492
transform -1 0 43608 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input123
timestamp 1624635492
transform -1 0 42872 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input119
timestamp 1624635492
transform 1 0 43332 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1572
timestamp 1624635492
transform 1 0 42872 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_469
timestamp 1624635492
transform 1 0 44252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_462
timestamp 1624635492
transform 1 0 43608 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_469
timestamp 1624635492
transform 1 0 44252 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_462
timestamp 1624635492
transform 1 0 43608 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input243
timestamp 1624635492
transform -1 0 44896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input231
timestamp 1624635492
transform 1 0 43976 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input132
timestamp 1624635492
transform -1 0 44896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input126
timestamp 1624635492
transform 1 0 43976 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_484
timestamp 1624635492
transform 1 0 45632 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_482
timestamp 1624635492
transform 1 0 45448 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_476
timestamp 1624635492
transform 1 0 44896 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_483
timestamp 1624635492
transform 1 0 45540 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_476
timestamp 1624635492
transform 1 0 44896 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input240
timestamp 1624635492
transform -1 0 45540 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1578
timestamp 1624635492
transform 1 0 45540 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_498
timestamp 1624635492
transform 1 0 46920 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_491
timestamp 1624635492
transform 1 0 46276 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_497
timestamp 1624635492
transform 1 0 46828 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_490
timestamp 1624635492
transform 1 0 46184 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input263
timestamp 1624635492
transform 1 0 46644 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input257
timestamp 1624635492
transform 1 0 46000 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input251
timestamp 1624635492
transform -1 0 46828 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input248
timestamp 1624635492
transform -1 0 46184 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_511
timestamp 1624635492
transform 1 0 48116 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1624635492
transform 1 0 47564 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_510
timestamp 1624635492
transform 1 0 48024 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_504
timestamp 1624635492
transform 1 0 47472 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1624635492
transform -1 0 48116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1624635492
transform -1 0 48392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input264
timestamp 1624635492
transform -1 0 47564 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input259
timestamp 1624635492
transform 1 0 47196 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1573
timestamp 1624635492
transform 1 0 48116 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_523
timestamp 1624635492
transform 1 0 49220 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_517
timestamp 1624635492
transform 1 0 48668 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_520
timestamp 1624635492
transform 1 0 48944 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_514
timestamp 1624635492
transform 1 0 48392 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1624635492
transform -1 0 49220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1624635492
transform -1 0 48668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1624635492
transform -1 0 49496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1624635492
transform -1 0 48944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_535
timestamp 1624635492
transform 1 0 50324 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_529
timestamp 1624635492
transform 1 0 49772 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_535
timestamp 1624635492
transform 1 0 50324 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_526
timestamp 1624635492
transform 1 0 49496 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1624635492
transform -1 0 50324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1624635492
transform -1 0 49772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input271
timestamp 1624635492
transform -1 0 50324 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_543
timestamp 1624635492
transform 1 0 51060 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_539
timestamp 1624635492
transform 1 0 50692 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_542
timestamp 1624635492
transform 1 0 50968 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input147_A
timestamp 1624635492
transform -1 0 51060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input273
timestamp 1624635492
transform -1 0 50968 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1579
timestamp 1624635492
transform 1 0 50784 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_417
timestamp 1624635492
transform 1 0 39468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_410
timestamp 1624635492
transform 1 0 38824 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1624635492
transform -1 0 40112 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1624635492
transform -1 0 39468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_434
timestamp 1624635492
transform 1 0 41032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_430
timestamp 1624635492
transform 1 0 40664 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_424
timestamp 1624635492
transform 1 0 40112 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1624635492
transform 1 0 40756 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_448
timestamp 1624635492
transform 1 0 42320 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_441
timestamp 1624635492
transform 1 0 41676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input222
timestamp 1624635492
transform -1 0 42320 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input221
timestamp 1624635492
transform 1 0 41400 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_455
timestamp 1624635492
transform 1 0 42964 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input227
timestamp 1624635492
transform 1 0 43332 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1583
timestamp 1624635492
transform 1 0 42872 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_469
timestamp 1624635492
transform 1 0 44252 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_462
timestamp 1624635492
transform 1 0 43608 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input252
timestamp 1624635492
transform -1 0 44896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input236
timestamp 1624635492
transform -1 0 44252 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_483
timestamp 1624635492
transform 1 0 45540 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_476
timestamp 1624635492
transform 1 0 44896 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input258
timestamp 1624635492
transform -1 0 45540 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_495
timestamp 1624635492
transform 1 0 46644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_489
timestamp 1624635492
transform 1 0 46092 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1624635492
transform -1 0 47196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1624635492
transform -1 0 46644 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1624635492
transform -1 0 46092 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_507
timestamp 1624635492
transform 1 0 47748 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_501
timestamp 1624635492
transform 1 0 47196 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1624635492
transform -1 0 48392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1624635492
transform -1 0 47748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1584
timestamp 1624635492
transform 1 0 48116 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_520
timestamp 1624635492
transform 1 0 48944 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_514
timestamp 1624635492
transform 1 0 48392 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1624635492
transform -1 0 49496 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1624635492
transform -1 0 48944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_538
timestamp 1624635492
transform 1 0 50600 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_532
timestamp 1624635492
transform 1 0 50048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_526
timestamp 1624635492
transform 1 0 49496 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input266_A
timestamp 1624635492
transform -1 0 50600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input146_A
timestamp 1624635492
transform -1 0 50048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_544
timestamp 1624635492
transform 1 0 51152 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input270_A
timestamp 1624635492
transform -1 0 51152 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_417
timestamp 1624635492
transform 1 0 39468 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_410
timestamp 1624635492
transform 1 0 38824 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1624635492
transform -1 0 39468 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_434
timestamp 1624635492
transform 1 0 41032 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_427
timestamp 1624635492
transform 1 0 40388 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_425
timestamp 1624635492
transform 1 0 40204 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1624635492
transform -1 0 41032 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1588
timestamp 1624635492
transform 1 0 40296 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_448
timestamp 1624635492
transform 1 0 42320 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_441
timestamp 1624635492
transform 1 0 41676 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input225
timestamp 1624635492
transform -1 0 42320 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input223
timestamp 1624635492
transform -1 0 41676 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_455
timestamp 1624635492
transform 1 0 42964 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input241
timestamp 1624635492
transform -1 0 43608 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input237
timestamp 1624635492
transform -1 0 42964 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_469
timestamp 1624635492
transform 1 0 44252 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_462
timestamp 1624635492
transform 1 0 43608 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input256
timestamp 1624635492
transform 1 0 44620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input255
timestamp 1624635492
transform 1 0 43976 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_486
timestamp 1624635492
transform 1 0 45816 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_482
timestamp 1624635492
transform 1 0 45448 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_476
timestamp 1624635492
transform 1 0 44896 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1624635492
transform -1 0 45816 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1589
timestamp 1624635492
transform 1 0 45540 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_498
timestamp 1624635492
transform 1 0 46920 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_492
timestamp 1624635492
transform 1 0 46368 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1624635492
transform -1 0 46920 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1624635492
transform -1 0 46368 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_510
timestamp 1624635492
transform 1 0 48024 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_504
timestamp 1624635492
transform 1 0 47472 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input251_A
timestamp 1624635492
transform -1 0 48024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input248_A
timestamp 1624635492
transform -1 0 47472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_522
timestamp 1624635492
transform 1 0 49128 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_516
timestamp 1624635492
transform 1 0 48576 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input262_A
timestamp 1624635492
transform -1 0 49128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input253_A
timestamp 1624635492
transform -1 0 48576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_534
timestamp 1624635492
transform 1 0 50232 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_528
timestamp 1624635492
transform 1 0 49680 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input268_A
timestamp 1624635492
transform -1 0 50232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input267_A
timestamp 1624635492
transform -1 0 49680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_543
timestamp 1624635492
transform 1 0 51060 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input273_A
timestamp 1624635492
transform -1 0 51060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1590
timestamp 1624635492
transform 1 0 50784 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_417
timestamp 1624635492
transform 1 0 39468 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_410
timestamp 1624635492
transform 1 0 38824 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input220
timestamp 1624635492
transform -1 0 40112 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input219
timestamp 1624635492
transform -1 0 39468 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_431
timestamp 1624635492
transform 1 0 40756 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_424
timestamp 1624635492
transform 1 0 40112 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input232
timestamp 1624635492
transform 1 0 40480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_448
timestamp 1624635492
transform 1 0 42320 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_441
timestamp 1624635492
transform 1 0 41676 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_437
timestamp 1624635492
transform 1 0 41308 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input247
timestamp 1624635492
transform -1 0 42320 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input234
timestamp 1624635492
transform 1 0 41400 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_455
timestamp 1624635492
transform 1 0 42964 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input249
timestamp 1624635492
transform -1 0 43608 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1594
timestamp 1624635492
transform 1 0 42872 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_468
timestamp 1624635492
transform 1 0 44160 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_462
timestamp 1624635492
transform 1 0 43608 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1624635492
transform -1 0 44712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1624635492
transform -1 0 44160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_486
timestamp 1624635492
transform 1 0 45816 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_480
timestamp 1624635492
transform 1 0 45264 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_474
timestamp 1624635492
transform 1 0 44712 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1624635492
transform -1 0 45816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1624635492
transform -1 0 45264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_498
timestamp 1624635492
transform 1 0 46920 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_492
timestamp 1624635492
transform 1 0 46368 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input245_A
timestamp 1624635492
transform -1 0 46920 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input241_A
timestamp 1624635492
transform -1 0 46368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_510
timestamp 1624635492
transform 1 0 48024 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_504
timestamp 1624635492
transform 1 0 47472 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input260_A
timestamp 1624635492
transform -1 0 48392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input254_A
timestamp 1624635492
transform -1 0 47472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1595
timestamp 1624635492
transform 1 0 48116 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_520
timestamp 1624635492
transform 1 0 48944 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_514
timestamp 1624635492
transform 1 0 48392 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input269_A
timestamp 1624635492
transform -1 0 49496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input265_A
timestamp 1624635492
transform -1 0 48944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_536
timestamp 1624635492
transform 1 0 50416 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_526
timestamp 1624635492
transform 1 0 49496 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A2
timestamp 1624635492
transform 1 0 50232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_542
timestamp 1624635492
transform 1 0 50968 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A1
timestamp 1624635492
transform 1 0 50784 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _113_
timestamp 1624635492
transform 1 0 51336 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_419
timestamp 1624635492
transform 1 0 39652 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_412
timestamp 1624635492
transform 1 0 39008 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input229
timestamp 1624635492
transform -1 0 39652 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_429
timestamp 1624635492
transform 1 0 40572 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_425
timestamp 1624635492
transform 1 0 40204 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1624635492
transform -1 0 40572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input235
timestamp 1624635492
transform 1 0 41124 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1599
timestamp 1624635492
transform 1 0 40296 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_444
timestamp 1624635492
transform 1 0 41952 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_438
timestamp 1624635492
transform 1 0 41400 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1624635492
transform -1 0 42504 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1624635492
transform -1 0 41952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_456
timestamp 1624635492
transform 1 0 43056 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_450
timestamp 1624635492
transform 1 0 42504 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1624635492
transform -1 0 43608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1624635492
transform -1 0 43056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_468
timestamp 1624635492
transform 1 0 44160 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_462
timestamp 1624635492
transform 1 0 43608 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input224_A
timestamp 1624635492
transform -1 0 44712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1624635492
transform -1 0 44160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_486
timestamp 1624635492
transform 1 0 45816 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_482
timestamp 1624635492
transform 1 0 45448 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_474
timestamp 1624635492
transform 1 0 44712 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input240_A
timestamp 1624635492
transform -1 0 45816 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1600
timestamp 1624635492
transform 1 0 45540 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_498
timestamp 1624635492
transform 1 0 46920 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_492
timestamp 1624635492
transform 1 0 46368 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input258_A
timestamp 1624635492
transform -1 0 46920 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input252_A
timestamp 1624635492
transform -1 0 46368 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_510
timestamp 1624635492
transform 1 0 48024 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_504
timestamp 1624635492
transform 1 0 47472 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input264_A
timestamp 1624635492
transform -1 0 48024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input259_A
timestamp 1624635492
transform -1 0 47472 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_522
timestamp 1624635492
transform 1 0 49128 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_516
timestamp 1624635492
transform 1 0 48576 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output536_A
timestamp 1624635492
transform -1 0 49128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output526_A
timestamp 1624635492
transform 1 0 48392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_534
timestamp 1624635492
transform 1 0 50232 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1624635492
transform 1 0 49680 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output541_A
timestamp 1624635492
transform 1 0 50048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output540_A
timestamp 1624635492
transform 1 0 49496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_543
timestamp 1624635492
transform 1 0 51060 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A3
timestamp 1624635492
transform 1 0 50876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1601
timestamp 1624635492
transform 1 0 50784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_417
timestamp 1624635492
transform 1 0 39468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_410
timestamp 1624635492
transform 1 0 38824 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input244
timestamp 1624635492
transform -1 0 40112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input233
timestamp 1624635492
transform -1 0 39468 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_434
timestamp 1624635492
transform 1 0 41032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_430
timestamp 1624635492
transform 1 0 40664 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_424
timestamp 1624635492
transform 1 0 40112 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input246
timestamp 1624635492
transform -1 0 41032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_446
timestamp 1624635492
transform 1 0 42136 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_440
timestamp 1624635492
transform 1 0 41584 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1624635492
transform -1 0 42136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1624635492
transform -1 0 41584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_457
timestamp 1624635492
transform 1 0 43148 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input222_A
timestamp 1624635492
transform -1 0 43700 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1624635492
transform -1 0 43148 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1605
timestamp 1624635492
transform 1 0 42872 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_469
timestamp 1624635492
transform 1 0 44252 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_463
timestamp 1624635492
transform 1 0 43700 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input236_A
timestamp 1624635492
transform -1 0 44804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input231_A
timestamp 1624635492
transform -1 0 44252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_485
timestamp 1624635492
transform 1 0 45724 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_481
timestamp 1624635492
transform 1 0 45356 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_475
timestamp 1624635492
transform 1 0 44804 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input257_A
timestamp 1624635492
transform -1 0 46000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input243_A
timestamp 1624635492
transform -1 0 45356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_495
timestamp 1624635492
transform 1 0 46644 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_492
timestamp 1624635492
transform 1 0 46368 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_488
timestamp 1624635492
transform 1 0 46000 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output511_A
timestamp 1624635492
transform -1 0 47196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input263_A
timestamp 1624635492
transform -1 0 46644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1624635492
transform 1 0 48208 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_507
timestamp 1624635492
transform 1 0 47748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_501
timestamp 1624635492
transform 1 0 47196 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output530_A
timestamp 1624635492
transform -1 0 47748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1606
timestamp 1624635492
transform 1 0 48116 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_524
timestamp 1624635492
transform 1 0 49312 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_518
timestamp 1624635492
transform 1 0 48760 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output546_A
timestamp 1624635492
transform -1 0 49312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output537_A
timestamp 1624635492
transform 1 0 48576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_536
timestamp 1624635492
transform 1 0 50416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_530
timestamp 1624635492
transform 1 0 49864 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output551_A
timestamp 1624635492
transform -1 0 50416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output548_A
timestamp 1624635492
transform 1 0 49680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_421
timestamp 1624635492
transform 1 0 39836 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_415
timestamp 1624635492
transform 1 0 39284 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_422
timestamp 1624635492
transform 1 0 39928 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1624635492
transform 1 0 39376 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_410
timestamp 1624635492
transform 1 0 38824 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1624635492
transform -1 0 39836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1624635492
transform -1 0 39928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1624635492
transform -1 0 39284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_adc.COMP_INN
timestamp 1624635492
transform 1 0 39192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1610
timestamp 1624635492
transform 1 0 40296 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1624635492
transform -1 0 40388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_427
timestamp 1624635492
transform 1 0 40388 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_427
timestamp 1624635492
transform 1 0 40388 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1624635492
transform -1 0 40664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1624635492
transform -1 0 40940 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_430
timestamp 1624635492
transform 1 0 40664 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1624635492
transform -1 0 41308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_434
timestamp 1624635492
transform 1 0 41032 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_433
timestamp 1624635492
transform 1 0 40940 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_445
timestamp 1624635492
transform 1 0 42044 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_439
timestamp 1624635492
transform 1 0 41492 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_443
timestamp 1624635492
transform 1 0 41860 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_437
timestamp 1624635492
transform 1 0 41308 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input223_A
timestamp 1624635492
transform -1 0 42044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input221_A
timestamp 1624635492
transform -1 0 41492 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1624635492
transform -1 0 42412 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1624635492
transform -1 0 41860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1616
timestamp 1624635492
transform 1 0 42872 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input225_A
timestamp 1624635492
transform -1 0 42964 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_449
timestamp 1624635492
transform 1 0 42412 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_453
timestamp 1624635492
transform 1 0 42780 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input227_A
timestamp 1624635492
transform -1 0 43516 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input237_A
timestamp 1624635492
transform -1 0 43148 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input249_A
timestamp 1624635492
transform -1 0 43700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_455
timestamp 1624635492
transform 1 0 42964 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_457
timestamp 1624635492
transform 1 0 43148 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_461
timestamp 1624635492
transform 1 0 43516 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_469
timestamp 1624635492
transform 1 0 44252 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_463
timestamp 1624635492
transform 1 0 43700 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_470
timestamp 1624635492
transform 1 0 44344 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output507_A
timestamp 1624635492
transform 1 0 44620 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input255_A
timestamp 1624635492
transform -1 0 44252 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _314_
timestamp 1624635492
transform -1 0 44344 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input256_A
timestamp 1624635492
transform -1 0 44896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output520_A
timestamp 1624635492
transform -1 0 45356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_475
timestamp 1624635492
transform 1 0 44804 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1611
timestamp 1624635492
transform 1 0 45540 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output509_A
timestamp 1624635492
transform 1 0 45632 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output528_A
timestamp 1624635492
transform 1 0 45724 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_482
timestamp 1624635492
transform 1 0 45448 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_486
timestamp 1624635492
transform 1 0 45816 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_481
timestamp 1624635492
transform 1 0 45356 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_476
timestamp 1624635492
transform 1 0 44896 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_499
timestamp 1624635492
transform 1 0 47012 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_493
timestamp 1624635492
transform 1 0 46460 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_487
timestamp 1624635492
transform 1 0 45908 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_498
timestamp 1624635492
transform 1 0 46920 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_492
timestamp 1624635492
transform 1 0 46368 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output539_A
timestamp 1624635492
transform -1 0 47012 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output534_A
timestamp 1624635492
transform -1 0 46460 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output529_A
timestamp 1624635492
transform 1 0 46736 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output522_A
timestamp 1624635492
transform -1 0 46368 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_512
timestamp 1624635492
transform 1 0 48208 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_505
timestamp 1624635492
transform 1 0 47564 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_510
timestamp 1624635492
transform 1 0 48024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_504
timestamp 1624635492
transform 1 0 47472 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output543_A
timestamp 1624635492
transform 1 0 47380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output542_A
timestamp 1624635492
transform -1 0 48024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output535_A
timestamp 1624635492
transform -1 0 47472 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1617
timestamp 1624635492
transform 1 0 48116 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_524
timestamp 1624635492
transform 1 0 49312 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_522
timestamp 1624635492
transform 1 0 49128 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_536
timestamp 1624635492
transform 1 0 50416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_534
timestamp 1624635492
transform 1 0 50232 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_541
timestamp 1624635492
transform 1 0 50876 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1612
timestamp 1624635492
transform 1 0 50784 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_421
timestamp 1624635492
transform 1 0 39836 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_415
timestamp 1624635492
transform 1 0 39284 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1624635492
transform -1 0 39836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1624635492
transform -1 0 39284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_435
timestamp 1624635492
transform 1 0 41124 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1624635492
transform 1 0 40572 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_425
timestamp 1624635492
transform 1 0 40204 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input229_A
timestamp 1624635492
transform -1 0 41124 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input220_A
timestamp 1624635492
transform -1 0 40572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1621
timestamp 1624635492
transform 1 0 40296 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_447
timestamp 1624635492
transform 1 0 42228 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_441
timestamp 1624635492
transform 1 0 41676 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input246_A
timestamp 1624635492
transform -1 0 42228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input234_A
timestamp 1624635492
transform -1 0 41676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_459
timestamp 1624635492
transform 1 0 43332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_453
timestamp 1624635492
transform 1 0 42780 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output496_A
timestamp 1624635492
transform -1 0 43332 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input247_A
timestamp 1624635492
transform -1 0 42780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_471
timestamp 1624635492
transform 1 0 44436 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_465
timestamp 1624635492
transform 1 0 43884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output519_A
timestamp 1624635492
transform -1 0 44436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output500_A
timestamp 1624635492
transform -1 0 43884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_486
timestamp 1624635492
transform 1 0 45816 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1624635492
transform 1 0 44988 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output533_A
timestamp 1624635492
transform -1 0 45816 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output525_A
timestamp 1624635492
transform 1 0 44804 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1622
timestamp 1624635492
transform 1 0 45540 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_498
timestamp 1624635492
transform 1 0 46920 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_510
timestamp 1624635492
transform 1 0 48024 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _141_
timestamp 1624635492
transform 1 0 48116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_514
timestamp 1624635492
transform 1 0 48392 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_538
timestamp 1624635492
transform 1 0 50600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_526
timestamp 1624635492
transform 1 0 49496 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_541
timestamp 1624635492
transform 1 0 50876 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1623
timestamp 1624635492
transform 1 0 50784 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_421
timestamp 1624635492
transform 1 0 39836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_415
timestamp 1624635492
transform 1 0 39284 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input219_A
timestamp 1624635492
transform -1 0 39836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input216_A
timestamp 1624635492
transform -1 0 39284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_435
timestamp 1624635492
transform 1 0 41124 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_432
timestamp 1624635492
transform 1 0 40848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_428
timestamp 1624635492
transform 1 0 40480 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_425
timestamp 1624635492
transform 1 0 40204 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input235_A
timestamp 1624635492
transform -1 0 41124 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input232_A
timestamp 1624635492
transform -1 0 40480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_445
timestamp 1624635492
transform 1 0 42044 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output492_A
timestamp 1624635492
transform 1 0 41860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_457
timestamp 1624635492
transform 1 0 43148 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_453
timestamp 1624635492
transform 1 0 42780 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output512_A
timestamp 1624635492
transform -1 0 43700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output504_A
timestamp 1624635492
transform 1 0 42964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1627
timestamp 1624635492
transform 1 0 42872 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_469
timestamp 1624635492
transform 1 0 44252 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_463
timestamp 1624635492
transform 1 0 43700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output531_A
timestamp 1624635492
transform -1 0 44804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output523_A
timestamp 1624635492
transform 1 0 44068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_475
timestamp 1624635492
transform 1 0 44804 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_499
timestamp 1624635492
transform 1 0 47012 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_487
timestamp 1624635492
transform 1 0 45908 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_512
timestamp 1624635492
transform 1 0 48208 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1628
timestamp 1624635492
transform 1 0 48116 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_524
timestamp 1624635492
transform 1 0 49312 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_536
timestamp 1624635492
transform 1 0 50416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1624635492
transform 1 0 39836 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_415
timestamp 1624635492
transform 1 0 39284 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input233_A
timestamp 1624635492
transform -1 0 39836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input226_A
timestamp 1624635492
transform -1 0 39284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_435
timestamp 1624635492
transform 1 0 41124 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_429
timestamp 1624635492
transform 1 0 40572 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_425
timestamp 1624635492
transform 1 0 40204 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output490_A
timestamp 1624635492
transform -1 0 41124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input244_A
timestamp 1624635492
transform -1 0 40572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1632
timestamp 1624635492
transform 1 0 40296 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_447
timestamp 1624635492
transform 1 0 42228 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_441
timestamp 1624635492
transform 1 0 41676 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output503_A
timestamp 1624635492
transform -1 0 42228 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output497_A
timestamp 1624635492
transform -1 0 41676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_459
timestamp 1624635492
transform 1 0 43332 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_453
timestamp 1624635492
transform 1 0 42780 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output521_A
timestamp 1624635492
transform -1 0 43332 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output508_A
timestamp 1624635492
transform -1 0 42780 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_471
timestamp 1624635492
transform 1 0 44436 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_484
timestamp 1624635492
transform 1 0 45632 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1633
timestamp 1624635492
transform 1 0 45540 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_496
timestamp 1624635492
transform 1 0 46736 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_511
timestamp 1624635492
transform 1 0 48116 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _245_
timestamp 1624635492
transform 1 0 47840 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_523
timestamp 1624635492
transform 1 0 49220 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_535
timestamp 1624635492
transform 1 0 50324 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_541
timestamp 1624635492
transform 1 0 50876 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_539
timestamp 1624635492
transform 1 0 50692 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1634
timestamp 1624635492
transform 1 0 50784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_420
timestamp 1624635492
transform 1 0 39744 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_414
timestamp 1624635492
transform 1 0 39192 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output487_A
timestamp 1624635492
transform -1 0 39744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1624635492
transform 1 0 39008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_434
timestamp 1624635492
transform 1 0 41032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_426
timestamp 1624635492
transform 1 0 40296 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output499_A
timestamp 1624635492
transform 1 0 40848 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output488_A
timestamp 1624635492
transform -1 0 40296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_446
timestamp 1624635492
transform 1 0 42136 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_440
timestamp 1624635492
transform 1 0 41584 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output514_A
timestamp 1624635492
transform 1 0 41952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output506_A
timestamp 1624635492
transform 1 0 41400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_455
timestamp 1624635492
transform 1 0 42964 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1638
timestamp 1624635492
transform 1 0 42872 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_467
timestamp 1624635492
transform 1 0 44068 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_479
timestamp 1624635492
transform 1 0 45172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_491
timestamp 1624635492
transform 1 0 46276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_512
timestamp 1624635492
transform 1 0 48208 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_503
timestamp 1624635492
transform 1 0 47380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1639
timestamp 1624635492
transform 1 0 48116 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_524
timestamp 1624635492
transform 1 0 49312 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_536
timestamp 1624635492
transform 1 0 50416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_422
timestamp 1624635492
transform 1 0 39928 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1624635492
transform 1 0 39376 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_410
timestamp 1624635492
transform 1 0 38824 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output501_A
timestamp 1624635492
transform -1 0 39928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output495_A
timestamp 1624635492
transform -1 0 39376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_435
timestamp 1624635492
transform 1 0 41124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_429
timestamp 1624635492
transform 1 0 40572 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output515_A
timestamp 1624635492
transform -1 0 41124 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output502_A
timestamp 1624635492
transform 1 0 40388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1643
timestamp 1624635492
transform 1 0 40296 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_441
timestamp 1624635492
transform 1 0 41676 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output524_A
timestamp 1624635492
transform -1 0 41676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_453
timestamp 1624635492
transform 1 0 42780 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_465
timestamp 1624635492
transform 1 0 43884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_484
timestamp 1624635492
transform 1 0 45632 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_477
timestamp 1624635492
transform 1 0 44988 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1644
timestamp 1624635492
transform 1 0 45540 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_496
timestamp 1624635492
transform 1 0 46736 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_508
timestamp 1624635492
transform 1 0 47840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_520
timestamp 1624635492
transform 1 0 48944 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_532
timestamp 1624635492
transform 1 0 50048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_541
timestamp 1624635492
transform 1 0 50876 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1645
timestamp 1624635492
transform 1 0 50784 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_416
timestamp 1624635492
transform 1 0 39376 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_421
timestamp 1624635492
transform 1 0 39836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_415
timestamp 1624635492
transform 1 0 39284 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output510_A
timestamp 1624635492
transform 1 0 39652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output498_A
timestamp 1624635492
transform -1 0 39284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_427
timestamp 1624635492
transform 1 0 40388 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_424
timestamp 1624635492
transform 1 0 40112 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_433
timestamp 1624635492
transform 1 0 40940 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1654
timestamp 1624635492
transform 1 0 40296 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_439
timestamp 1624635492
transform 1 0 41492 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_445
timestamp 1624635492
transform 1 0 42044 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_451
timestamp 1624635492
transform 1 0 42596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_455
timestamp 1624635492
transform 1 0 42964 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_453
timestamp 1624635492
transform 1 0 42780 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1649
timestamp 1624635492
transform 1 0 42872 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_463
timestamp 1624635492
transform 1 0 43700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_467
timestamp 1624635492
transform 1 0 44068 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_484
timestamp 1624635492
transform 1 0 45632 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_475
timestamp 1624635492
transform 1 0 44804 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_479
timestamp 1624635492
transform 1 0 45172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1655
timestamp 1624635492
transform 1 0 45540 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_496
timestamp 1624635492
transform 1 0 46736 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_491
timestamp 1624635492
transform 1 0 46276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_508
timestamp 1624635492
transform 1 0 47840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_512
timestamp 1624635492
transform 1 0 48208 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_503
timestamp 1624635492
transform 1 0 47380 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1650
timestamp 1624635492
transform 1 0 48116 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_520
timestamp 1624635492
transform 1 0 48944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_524
timestamp 1624635492
transform 1 0 49312 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_532
timestamp 1624635492
transform 1 0 50048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_536
timestamp 1624635492
transform 1 0 50416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_541
timestamp 1624635492
transform 1 0 50876 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1656
timestamp 1624635492
transform 1 0 50784 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_412
timestamp 1624635492
transform 1 0 39008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_424
timestamp 1624635492
transform 1 0 40112 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_448
timestamp 1624635492
transform 1 0 42320 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_436
timestamp 1624635492
transform 1 0 41216 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_455
timestamp 1624635492
transform 1 0 42964 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1660
timestamp 1624635492
transform 1 0 42872 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_467
timestamp 1624635492
transform 1 0 44068 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_479
timestamp 1624635492
transform 1 0 45172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_491
timestamp 1624635492
transform 1 0 46276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_512
timestamp 1624635492
transform 1 0 48208 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_503
timestamp 1624635492
transform 1 0 47380 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1661
timestamp 1624635492
transform 1 0 48116 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_524
timestamp 1624635492
transform 1 0 49312 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_536
timestamp 1624635492
transform 1 0 50416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_412
timestamp 1624635492
transform 1 0 39008 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_427
timestamp 1624635492
transform 1 0 40388 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_424
timestamp 1624635492
transform 1 0 40112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1665
timestamp 1624635492
transform 1 0 40296 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_439
timestamp 1624635492
transform 1 0 41492 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_451
timestamp 1624635492
transform 1 0 42596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_463
timestamp 1624635492
transform 1 0 43700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_484
timestamp 1624635492
transform 1 0 45632 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_475
timestamp 1624635492
transform 1 0 44804 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1666
timestamp 1624635492
transform 1 0 45540 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_496
timestamp 1624635492
transform 1 0 46736 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_508
timestamp 1624635492
transform 1 0 47840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_520
timestamp 1624635492
transform 1 0 48944 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_532
timestamp 1624635492
transform 1 0 50048 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_541
timestamp 1624635492
transform 1 0 50876 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1667
timestamp 1624635492
transform 1 0 50784 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_412
timestamp 1624635492
transform 1 0 39008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_424
timestamp 1624635492
transform 1 0 40112 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_448
timestamp 1624635492
transform 1 0 42320 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_436
timestamp 1624635492
transform 1 0 41216 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_455
timestamp 1624635492
transform 1 0 42964 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1671
timestamp 1624635492
transform 1 0 42872 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_467
timestamp 1624635492
transform 1 0 44068 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_479
timestamp 1624635492
transform 1 0 45172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_491
timestamp 1624635492
transform 1 0 46276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_512
timestamp 1624635492
transform 1 0 48208 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_503
timestamp 1624635492
transform 1 0 47380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1672
timestamp 1624635492
transform 1 0 48116 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_524
timestamp 1624635492
transform 1 0 49312 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_536
timestamp 1624635492
transform 1 0 50416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_412
timestamp 1624635492
transform 1 0 39008 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_427
timestamp 1624635492
transform 1 0 40388 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_424
timestamp 1624635492
transform 1 0 40112 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1676
timestamp 1624635492
transform 1 0 40296 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_439
timestamp 1624635492
transform 1 0 41492 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_451
timestamp 1624635492
transform 1 0 42596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_463
timestamp 1624635492
transform 1 0 43700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_484
timestamp 1624635492
transform 1 0 45632 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_475
timestamp 1624635492
transform 1 0 44804 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1677
timestamp 1624635492
transform 1 0 45540 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_496
timestamp 1624635492
transform 1 0 46736 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_508
timestamp 1624635492
transform 1 0 47840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_520
timestamp 1624635492
transform 1 0 48944 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_532
timestamp 1624635492
transform 1 0 50048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_541
timestamp 1624635492
transform 1 0 50876 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1678
timestamp 1624635492
transform 1 0 50784 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_559
timestamp 1624635492
transform 1 0 52532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_551
timestamp 1624635492
transform 1 0 51796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output547
timestamp 1624635492
transform -1 0 52532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output544
timestamp 1624635492
transform -1 0 51796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_567
timestamp 1624635492
transform 1 0 53268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output550
timestamp 1624635492
transform -1 0 53268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1533
timestamp 1624635492
transform 1 0 53636 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_580
timestamp 1624635492
transform 1 0 54464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_572
timestamp 1624635492
transform 1 0 53728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output555
timestamp 1624635492
transform -1 0 55200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output553
timestamp 1624635492
transform -1 0 54464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_596
timestamp 1624635492
transform 1 0 55936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_588
timestamp 1624635492
transform 1 0 55200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output557
timestamp 1624635492
transform -1 0 55936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_610
timestamp 1624635492
transform 1 0 57224 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_605
timestamp 1624635492
transform 1 0 56764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_601
timestamp 1624635492
transform 1 0 56396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output449
timestamp 1624635492
transform 1 0 56856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1534
timestamp 1624635492
transform 1 0 56304 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_618
timestamp 1624635492
transform 1 0 57960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output445
timestamp 1624635492
transform -1 0 57960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1624635492
transform -1 0 58604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_630
timestamp 1624635492
transform 1 0 59064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_625
timestamp 1624635492
transform 1 0 58604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output446
timestamp 1624635492
transform -1 0 59800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1535
timestamp 1624635492
transform 1 0 58972 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_646
timestamp 1624635492
transform 1 0 60536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_638
timestamp 1624635492
transform 1 0 59800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output447
timestamp 1624635492
transform -1 0 60536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_659
timestamp 1624635492
transform 1 0 61732 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_654
timestamp 1624635492
transform 1 0 61272 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output448
timestamp 1624635492
transform -1 0 61272 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1536
timestamp 1624635492
transform 1 0 61640 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_667
timestamp 1624635492
transform 1 0 62468 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output451
timestamp 1624635492
transform -1 0 63204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output450
timestamp 1624635492
transform -1 0 62468 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_675
timestamp 1624635492
transform 1 0 63204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output452
timestamp 1624635492
transform -1 0 63940 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_555
timestamp 1624635492
transform 1 0 52164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_548
timestamp 1624635492
transform 1 0 51520 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_552
timestamp 1624635492
transform 1 0 51888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output558
timestamp 1624635492
transform -1 0 52900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output556
timestamp 1624635492
transform -1 0 52624 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output554
timestamp 1624635492
transform -1 0 51888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1624635492
transform 1 0 51888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_567
timestamp 1624635492
transform 1 0 53268 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_563
timestamp 1624635492
transform 1 0 52900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_569
timestamp 1624635492
transform 1 0 53452 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_560
timestamp 1624635492
transform 1 0 52624 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output561
timestamp 1624635492
transform -1 0 53728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1541
timestamp 1624635492
transform 1 0 53360 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_582
timestamp 1624635492
transform 1 0 54648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_572
timestamp 1624635492
transform 1 0 53728 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_577
timestamp 1624635492
transform 1 0 54188 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output563
timestamp 1624635492
transform -1 0 54648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output562
timestamp 1624635492
transform -1 0 54924 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output559
timestamp 1624635492
transform -1 0 54188 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_591
timestamp 1624635492
transform 1 0 55476 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_586
timestamp 1624635492
transform 1 0 55016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_593
timestamp 1624635492
transform 1 0 55660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1624635492
transform 1 0 54924 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output566
timestamp 1624635492
transform -1 0 56396 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output565
timestamp 1624635492
transform -1 0 55476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output564
timestamp 1624635492
transform -1 0 55660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1547
timestamp 1624635492
transform 1 0 56028 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1624635492
transform 1 0 56856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_598
timestamp 1624635492
transform 1 0 56120 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_609
timestamp 1624635492
transform 1 0 57132 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_601
timestamp 1624635492
transform 1 0 56396 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output570
timestamp 1624635492
transform -1 0 57592 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output568
timestamp 1624635492
transform -1 0 56856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output567
timestamp 1624635492
transform -1 0 57132 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_621
timestamp 1624635492
transform 1 0 58236 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_614
timestamp 1624635492
transform 1 0 57592 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_617
timestamp 1624635492
transform 1 0 57868 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output569
timestamp 1624635492
transform -1 0 57868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform -1 0 58236 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_630
timestamp 1624635492
transform 1 0 59064 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_633
timestamp 1624635492
transform 1 0 59340 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_626
timestamp 1624635492
transform 1 0 58696 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1624635492
transform 1 0 59432 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1624635492
transform -1 0 59064 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1624635492
transform -1 0 59340 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1542
timestamp 1624635492
transform 1 0 58604 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_644
timestamp 1624635492
transform 1 0 60352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_637
timestamp 1624635492
transform 1 0 59708 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_647
timestamp 1624635492
transform 1 0 60628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_640
timestamp 1624635492
transform 1 0 59984 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 60904 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1624635492
transform -1 0 60352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1624635492
transform 1 0 60352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1624635492
transform -1 0 59984 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_655
timestamp 1624635492
transform 1 0 61364 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_650
timestamp 1624635492
transform 1 0 60904 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_661
timestamp 1624635492
transform 1 0 61916 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_655
timestamp 1624635492
transform 1 0 61364 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 61916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output453
timestamp 1624635492
transform -1 0 61364 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1624635492
transform -1 0 62008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1548
timestamp 1624635492
transform 1 0 61272 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_669
timestamp 1624635492
transform 1 0 62652 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_662
timestamp 1624635492
transform 1 0 62008 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_673
timestamp 1624635492
transform 1 0 63020 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_669
timestamp 1624635492
transform 1 0 62652 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output459
timestamp 1624635492
transform 1 0 63112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output457
timestamp 1624635492
transform -1 0 62652 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1624635492
transform 1 0 63020 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1624635492
transform 1 0 62376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_676
timestamp 1624635492
transform 1 0 63296 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_678
timestamp 1624635492
transform 1 0 63480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1543
timestamp 1624635492
transform 1 0 63848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_554
timestamp 1624635492
transform 1 0 52072 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_547
timestamp 1624635492
transform 1 0 51428 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1624635492
transform 1 0 52440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1624635492
transform -1 0 52072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_569
timestamp 1624635492
transform 1 0 53452 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_567
timestamp 1624635492
transform 1 0 53268 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_561
timestamp 1624635492
transform 1 0 52716 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1552
timestamp 1624635492
transform 1 0 53360 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_583
timestamp 1624635492
transform 1 0 54740 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_576
timestamp 1624635492
transform 1 0 54096 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input156
timestamp 1624635492
transform 1 0 54464 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input153
timestamp 1624635492
transform 1 0 53820 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_597
timestamp 1624635492
transform 1 0 56028 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_590
timestamp 1624635492
transform 1 0 55384 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1624635492
transform 1 0 55752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1624635492
transform 1 0 55108 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_604
timestamp 1624635492
transform 1 0 56672 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1624635492
transform -1 0 57316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input162
timestamp 1624635492
transform -1 0 56672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_620
timestamp 1624635492
transform 1 0 58144 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_611
timestamp 1624635492
transform 1 0 57316 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _295_
timestamp 1624635492
transform 1 0 57868 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_633
timestamp 1624635492
transform 1 0 59340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_626
timestamp 1624635492
transform 1 0 58696 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_624
timestamp 1624635492
transform 1 0 58512 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input169
timestamp 1624635492
transform 1 0 59064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1553
timestamp 1624635492
transform 1 0 58604 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_648
timestamp 1624635492
transform 1 0 60720 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_644
timestamp 1624635492
transform 1 0 60352 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_640
timestamp 1624635492
transform 1 0 59984 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1624635492
transform 1 0 59708 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1624635492
transform -1 0 60720 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_658
timestamp 1624635492
transform 1 0 61640 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_654
timestamp 1624635492
transform 1 0 61272 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1624635492
transform -1 0 61640 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_671
timestamp 1624635492
transform 1 0 62836 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_664
timestamp 1624635492
transform 1 0 62192 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 62192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1624635492
transform -1 0 62836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_678
timestamp 1624635492
transform 1 0 63480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1624635492
transform -1 0 63480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1554
timestamp 1624635492
transform 1 0 63848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_555
timestamp 1624635492
transform 1 0 52164 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_548
timestamp 1624635492
transform 1 0 51520 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input275
timestamp 1624635492
transform -1 0 52164 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_571
timestamp 1624635492
transform 1 0 53636 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_564
timestamp 1624635492
transform 1 0 52992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input154
timestamp 1624635492
transform 1 0 53360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _243_
timestamp 1624635492
transform -1 0 52992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_578
timestamp 1624635492
transform 1 0 54280 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1624635492
transform 1 0 54648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input157
timestamp 1624635492
transform 1 0 54004 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_593
timestamp 1624635492
transform 1 0 55660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_589
timestamp 1624635492
transform 1 0 55292 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_585
timestamp 1624635492
transform 1 0 54924 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input161
timestamp 1624635492
transform -1 0 55660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1558
timestamp 1624635492
transform 1 0 56028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_607
timestamp 1624635492
transform 1 0 56948 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_600
timestamp 1624635492
transform 1 0 56304 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input151_A
timestamp 1624635492
transform -1 0 56304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input164
timestamp 1624635492
transform -1 0 56948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1624635492
transform 1 0 58236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_614
timestamp 1624635492
transform 1 0 57592 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input292
timestamp 1624635492
transform 1 0 57960 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input165
timestamp 1624635492
transform -1 0 57592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_634
timestamp 1624635492
transform 1 0 59432 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_628
timestamp 1624635492
transform 1 0 58880 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input172
timestamp 1624635492
transform -1 0 59800 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input170
timestamp 1624635492
transform -1 0 58880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_645
timestamp 1624635492
transform 1 0 60444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_638
timestamp 1624635492
transform 1 0 59800 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _137_
timestamp 1624635492
transform -1 0 60444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_655
timestamp 1624635492
transform 1 0 61364 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_653
timestamp 1624635492
transform 1 0 61180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1559
timestamp 1624635492
transform 1 0 61272 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _216_
timestamp 1624635492
transform -1 0 62008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_669
timestamp 1624635492
transform 1 0 62652 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_662
timestamp 1624635492
transform 1 0 62008 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input180
timestamp 1624635492
transform -1 0 63296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input177
timestamp 1624635492
transform 1 0 62376 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_676
timestamp 1624635492
transform 1 0 63296 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1624635492
transform -1 0 64124 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_558
timestamp 1624635492
transform 1 0 52440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_551
timestamp 1624635492
transform 1 0 51796 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input277
timestamp 1624635492
transform 1 0 52164 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_569
timestamp 1624635492
transform 1 0 53452 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_564
timestamp 1624635492
transform 1 0 52992 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1624635492
transform -1 0 52992 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1563
timestamp 1624635492
transform 1 0 53360 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_583
timestamp 1624635492
transform 1 0 54740 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_576
timestamp 1624635492
transform 1 0 54096 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input284
timestamp 1624635492
transform 1 0 54464 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input280
timestamp 1624635492
transform -1 0 54096 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_597
timestamp 1624635492
transform 1 0 56028 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_590
timestamp 1624635492
transform 1 0 55384 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input288
timestamp 1624635492
transform -1 0 56028 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input286
timestamp 1624635492
transform -1 0 55384 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_604
timestamp 1624635492
transform 1 0 56672 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input291
timestamp 1624635492
transform -1 0 57316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input289
timestamp 1624635492
transform 1 0 56396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_618
timestamp 1624635492
transform 1 0 57960 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_611
timestamp 1624635492
transform 1 0 57316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input293
timestamp 1624635492
transform -1 0 57960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_634
timestamp 1624635492
transform 1 0 59432 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_628
timestamp 1624635492
transform 1 0 58880 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_624
timestamp 1624635492
transform 1 0 58512 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 59432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 58880 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1564
timestamp 1624635492
transform 1 0 58604 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_642
timestamp 1624635492
transform 1 0 60168 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_638
timestamp 1624635492
transform 1 0 59800 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input174
timestamp 1624635492
transform 1 0 60536 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input173
timestamp 1624635492
transform -1 0 60168 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_656
timestamp 1624635492
transform 1 0 61456 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_649
timestamp 1624635492
transform 1 0 60812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input176
timestamp 1624635492
transform 1 0 61824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input175
timestamp 1624635492
transform -1 0 61456 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_670
timestamp 1624635492
transform 1 0 62744 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_663
timestamp 1624635492
transform 1 0 62100 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input181
timestamp 1624635492
transform 1 0 63112 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input179
timestamp 1624635492
transform -1 0 62744 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_681
timestamp 1624635492
transform 1 0 63756 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_677
timestamp 1624635492
transform 1 0 63388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1565
timestamp 1624635492
transform 1 0 63848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_555
timestamp 1624635492
transform 1 0 52164 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_548
timestamp 1624635492
transform 1 0 51520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input279
timestamp 1624635492
transform -1 0 52808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input278
timestamp 1624635492
transform -1 0 52164 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_569
timestamp 1624635492
transform 1 0 53452 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_562
timestamp 1624635492
transform 1 0 52808 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input281
timestamp 1624635492
transform 1 0 53176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_583
timestamp 1624635492
transform 1 0 54740 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_576
timestamp 1624635492
transform 1 0 54096 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input285
timestamp 1624635492
transform -1 0 54740 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input282
timestamp 1624635492
transform -1 0 54096 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_596
timestamp 1624635492
transform 1 0 55936 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_590
timestamp 1624635492
transform 1 0 55384 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input287
timestamp 1624635492
transform -1 0 55384 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1569
timestamp 1624635492
transform 1 0 56028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_605
timestamp 1624635492
transform 1 0 56764 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_598
timestamp 1624635492
transform 1 0 56120 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input162_A
timestamp 1624635492
transform -1 0 57316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input290
timestamp 1624635492
transform -1 0 56764 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_617
timestamp 1624635492
transform 1 0 57868 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_611
timestamp 1624635492
transform 1 0 57316 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input163_A
timestamp 1624635492
transform -1 0 57868 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_634
timestamp 1624635492
transform 1 0 59432 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_628
timestamp 1624635492
transform 1 0 58880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_625
timestamp 1624635492
transform 1 0 58604 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input169_A
timestamp 1624635492
transform -1 0 58880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input168_A
timestamp 1624635492
transform -1 0 59432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_644
timestamp 1624635492
transform 1 0 60352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 60904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 60352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_657
timestamp 1624635492
transform 1 0 61548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_650
timestamp 1624635492
transform 1 0 60904 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 62100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 61548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1570
timestamp 1624635492
transform 1 0 61272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_672
timestamp 1624635492
transform 1 0 62928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_663
timestamp 1624635492
transform 1 0 62100 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input295
timestamp 1624635492
transform -1 0 62928 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_679
timestamp 1624635492
transform 1 0 63572 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input182
timestamp 1624635492
transform -1 0 63572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_555
timestamp 1624635492
transform 1 0 52164 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_549
timestamp 1624635492
transform 1 0 51612 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_554
timestamp 1624635492
transform 1 0 52072 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_550
timestamp 1624635492
transform 1 0 51704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input152_A
timestamp 1624635492
transform -1 0 52716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input150_A
timestamp 1624635492
transform -1 0 52164 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input149_A
timestamp 1624635492
transform -1 0 52624 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input148_A
timestamp 1624635492
transform -1 0 51612 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _263_
timestamp 1624635492
transform 1 0 51796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_568
timestamp 1624635492
transform 1 0 53360 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_565
timestamp 1624635492
transform 1 0 53084 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_561
timestamp 1624635492
transform 1 0 52716 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_569
timestamp 1624635492
transform 1 0 53452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_560
timestamp 1624635492
transform 1 0 52624 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input154_A
timestamp 1624635492
transform -1 0 53360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input153_A
timestamp 1624635492
transform -1 0 53820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1574
timestamp 1624635492
transform 1 0 53360 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input157_A
timestamp 1624635492
transform -1 0 54004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_573
timestamp 1624635492
transform 1 0 53820 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_572
timestamp 1624635492
transform 1 0 53728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_575
timestamp 1624635492
transform 1 0 54004 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input156_A
timestamp 1624635492
transform -1 0 54464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input159_A
timestamp 1624635492
transform -1 0 54648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_577
timestamp 1624635492
transform 1 0 54188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_580
timestamp 1624635492
transform 1 0 54464 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_579
timestamp 1624635492
transform 1 0 54372 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_584
timestamp 1624635492
transform 1 0 54832 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_582
timestamp 1624635492
transform 1 0 54648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_596
timestamp 1624635492
transform 1 0 55936 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_588
timestamp 1624635492
transform 1 0 55200 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_594
timestamp 1624635492
transform 1 0 55752 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_591
timestamp 1624635492
transform 1 0 55476 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_587
timestamp 1624635492
transform 1 0 55108 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input282_A
timestamp 1624635492
transform -1 0 55200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input160_A
timestamp 1624635492
transform -1 0 55752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input158_A
timestamp 1624635492
transform -1 0 55108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1580
timestamp 1624635492
transform 1 0 56028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input161_A
timestamp 1624635492
transform -1 0 56304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input286_A
timestamp 1624635492
transform -1 0 56304 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input288_A
timestamp 1624635492
transform -1 0 56856 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_600
timestamp 1624635492
transform 1 0 56304 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input164_A
timestamp 1624635492
transform -1 0 57132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input291_A
timestamp 1624635492
transform -1 0 57408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_606
timestamp 1624635492
transform 1 0 56856 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_609
timestamp 1624635492
transform 1 0 57132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_606
timestamp 1624635492
transform 1 0 56856 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_600
timestamp 1624635492
transform 1 0 56304 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_618
timestamp 1624635492
transform 1 0 57960 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_612
timestamp 1624635492
transform 1 0 57408 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1624635492
transform 1 0 58236 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_615
timestamp 1624635492
transform 1 0 57684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input293_A
timestamp 1624635492
transform -1 0 58512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input292_A
timestamp 1624635492
transform -1 0 57960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input290_A
timestamp 1624635492
transform -1 0 58236 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input165_A
timestamp 1624635492
transform -1 0 57684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_634
timestamp 1624635492
transform 1 0 59432 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_624
timestamp 1624635492
transform 1 0 58512 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_634
timestamp 1624635492
transform 1 0 59432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_630
timestamp 1624635492
transform 1 0 59064 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_626
timestamp 1624635492
transform 1 0 58696 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output446_A
timestamp 1624635492
transform 1 0 59248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input171_A
timestamp 1624635492
transform -1 0 59708 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input170_A
timestamp 1624635492
transform -1 0 59064 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1575
timestamp 1624635492
transform 1 0 58604 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_646
timestamp 1624635492
transform 1 0 60536 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_640
timestamp 1624635492
transform 1 0 59984 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_643
timestamp 1624635492
transform 1 0 60260 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_637
timestamp 1624635492
transform 1 0 59708 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output447_A
timestamp 1624635492
transform -1 0 59984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input174_A
timestamp 1624635492
transform -1 0 60536 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input173_A
timestamp 1624635492
transform -1 0 60812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input172_A
timestamp 1624635492
transform -1 0 60260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_657
timestamp 1624635492
transform 1 0 61548 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_660
timestamp 1624635492
transform 1 0 61824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_657
timestamp 1624635492
transform 1 0 61548 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_649
timestamp 1624635492
transform 1 0 60812 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input176_A
timestamp 1624635492
transform -1 0 62100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input175_A
timestamp 1624635492
transform -1 0 61548 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 61824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1581
timestamp 1624635492
transform 1 0 61272 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_673
timestamp 1624635492
transform 1 0 63020 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_663
timestamp 1624635492
transform 1 0 62100 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_673
timestamp 1624635492
transform 1 0 63020 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_670
timestamp 1624635492
transform 1 0 62744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_666
timestamp 1624635492
transform 1 0 62376 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 63020 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 63020 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 62376 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_679
timestamp 1624635492
transform 1 0 63572 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_681
timestamp 1624635492
transform 1 0 63756 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 63572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1576
timestamp 1624635492
transform 1 0 63848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_556
timestamp 1624635492
transform 1 0 52256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_550
timestamp 1624635492
transform 1 0 51704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input275_A
timestamp 1624635492
transform -1 0 52256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input271_A
timestamp 1624635492
transform -1 0 51704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_571
timestamp 1624635492
transform 1 0 53636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_562
timestamp 1624635492
transform 1 0 52808 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input279_A
timestamp 1624635492
transform -1 0 53636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input276_A
timestamp 1624635492
transform -1 0 52808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1585
timestamp 1624635492
transform 1 0 53360 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_583
timestamp 1624635492
transform 1 0 54740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_577
timestamp 1624635492
transform 1 0 54188 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input284_A
timestamp 1624635492
transform -1 0 54740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input280_A
timestamp 1624635492
transform -1 0 54188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_595
timestamp 1624635492
transform 1 0 55844 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_589
timestamp 1624635492
transform 1 0 55292 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input287_A
timestamp 1624635492
transform -1 0 55844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input285_A
timestamp 1624635492
transform -1 0 55292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_607
timestamp 1624635492
transform 1 0 56948 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_601
timestamp 1624635492
transform 1 0 56396 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output449_A
timestamp 1624635492
transform 1 0 56764 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input289_A
timestamp 1624635492
transform -1 0 56396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_620
timestamp 1624635492
transform 1 0 58144 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_617
timestamp 1624635492
transform 1 0 57868 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_613
timestamp 1624635492
transform 1 0 57500 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output568_A
timestamp 1624635492
transform -1 0 57500 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output445_A
timestamp 1624635492
transform 1 0 57960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_634
timestamp 1624635492
transform 1 0 59432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_626
timestamp 1624635492
transform 1 0 58696 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_624
timestamp 1624635492
transform 1 0 58512 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output474_A
timestamp 1624635492
transform -1 0 59800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1586
timestamp 1624635492
transform 1 0 58604 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_644
timestamp 1624635492
transform 1 0 60352 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_638
timestamp 1624635492
transform 1 0 59800 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output453_A
timestamp 1624635492
transform 1 0 60168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output448_A
timestamp 1624635492
transform 1 0 60720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_660
timestamp 1624635492
transform 1 0 61824 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_650
timestamp 1624635492
transform 1 0 60904 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output450_A
timestamp 1624635492
transform 1 0 61640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_672
timestamp 1624635492
transform 1 0 62928 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_666
timestamp 1624635492
transform 1 0 62376 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input179_A
timestamp 1624635492
transform -1 0 62928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input177_A
timestamp 1624635492
transform -1 0 62376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_678
timestamp 1624635492
transform 1 0 63480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input180_A
timestamp 1624635492
transform -1 0 63480 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1587
timestamp 1624635492
transform 1 0 63848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_555
timestamp 1624635492
transform 1 0 52164 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_549
timestamp 1624635492
transform 1 0 51612 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input278_A
timestamp 1624635492
transform -1 0 52716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input277_A
timestamp 1624635492
transform -1 0 52164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input274_A
timestamp 1624635492
transform -1 0 51612 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_567
timestamp 1624635492
transform 1 0 53268 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_561
timestamp 1624635492
transform 1 0 52716 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output550_A
timestamp 1624635492
transform 1 0 53636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input281_A
timestamp 1624635492
transform -1 0 53268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_582
timestamp 1624635492
transform 1 0 54648 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_579
timestamp 1624635492
transform 1 0 54372 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_573
timestamp 1624635492
transform 1 0 53820 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output553_A
timestamp 1624635492
transform 1 0 54464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_596
timestamp 1624635492
transform 1 0 55936 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_590
timestamp 1624635492
transform 1 0 55384 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output555_A
timestamp 1624635492
transform 1 0 55200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1591
timestamp 1624635492
transform 1 0 56028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_610
timestamp 1624635492
transform 1 0 57224 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_606
timestamp 1624635492
transform 1 0 56856 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_600
timestamp 1624635492
transform 1 0 56304 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output566_A
timestamp 1624635492
transform -1 0 56856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output557_A
timestamp 1624635492
transform -1 0 56304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_619
timestamp 1624635492
transform 1 0 58052 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_613
timestamp 1624635492
transform 1 0 57500 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output570_A
timestamp 1624635492
transform -1 0 58052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output569_A
timestamp 1624635492
transform 1 0 57316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_631
timestamp 1624635492
transform 1 0 59156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_647
timestamp 1624635492
transform 1 0 60628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_643
timestamp 1624635492
transform 1 0 60260 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output473_A
timestamp 1624635492
transform 1 0 60720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_659
timestamp 1624635492
transform 1 0 61732 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_655
timestamp 1624635492
transform 1 0 61364 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_650
timestamp 1624635492
transform 1 0 60904 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output451_A
timestamp 1624635492
transform 1 0 61824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1592
timestamp 1624635492
transform 1 0 61272 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_674
timestamp 1624635492
transform 1 0 63112 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_668
timestamp 1624635492
transform 1 0 62560 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_662
timestamp 1624635492
transform 1 0 62008 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output417_A
timestamp 1624635492
transform 1 0 62376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input181_A
timestamp 1624635492
transform -1 0 63112 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_681
timestamp 1624635492
transform 1 0 63756 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_678
timestamp 1624635492
transform 1 0 63480 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input195_A
timestamp 1624635492
transform -1 0 63756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_555
timestamp 1624635492
transform 1 0 52164 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_549
timestamp 1624635492
transform 1 0 51612 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output554_A
timestamp 1624635492
transform -1 0 52716 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B1
timestamp 1624635492
transform -1 0 52164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_571
timestamp 1624635492
transform 1 0 53636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_567
timestamp 1624635492
transform 1 0 53268 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_561
timestamp 1624635492
transform 1 0 52716 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output558_A
timestamp 1624635492
transform -1 0 53636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1596
timestamp 1624635492
transform 1 0 53360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_583
timestamp 1624635492
transform 1 0 54740 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_577
timestamp 1624635492
transform 1 0 54188 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output562_A
timestamp 1624635492
transform 1 0 54556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output559_A
timestamp 1624635492
transform -1 0 54188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_595
timestamp 1624635492
transform 1 0 55844 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_589
timestamp 1624635492
transform 1 0 55292 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output565_A
timestamp 1624635492
transform -1 0 55844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output564_A
timestamp 1624635492
transform 1 0 55108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_607
timestamp 1624635492
transform 1 0 56948 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_619
timestamp 1624635492
transform 1 0 58052 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_626
timestamp 1624635492
transform 1 0 58696 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1597
timestamp 1624635492
transform 1 0 58604 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_638
timestamp 1624635492
transform 1 0 59800 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_658
timestamp 1624635492
transform 1 0 61640 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_654
timestamp 1624635492
transform 1 0 61272 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_650
timestamp 1624635492
transform 1 0 60904 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _200_
timestamp 1624635492
transform -1 0 61640 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_674
timestamp 1624635492
transform 1 0 63112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1624635492
transform 1 0 62836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1624635492
transform 1 0 62284 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_662
timestamp 1624635492
transform 1 0 62008 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output457_A
timestamp 1624635492
transform 1 0 62100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input295_A
timestamp 1624635492
transform -1 0 63112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1598
timestamp 1624635492
transform 1 0 63848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_555
timestamp 1624635492
transform 1 0 52164 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_549
timestamp 1624635492
transform 1 0 51612 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output556_A
timestamp 1624635492
transform -1 0 52716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output552_A
timestamp 1624635492
transform -1 0 52164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output544_A
timestamp 1624635492
transform 1 0 51428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_568
timestamp 1624635492
transform 1 0 53360 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_565
timestamp 1624635492
transform 1 0 53084 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_561
timestamp 1624635492
transform 1 0 52716 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output561_A
timestamp 1624635492
transform 1 0 53176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_578
timestamp 1624635492
transform 1 0 54280 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output563_A
timestamp 1624635492
transform 1 0 54096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_596
timestamp 1624635492
transform 1 0 55936 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_590
timestamp 1624635492
transform 1 0 55384 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1602
timestamp 1624635492
transform 1 0 56028 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_610
timestamp 1624635492
transform 1 0 57224 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_598
timestamp 1624635492
transform 1 0 56120 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_622
timestamp 1624635492
transform 1 0 58328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_634
timestamp 1624635492
transform 1 0 59432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_646
timestamp 1624635492
transform 1 0 60536 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_655
timestamp 1624635492
transform 1 0 61364 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1603
timestamp 1624635492
transform 1 0 61272 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_673
timestamp 1624635492
transform 1 0 63020 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_667
timestamp 1624635492
transform 1 0 62468 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_663
timestamp 1624635492
transform 1 0 62100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output472_A
timestamp 1624635492
transform 1 0 62284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output459_A
timestamp 1624635492
transform 1 0 62836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_679
timestamp 1624635492
transform 1 0 63572 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output452_A
timestamp 1624635492
transform 1 0 63388 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_548
timestamp 1624635492
transform 1 0 51520 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_569
timestamp 1624635492
transform 1 0 53452 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_560
timestamp 1624635492
transform 1 0 52624 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1607
timestamp 1624635492
transform 1 0 53360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_581
timestamp 1624635492
transform 1 0 54556 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_593
timestamp 1624635492
transform 1 0 55660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_605
timestamp 1624635492
transform 1 0 56764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1624635492
transform 1 0 57868 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_626
timestamp 1624635492
transform 1 0 58696 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1608
timestamp 1624635492
transform 1 0 58604 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_638
timestamp 1624635492
transform 1 0 59800 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_650
timestamp 1624635492
transform 1 0 60904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_674
timestamp 1624635492
transform 1 0 63112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_662
timestamp 1624635492
transform 1 0 62008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_678
timestamp 1624635492
transform 1 0 63480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output471_A
timestamp 1624635492
transform 1 0 63296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1609
timestamp 1624635492
transform 1 0 63848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_548
timestamp 1624635492
transform 1 0 51520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_553
timestamp 1624635492
transform 1 0 51980 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_569
timestamp 1624635492
transform 1 0 53452 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_560
timestamp 1624635492
transform 1 0 52624 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_565
timestamp 1624635492
transform 1 0 53084 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1618
timestamp 1624635492
transform 1 0 53360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_581
timestamp 1624635492
transform 1 0 54556 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_577
timestamp 1624635492
transform 1 0 54188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_593
timestamp 1624635492
transform 1 0 55660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_589
timestamp 1624635492
transform 1 0 55292 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1613
timestamp 1624635492
transform 1 0 56028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_605
timestamp 1624635492
transform 1 0 56764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_610
timestamp 1624635492
transform 1 0 57224 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_598
timestamp 1624635492
transform 1 0 56120 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1624635492
transform 1 0 57868 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_622
timestamp 1624635492
transform 1 0 58328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_626
timestamp 1624635492
transform 1 0 58696 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_634
timestamp 1624635492
transform 1 0 59432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1619
timestamp 1624635492
transform 1 0 58604 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_638
timestamp 1624635492
transform 1 0 59800 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_646
timestamp 1624635492
transform 1 0 60536 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_650
timestamp 1624635492
transform 1 0 60904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_655
timestamp 1624635492
transform 1 0 61364 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1614
timestamp 1624635492
transform 1 0 61272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_674
timestamp 1624635492
transform 1 0 63112 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_662
timestamp 1624635492
transform 1 0 62008 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_667
timestamp 1624635492
transform 1 0 62468 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_679
timestamp 1624635492
transform 1 0 63572 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output461_A
timestamp 1624635492
transform 1 0 63848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1620
timestamp 1624635492
transform 1 0 63848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_553
timestamp 1624635492
transform 1 0 51980 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_565
timestamp 1624635492
transform 1 0 53084 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_577
timestamp 1624635492
transform 1 0 54188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_589
timestamp 1624635492
transform 1 0 55292 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1624
timestamp 1624635492
transform 1 0 56028 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_610
timestamp 1624635492
transform 1 0 57224 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_598
timestamp 1624635492
transform 1 0 56120 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_622
timestamp 1624635492
transform 1 0 58328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_634
timestamp 1624635492
transform 1 0 59432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_646
timestamp 1624635492
transform 1 0 60536 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_655
timestamp 1624635492
transform 1 0 61364 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1625
timestamp 1624635492
transform 1 0 61272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_667
timestamp 1624635492
transform 1 0 62468 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_679
timestamp 1624635492
transform 1 0 63572 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_548
timestamp 1624635492
transform 1 0 51520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_569
timestamp 1624635492
transform 1 0 53452 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_560
timestamp 1624635492
transform 1 0 52624 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1629
timestamp 1624635492
transform 1 0 53360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_581
timestamp 1624635492
transform 1 0 54556 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_593
timestamp 1624635492
transform 1 0 55660 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_605
timestamp 1624635492
transform 1 0 56764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1624635492
transform 1 0 57868 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_626
timestamp 1624635492
transform 1 0 58696 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1630
timestamp 1624635492
transform 1 0 58604 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_638
timestamp 1624635492
transform 1 0 59800 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_650
timestamp 1624635492
transform 1 0 60904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_674
timestamp 1624635492
transform 1 0 63112 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_662
timestamp 1624635492
transform 1 0 62008 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1631
timestamp 1624635492
transform 1 0 63848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_553
timestamp 1624635492
transform 1 0 51980 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_565
timestamp 1624635492
transform 1 0 53084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_577
timestamp 1624635492
transform 1 0 54188 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_589
timestamp 1624635492
transform 1 0 55292 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1635
timestamp 1624635492
transform 1 0 56028 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_610
timestamp 1624635492
transform 1 0 57224 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_598
timestamp 1624635492
transform 1 0 56120 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_622
timestamp 1624635492
transform 1 0 58328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_634
timestamp 1624635492
transform 1 0 59432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_646
timestamp 1624635492
transform 1 0 60536 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_655
timestamp 1624635492
transform 1 0 61364 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1636
timestamp 1624635492
transform 1 0 61272 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_667
timestamp 1624635492
transform 1 0 62468 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_679
timestamp 1624635492
transform 1 0 63572 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_548
timestamp 1624635492
transform 1 0 51520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_569
timestamp 1624635492
transform 1 0 53452 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_560
timestamp 1624635492
transform 1 0 52624 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1640
timestamp 1624635492
transform 1 0 53360 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_576
timestamp 1624635492
transform 1 0 54096 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _326_
timestamp 1624635492
transform -1 0 54096 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_588
timestamp 1624635492
transform 1 0 55200 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_600
timestamp 1624635492
transform 1 0 56304 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_612
timestamp 1624635492
transform 1 0 57408 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_626
timestamp 1624635492
transform 1 0 58696 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_624
timestamp 1624635492
transform 1 0 58512 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1641
timestamp 1624635492
transform 1 0 58604 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_638
timestamp 1624635492
transform 1 0 59800 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_650
timestamp 1624635492
transform 1 0 60904 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_674
timestamp 1624635492
transform 1 0 63112 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_662
timestamp 1624635492
transform 1 0 62008 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1642
timestamp 1624635492
transform 1 0 63848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_553
timestamp 1624635492
transform 1 0 51980 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_565
timestamp 1624635492
transform 1 0 53084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_577
timestamp 1624635492
transform 1 0 54188 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_589
timestamp 1624635492
transform 1 0 55292 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1646
timestamp 1624635492
transform 1 0 56028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_610
timestamp 1624635492
transform 1 0 57224 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_598
timestamp 1624635492
transform 1 0 56120 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_622
timestamp 1624635492
transform 1 0 58328 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_634
timestamp 1624635492
transform 1 0 59432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_646
timestamp 1624635492
transform 1 0 60536 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_655
timestamp 1624635492
transform 1 0 61364 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1647
timestamp 1624635492
transform 1 0 61272 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_667
timestamp 1624635492
transform 1 0 62468 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_679
timestamp 1624635492
transform 1 0 63572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_553
timestamp 1624635492
transform 1 0 51980 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_548
timestamp 1624635492
transform 1 0 51520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_565
timestamp 1624635492
transform 1 0 53084 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_569
timestamp 1624635492
transform 1 0 53452 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_560
timestamp 1624635492
transform 1 0 52624 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1651
timestamp 1624635492
transform 1 0 53360 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_577
timestamp 1624635492
transform 1 0 54188 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_581
timestamp 1624635492
transform 1 0 54556 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_589
timestamp 1624635492
transform 1 0 55292 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_593
timestamp 1624635492
transform 1 0 55660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1657
timestamp 1624635492
transform 1 0 56028 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_610
timestamp 1624635492
transform 1 0 57224 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_598
timestamp 1624635492
transform 1 0 56120 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_605
timestamp 1624635492
transform 1 0 56764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_622
timestamp 1624635492
transform 1 0 58328 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1624635492
transform 1 0 57868 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_634
timestamp 1624635492
transform 1 0 59432 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_626
timestamp 1624635492
transform 1 0 58696 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1652
timestamp 1624635492
transform 1 0 58604 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_646
timestamp 1624635492
transform 1 0 60536 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_638
timestamp 1624635492
transform 1 0 59800 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_655
timestamp 1624635492
transform 1 0 61364 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_650
timestamp 1624635492
transform 1 0 60904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1658
timestamp 1624635492
transform 1 0 61272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_667
timestamp 1624635492
transform 1 0 62468 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_674
timestamp 1624635492
transform 1 0 63112 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_662
timestamp 1624635492
transform 1 0 62008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_679
timestamp 1624635492
transform 1 0 63572 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1653
timestamp 1624635492
transform 1 0 63848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_548
timestamp 1624635492
transform 1 0 51520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_569
timestamp 1624635492
transform 1 0 53452 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_560
timestamp 1624635492
transform 1 0 52624 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1662
timestamp 1624635492
transform 1 0 53360 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_581
timestamp 1624635492
transform 1 0 54556 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_593
timestamp 1624635492
transform 1 0 55660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_605
timestamp 1624635492
transform 1 0 56764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1624635492
transform 1 0 57868 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_626
timestamp 1624635492
transform 1 0 58696 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1663
timestamp 1624635492
transform 1 0 58604 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_638
timestamp 1624635492
transform 1 0 59800 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_650
timestamp 1624635492
transform 1 0 60904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_674
timestamp 1624635492
transform 1 0 63112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_662
timestamp 1624635492
transform 1 0 62008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1664
timestamp 1624635492
transform 1 0 63848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_553
timestamp 1624635492
transform 1 0 51980 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_565
timestamp 1624635492
transform 1 0 53084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_577
timestamp 1624635492
transform 1 0 54188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_589
timestamp 1624635492
transform 1 0 55292 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1668
timestamp 1624635492
transform 1 0 56028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_610
timestamp 1624635492
transform 1 0 57224 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_598
timestamp 1624635492
transform 1 0 56120 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_622
timestamp 1624635492
transform 1 0 58328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_634
timestamp 1624635492
transform 1 0 59432 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_646
timestamp 1624635492
transform 1 0 60536 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_655
timestamp 1624635492
transform 1 0 61364 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1669
timestamp 1624635492
transform 1 0 61272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_667
timestamp 1624635492
transform 1 0 62468 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_679
timestamp 1624635492
transform 1 0 63572 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_548
timestamp 1624635492
transform 1 0 51520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_569
timestamp 1624635492
transform 1 0 53452 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_560
timestamp 1624635492
transform 1 0 52624 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1673
timestamp 1624635492
transform 1 0 53360 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_581
timestamp 1624635492
transform 1 0 54556 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_597
timestamp 1624635492
transform 1 0 56028 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_593
timestamp 1624635492
transform 1 0 55660 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_600
timestamp 1624635492
transform 1 0 56304 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__B
timestamp 1624635492
transform 1 0 56120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_612
timestamp 1624635492
transform 1 0 57408 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_626
timestamp 1624635492
transform 1 0 58696 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_624
timestamp 1624635492
transform 1 0 58512 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1674
timestamp 1624635492
transform 1 0 58604 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_638
timestamp 1624635492
transform 1 0 59800 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_650
timestamp 1624635492
transform 1 0 60904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_674
timestamp 1624635492
transform 1 0 63112 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_662
timestamp 1624635492
transform 1 0 62008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1675
timestamp 1624635492
transform 1 0 63848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_553
timestamp 1624635492
transform 1 0 51980 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_565
timestamp 1624635492
transform 1 0 53084 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_577
timestamp 1624635492
transform 1 0 54188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_589
timestamp 1624635492
transform 1 0 55292 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1679
timestamp 1624635492
transform 1 0 56028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_605
timestamp 1624635492
transform 1 0 56764 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_598
timestamp 1624635492
transform 1 0 56120 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1624635492
transform 1 0 57132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 56488 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_623
timestamp 1624635492
transform 1 0 58420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_611
timestamp 1624635492
transform 1 0 57316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_635
timestamp 1624635492
transform 1 0 59524 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_647
timestamp 1624635492
transform 1 0 60628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_655
timestamp 1624635492
transform 1 0 61364 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_653
timestamp 1624635492
transform 1 0 61180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1680
timestamp 1624635492
transform 1 0 61272 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_667
timestamp 1624635492
transform 1 0 62468 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_679
timestamp 1624635492
transform 1 0 63572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_688
timestamp 1624635492
transform 1 0 64400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_683
timestamp 1624635492
transform 1 0 63940 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output454
timestamp 1624635492
transform -1 0 65136 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1537
timestamp 1624635492
transform 1 0 64308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_704
timestamp 1624635492
transform 1 0 65872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_696
timestamp 1624635492
transform 1 0 65136 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output458
timestamp 1624635492
transform -1 0 66608 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output456
timestamp 1624635492
transform -1 0 65872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_719
timestamp 1624635492
transform 1 0 67252 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_712
timestamp 1624635492
transform 1 0 66608 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 67252 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1538
timestamp 1624635492
transform 1 0 66976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1624635492
transform 1 0 68172 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output406
timestamp 1624635492
transform 1 0 67804 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1624635492
transform -1 0 68816 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_692
timestamp 1624635492
transform 1 0 64768 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_688
timestamp 1624635492
transform 1 0 64400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_691
timestamp 1624635492
transform 1 0 64676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_683
timestamp 1624635492
transform 1 0 63940 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output463
timestamp 1624635492
transform -1 0 65228 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output462
timestamp 1624635492
transform -1 0 65412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output461
timestamp 1624635492
transform -1 0 64400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output460
timestamp 1624635492
transform -1 0 64676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_707
timestamp 1624635492
transform 1 0 66148 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_697
timestamp 1624635492
transform 1 0 65228 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_707
timestamp 1624635492
transform 1 0 66148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_699
timestamp 1624635492
transform 1 0 65412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output472
timestamp 1624635492
transform 1 0 65780 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output464
timestamp 1624635492
transform -1 0 66148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_720
timestamp 1624635492
transform 1 0 67344 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_712
timestamp 1624635492
transform 1 0 66608 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_721
timestamp 1624635492
transform 1 0 67436 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_715
timestamp 1624635492
transform 1 0 66884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform 1 0 67252 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output467
timestamp 1624635492
transform -1 0 67344 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output465
timestamp 1624635492
transform -1 0 66884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1549
timestamp 1624635492
transform 1 0 66516 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_732
timestamp 1624635492
transform 1 0 68448 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_728
timestamp 1624635492
transform 1 0 68080 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1624635492
transform 1 0 68172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output469
timestamp 1624635492
transform -1 0 68080 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output368
timestamp 1624635492
transform 1 0 67804 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1624635492
transform -1 0 68816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1624635492
transform -1 0 68816 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_690
timestamp 1624635492
transform 1 0 64584 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_683
timestamp 1624635492
transform 1 0 63940 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1624635492
transform 1 0 64308 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_708
timestamp 1624635492
transform 1 0 66240 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_700
timestamp 1624635492
transform 1 0 65504 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_696
timestamp 1624635492
transform 1 0 65136 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output572
timestamp 1624635492
transform 1 0 65872 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform -1 0 65504 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_720
timestamp 1624635492
transform 1 0 67344 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_716
timestamp 1624635492
transform 1 0 66976 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output470
timestamp 1624635492
transform -1 0 67804 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output468
timestamp 1624635492
transform -1 0 66976 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_725
timestamp 1624635492
transform 1 0 67804 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1624635492
transform -1 0 68816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_692
timestamp 1624635492
transform 1 0 64768 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_685
timestamp 1624635492
transform 1 0 64124 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1624635492
transform -1 0 64768 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_706
timestamp 1624635492
transform 1 0 66056 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_699
timestamp 1624635492
transform 1 0 65412 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1624635492
transform -1 0 66056 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1624635492
transform 1 0 65136 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_721
timestamp 1624635492
transform 1 0 67436 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_716
timestamp 1624635492
transform 1 0 66976 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_712
timestamp 1624635492
transform 1 0 66608 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_710
timestamp 1624635492
transform 1 0 66424 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output474
timestamp 1624635492
transform 1 0 67068 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1560
timestamp 1624635492
transform 1 0 66516 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_729
timestamp 1624635492
transform 1 0 68172 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output471
timestamp 1624635492
transform -1 0 68172 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1624635492
transform -1 0 68816 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_690
timestamp 1624635492
transform 1 0 64584 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_683
timestamp 1624635492
transform 1 0 63940 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input183
timestamp 1624635492
transform 1 0 64308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1624635492
transform -1 0 65228 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_704
timestamp 1624635492
transform 1 0 65872 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_697
timestamp 1624635492
transform 1 0 65228 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1624635492
transform -1 0 66516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1624635492
transform -1 0 65872 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_721
timestamp 1624635492
transform 1 0 67436 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_711
timestamp 1624635492
transform 1 0 66516 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output573
timestamp 1624635492
transform 1 0 67068 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1624635492
transform 1 0 68172 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output473
timestamp 1624635492
transform 1 0 67804 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1624635492
transform -1 0 68816 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_688
timestamp 1624635492
transform 1 0 64400 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input184
timestamp 1624635492
transform -1 0 64400 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_707
timestamp 1624635492
transform 1 0 66148 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_700
timestamp 1624635492
transform 1 0 65504 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_696
timestamp 1624635492
transform 1 0 65136 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1624635492
transform -1 0 65504 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1624635492
transform -1 0 66148 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_721
timestamp 1624635492
transform 1 0 67436 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_716
timestamp 1624635492
transform 1 0 66976 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_712
timestamp 1624635492
transform 1 0 66608 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output574
timestamp 1624635492
transform 1 0 67068 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1571
timestamp 1624635492
transform 1 0 66516 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_729
timestamp 1624635492
transform 1 0 68172 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output417
timestamp 1624635492
transform 1 0 67804 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1624635492
transform -1 0 68816 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 64216 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 64308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_683
timestamp 1624635492
transform 1 0 63940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_686
timestamp 1624635492
transform 1 0 64216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_687
timestamp 1624635492
transform 1 0 64308 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input185
timestamp 1624635492
transform -1 0 64860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input195
timestamp 1624635492
transform -1 0 65044 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_691
timestamp 1624635492
transform 1 0 64676 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_693
timestamp 1624635492
transform 1 0 64860 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_695
timestamp 1624635492
transform 1 0 65044 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_702
timestamp 1624635492
transform 1 0 65688 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_706
timestamp 1624635492
transform 1 0 66056 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_700
timestamp 1624635492
transform 1 0 65504 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 66056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input187
timestamp 1624635492
transform -1 0 65688 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input186
timestamp 1624635492
transform 1 0 65228 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1582
timestamp 1624635492
transform 1 0 66516 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1624635492
transform -1 0 66700 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 66884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_713
timestamp 1624635492
transform 1 0 66700 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_710
timestamp 1624635492
transform 1 0 66424 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_712
timestamp 1624635492
transform 1 0 66608 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1624635492
transform 1 0 67068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1624635492
transform -1 0 67528 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_715
timestamp 1624635492
transform 1 0 66884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_720
timestamp 1624635492
transform 1 0 67344 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_729
timestamp 1624635492
transform 1 0 68172 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_722
timestamp 1624635492
transform 1 0 67528 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1624635492
transform 1 0 68172 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1624635492
transform 1 0 67896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1624635492
transform -1 0 68172 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1624635492
transform -1 0 68816 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1624635492
transform -1 0 68816 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_693
timestamp 1624635492
transform 1 0 64860 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_685
timestamp 1624635492
transform 1 0 64124 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input182_A
timestamp 1624635492
transform -1 0 64124 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 64860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_707
timestamp 1624635492
transform 1 0 66148 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_700
timestamp 1624635492
transform 1 0 65504 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input197
timestamp 1624635492
transform -1 0 65504 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input188
timestamp 1624635492
transform -1 0 66148 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_721
timestamp 1624635492
transform 1 0 67436 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_714
timestamp 1624635492
transform 1 0 66792 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input191
timestamp 1624635492
transform 1 0 67160 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input190
timestamp 1624635492
transform -1 0 66792 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1624635492
transform 1 0 68172 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output379
timestamp 1624635492
transform 1 0 67804 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1624635492
transform -1 0 68816 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_694
timestamp 1624635492
transform 1 0 64952 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_691
timestamp 1624635492
transform 1 0 64676 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_687
timestamp 1624635492
transform 1 0 64308 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input183_A
timestamp 1624635492
transform -1 0 64308 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1624635492
transform -1 0 64952 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_706
timestamp 1624635492
transform 1 0 66056 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_700
timestamp 1624635492
transform 1 0 65504 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1624635492
transform -1 0 65504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 66056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_721
timestamp 1624635492
transform 1 0 67436 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_714
timestamp 1624635492
transform 1 0 66792 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_710
timestamp 1624635492
transform 1 0 66424 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624635492
transform -1 0 66792 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input192
timestamp 1624635492
transform -1 0 67436 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1593
timestamp 1624635492
transform 1 0 66516 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_732
timestamp 1624635492
transform 1 0 68448 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_728
timestamp 1624635492
transform 1 0 68080 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input193
timestamp 1624635492
transform -1 0 68080 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1624635492
transform -1 0 68816 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_690
timestamp 1624635492
transform 1 0 64584 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_687
timestamp 1624635492
transform 1 0 64308 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_683
timestamp 1624635492
transform 1 0 63940 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input185_A
timestamp 1624635492
transform -1 0 65136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input184_A
timestamp 1624635492
transform -1 0 64584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_706
timestamp 1624635492
transform 1 0 66056 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_702
timestamp 1624635492
transform 1 0 65688 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_696
timestamp 1624635492
transform 1 0 65136 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1624635492
transform -1 0 65688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1624635492
transform -1 0 66332 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_715
timestamp 1624635492
transform 1 0 66884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_709
timestamp 1624635492
transform 1 0 66332 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1624635492
transform -1 0 66884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input194
timestamp 1624635492
transform -1 0 67528 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1624635492
transform 1 0 68172 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_722
timestamp 1624635492
transform 1 0 67528 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1624635492
transform -1 0 68172 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1624635492
transform -1 0 68816 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_691
timestamp 1624635492
transform 1 0 64676 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_685
timestamp 1624635492
transform 1 0 64124 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output406_A
timestamp 1624635492
transform 1 0 63940 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output379_A
timestamp 1624635492
transform 1 0 64492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input186_A
timestamp 1624635492
transform -1 0 65228 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_704
timestamp 1624635492
transform 1 0 65872 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_701
timestamp 1624635492
transform 1 0 65596 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_697
timestamp 1624635492
transform 1 0 65228 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input187_A
timestamp 1624635492
transform -1 0 65872 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_716
timestamp 1624635492
transform 1 0 66976 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_712
timestamp 1624635492
transform 1 0 66608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_710
timestamp 1624635492
transform 1 0 66424 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1624635492
transform -1 0 66976 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 67528 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1604
timestamp 1624635492
transform 1 0 66516 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_729
timestamp 1624635492
transform 1 0 68172 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_722
timestamp 1624635492
transform 1 0 67528 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input196
timestamp 1624635492
transform -1 0 68172 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1624635492
transform -1 0 68816 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_691
timestamp 1624635492
transform 1 0 64676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_685
timestamp 1624635492
transform 1 0 64124 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output460_A
timestamp 1624635492
transform 1 0 63940 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output454_A
timestamp 1624635492
transform 1 0 64492 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input197_A
timestamp 1624635492
transform -1 0 65228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_703
timestamp 1624635492
transform 1 0 65780 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_697
timestamp 1624635492
transform 1 0 65228 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input196_A
timestamp 1624635492
transform -1 0 65780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input188_A
timestamp 1624635492
transform -1 0 66332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_721
timestamp 1624635492
transform 1 0 67436 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_715
timestamp 1624635492
transform 1 0 66884 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_709
timestamp 1624635492
transform 1 0 66332 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input190_A
timestamp 1624635492
transform -1 0 66884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_732
timestamp 1624635492
transform 1 0 68448 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_724
timestamp 1624635492
transform 1 0 67712 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1624635492
transform -1 0 67712 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1624635492
transform -1 0 68816 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_693
timestamp 1624635492
transform 1 0 64860 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_683
timestamp 1624635492
transform 1 0 63940 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_694
timestamp 1624635492
transform 1 0 64952 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_684
timestamp 1624635492
transform 1 0 64032 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output463_A
timestamp 1624635492
transform 1 0 64676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output462_A
timestamp 1624635492
transform 1 0 64768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output456_A
timestamp 1624635492
transform -1 0 65504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output464_A
timestamp 1624635492
transform 1 0 65504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_700
timestamp 1624635492
transform 1 0 65504 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_699
timestamp 1624635492
transform 1 0 65412 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_702
timestamp 1624635492
transform 1 0 65688 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output368_A
timestamp 1624635492
transform 1 0 65964 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output458_A
timestamp 1624635492
transform 1 0 66056 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_704
timestamp 1624635492
transform 1 0 65872 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_707
timestamp 1624635492
transform 1 0 66148 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_708
timestamp 1624635492
transform 1 0 66240 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_717
timestamp 1624635492
transform 1 0 67068 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_714
timestamp 1624635492
transform 1 0 66792 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_718
timestamp 1624635492
transform 1 0 67160 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_712
timestamp 1624635492
transform 1 0 66608 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input194_A
timestamp 1624635492
transform -1 0 67068 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input192_A
timestamp 1624635492
transform -1 0 67620 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input191_A
timestamp 1624635492
transform -1 0 67160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1615
timestamp 1624635492
transform 1 0 66516 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1624635492
transform 1 0 68172 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_723
timestamp 1624635492
transform 1 0 67620 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_729
timestamp 1624635492
transform 1 0 68172 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_724
timestamp 1624635492
transform 1 0 67712 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input193_A
timestamp 1624635492
transform -1 0 68172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output428
timestamp 1624635492
transform 1 0 67804 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1624635492
transform -1 0 68816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1624635492
transform -1 0 68816 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_691
timestamp 1624635492
transform 1 0 64676 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_707
timestamp 1624635492
transform 1 0 66148 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_701
timestamp 1624635492
transform 1 0 65596 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output574_A
timestamp 1624635492
transform 1 0 65412 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output468_A
timestamp 1624635492
transform 1 0 65964 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_721
timestamp 1624635492
transform 1 0 67436 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_715
timestamp 1624635492
transform 1 0 66884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_712
timestamp 1624635492
transform 1 0 66608 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output467_A
timestamp 1624635492
transform 1 0 66700 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output390_A
timestamp 1624635492
transform -1 0 67436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1626
timestamp 1624635492
transform 1 0 66516 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_729
timestamp 1624635492
transform 1 0 68172 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output390
timestamp 1624635492
transform 1 0 67804 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1624635492
transform -1 0 68816 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_695
timestamp 1624635492
transform 1 0 65044 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_683
timestamp 1624635492
transform 1 0 63940 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_707
timestamp 1624635492
transform 1 0 66148 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_703
timestamp 1624635492
transform 1 0 65780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output573_A
timestamp 1624635492
transform 1 0 65964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_719
timestamp 1624635492
transform 1 0 67252 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_713
timestamp 1624635492
transform 1 0 66700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output470_A
timestamp 1624635492
transform -1 0 66700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output469_A
timestamp 1624635492
transform 1 0 67068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_725
timestamp 1624635492
transform 1 0 67804 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output428_A
timestamp 1624635492
transform -1 0 67804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1624635492
transform -1 0 68816 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_691
timestamp 1624635492
transform 1 0 64676 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_703
timestamp 1624635492
transform 1 0 65780 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_712
timestamp 1624635492
transform 1 0 66608 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 67528 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1637
timestamp 1624635492
transform 1 0 66516 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_729
timestamp 1624635492
transform 1 0 68172 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_722
timestamp 1624635492
transform 1 0 67528 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1624635492
transform -1 0 68172 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1624635492
transform -1 0 68816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_695
timestamp 1624635492
transform 1 0 65044 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_683
timestamp 1624635492
transform 1 0 63940 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_707
timestamp 1624635492
transform 1 0 66148 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_719
timestamp 1624635492
transform 1 0 67252 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_731
timestamp 1624635492
transform 1 0 68356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_279
timestamp 1624635492
transform -1 0 68816 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_691
timestamp 1624635492
transform 1 0 64676 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_703
timestamp 1624635492
transform 1 0 65780 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_712
timestamp 1624635492
transform 1 0 66608 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1648
timestamp 1624635492
transform 1 0 66516 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_732
timestamp 1624635492
transform 1 0 68448 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_724
timestamp 1624635492
transform 1 0 67712 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_281
timestamp 1624635492
transform -1 0 68816 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_691
timestamp 1624635492
transform 1 0 64676 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_695
timestamp 1624635492
transform 1 0 65044 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_683
timestamp 1624635492
transform 1 0 63940 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_703
timestamp 1624635492
transform 1 0 65780 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_707
timestamp 1624635492
transform 1 0 66148 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_712
timestamp 1624635492
transform 1 0 66608 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_721
timestamp 1624635492
transform 1 0 67436 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output437_A
timestamp 1624635492
transform 1 0 67252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1659
timestamp 1624635492
transform 1 0 66516 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_727
timestamp 1624635492
transform 1 0 67988 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1624635492
transform 1 0 68172 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output437
timestamp 1624635492
transform 1 0 67804 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_285
timestamp 1624635492
transform -1 0 68816 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_283
timestamp 1624635492
transform -1 0 68816 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _286_
timestamp 1624635492
transform -1 0 67988 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_695
timestamp 1624635492
transform 1 0 65044 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_683
timestamp 1624635492
transform 1 0 63940 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_707
timestamp 1624635492
transform 1 0 66148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_721
timestamp 1624635492
transform 1 0 67436 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_712
timestamp 1624635492
transform 1 0 66608 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _247_
timestamp 1624635492
transform -1 0 66608 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _206_
timestamp 1624635492
transform -1 0 67436 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1624635492
transform 1 0 68172 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output399
timestamp 1624635492
transform 1 0 67804 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_287
timestamp 1624635492
transform -1 0 68816 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_691
timestamp 1624635492
transform 1 0 64676 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_703
timestamp 1624635492
transform 1 0 65780 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_720
timestamp 1624635492
transform 1 0 67344 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_712
timestamp 1624635492
transform 1 0 66608 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1670
timestamp 1624635492
transform 1 0 66516 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1624635492
transform 1 0 67804 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output399_A
timestamp 1624635492
transform 1 0 67620 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_289
timestamp 1624635492
transform -1 0 68816 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_695
timestamp 1624635492
transform 1 0 65044 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_683
timestamp 1624635492
transform 1 0 63940 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_707
timestamp 1624635492
transform 1 0 66148 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_719
timestamp 1624635492
transform 1 0 67252 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_731
timestamp 1624635492
transform 1 0 68356 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_291
timestamp 1624635492
transform -1 0 68816 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_691
timestamp 1624635492
transform 1 0 64676 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_703
timestamp 1624635492
transform 1 0 65780 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_712
timestamp 1624635492
transform 1 0 66608 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 67528 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1681
timestamp 1624635492
transform 1 0 66516 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_729
timestamp 1624635492
transform 1 0 68172 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_722
timestamp 1624635492
transform 1 0 67528 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1624635492
transform -1 0 68172 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_293
timestamp 1624635492
transform -1 0 68816 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1624635492
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1624635492
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1624635492
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1624635492
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1624635492
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1624635492
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_94
timestamp 1624635492
transform 1 0 9752 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1624635492
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _282_
timestamp 1624635492
transform 1 0 9844 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_110
timestamp 1624635492
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_127
timestamp 1624635492
transform 1 0 12788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1624635492
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1624635492
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1624635492
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1624635492
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1624635492
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1624635492
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1624635492
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1624635492
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1624635492
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1624635492
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1624635492
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1624635492
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1624635492
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1624635492
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_51
timestamp 1624635492
transform 1 0 5796 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1624635492
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1624635492
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1624635492
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1624635492
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1624635492
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1624635492
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1624635492
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_17
timestamp 1624635492
transform 1 0 2668 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_11
timestamp 1624635492
transform 1 0 2116 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output394_A
timestamp 1624635492
transform -1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output394
timestamp 1624635492
transform -1 0 2116 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1624635492
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1624635492
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1624635492
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_54
timestamp 1624635492
transform 1 0 6072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1624635492
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1624635492
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1624635492
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1624635492
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1624635492
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1624635492
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_94
timestamp 1624635492
transform 1 0 9752 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _173_
timestamp 1624635492
transform -1 0 9752 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1624635492
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1624635492
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_118
timestamp 1624635492
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_106
timestamp 1624635492
transform 1 0 10856 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1624635492
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_130
timestamp 1624635492
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_17
timestamp 1624635492
transform 1 0 2668 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1624635492
transform 1 0 2116 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1624635492
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output432_A
timestamp 1624635492
transform -1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output432
timestamp 1624635492
transform -1 0 2116 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_59
timestamp 1624635492
transform 1 0 6532 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1624635492
transform 1 0 6072 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1624635492
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1624635492
transform 1 0 6440 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_71
timestamp 1624635492
transform 1 0 7636 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_88
timestamp 1624635492
transform 1 0 9200 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_83
timestamp 1624635492
transform 1 0 8740 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1624635492
transform 1 0 9108 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1624635492
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_112
timestamp 1624635492
transform 1 0 11408 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_100
timestamp 1624635492
transform 1 0 10304 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1624635492
transform 1 0 11776 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1624635492
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1624635492
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1624635492
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1624635492
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1624635492
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1624635492
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1624635492
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1624635492
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1624635492
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1624635492
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1624635492
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1624635492
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1624635492
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_17
timestamp 1624635492
transform 1 0 2668 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_5
timestamp 1624635492
transform 1 0 1564 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1624635492
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1624635492
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1624635492
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1624635492
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_78
timestamp 1624635492
transform 1 0 8280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1624635492
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1624635492
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1624635492
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1624635492
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1624635492
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1624635492
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1624635492
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1624635492
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_6
timestamp 1624635492
transform 1 0 1656 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1624635492
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1624635492
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _186_
timestamp 1624635492
transform 1 0 2208 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1624635492
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1624635492
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1624635492
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_51
timestamp 1624635492
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1624635492
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1624635492
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1624635492
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1624635492
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1624635492
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1624635492
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1624635492
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_131
timestamp 1624635492
transform 1 0 13156 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_127
timestamp 1624635492
transform 1 0 12788 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _159_
timestamp 1624635492
transform 1 0 12880 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1624635492
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1624635492
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1624635492
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1624635492
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1624635492
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1624635492
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1624635492
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1624635492
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1624635492
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1624635492
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_99
timestamp 1624635492
transform 1 0 10212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1624635492
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1624635492
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_111
timestamp 1624635492
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1624635492
transform 1 0 13524 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1624635492
transform 1 0 12420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1624635492
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1624635492
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1624635492
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1624635492
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1624635492
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1624635492
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1624635492
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1624635492
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1624635492
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1624635492
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1624635492
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1624635492
transform 1 0 6072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1624635492
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_58
timestamp 1624635492
transform 1 0 6440 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_51
timestamp 1624635492
transform 1 0 5796 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1624635492
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_78
timestamp 1624635492
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1624635492
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _346_
timestamp 1624635492
transform 1 0 6992 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_38_99
timestamp 1624635492
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_87
timestamp 1624635492
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_95
timestamp 1624635492
transform 1 0 9844 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_89
timestamp 1624635492
transform 1 0 9292 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_83
timestamp 1624635492
transform 1 0 8740 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__CLK
timestamp 1624635492
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__D
timestamp 1624635492
transform -1 0 9292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1624635492
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_116
timestamp 1624635492
transform 1 0 11776 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_111
timestamp 1624635492
transform 1 0 11316 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1624635492
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1624635492
transform 1 0 11500 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_107
timestamp 1624635492
transform 1 0 10948 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1624635492
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _259_
timestamp 1624635492
transform 1 0 11500 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_128
timestamp 1624635492
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_132
timestamp 1624635492
transform 1 0 13248 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1624635492
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _140_
timestamp 1624635492
transform 1 0 12972 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_17
timestamp 1624635492
transform 1 0 2668 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1624635492
transform 1 0 2116 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1624635492
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output393_A
timestamp 1624635492
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output393
timestamp 1624635492
transform -1 0 2116 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1624635492
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_29
timestamp 1624635492
transform 1 0 3772 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1624635492
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_53
timestamp 1624635492
transform 1 0 5980 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1624635492
transform 1 0 4876 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1624635492
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1624635492
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1624635492
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1624635492
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1624635492
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1624635492
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1624635492
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1624635492
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1624635492
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1624635492
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1624635492
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1624635492
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1624635492
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1624635492
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1624635492
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1624635492
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1624635492
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1624635492
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1624635492
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1624635492
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1624635492
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_119
timestamp 1624635492
transform 1 0 12052 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_111
timestamp 1624635492
transform 1 0 11316 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1624635492
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1624635492
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _196_
timestamp 1624635492
transform 1 0 12144 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1624635492
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1624635492
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1624635492
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1624635492
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1624635492
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1624635492
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_51
timestamp 1624635492
transform 1 0 5796 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1624635492
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1624635492
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1624635492
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1624635492
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_115
timestamp 1624635492
transform 1 0 11684 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1624635492
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1624635492
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1624635492
transform 1 0 12788 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_17
timestamp 1624635492
transform 1 0 2668 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1624635492
transform 1 0 2116 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1624635492
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output431_A
timestamp 1624635492
transform 1 0 2484 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output431
timestamp 1624635492
transform -1 0 2116 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1624635492
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1624635492
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1624635492
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1624635492
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1624635492
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1624635492
transform 1 0 8004 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_66
timestamp 1624635492
transform 1 0 7176 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _237_
timestamp 1624635492
transform 1 0 7728 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1624635492
transform 1 0 10212 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_87
timestamp 1624635492
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_83
timestamp 1624635492
transform 1 0 8740 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1624635492
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_119
timestamp 1624635492
transform 1 0 12052 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_113
timestamp 1624635492
transform 1 0 11500 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_103
timestamp 1624635492
transform 1 0 10580 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1624635492
transform 1 0 11868 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  _064_
timestamp 1624635492
transform -1 0 11500 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_42_131
timestamp 1624635492
transform 1 0 13156 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_8
timestamp 1624635492
transform 1 0 1840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1624635492
transform 1 0 1380 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1624635492
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1624635492
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1624635492
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1624635492
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _266_
timestamp 1624635492
transform 1 0 1564 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_30
timestamp 1624635492
transform 1 0 3864 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_28
timestamp 1624635492
transform 1 0 3680 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1624635492
transform 1 0 2944 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1624635492
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1624635492
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1624635492
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_54
timestamp 1624635492
transform 1 0 6072 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_42
timestamp 1624635492
transform 1 0 4968 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1624635492
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_51
timestamp 1624635492
transform 1 0 5796 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1624635492
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_78
timestamp 1624635492
transform 1 0 8280 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_66
timestamp 1624635492
transform 1 0 7176 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1624635492
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_99
timestamp 1624635492
transform 1 0 10212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_87
timestamp 1624635492
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1624635492
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1624635492
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1624635492
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_111
timestamp 1624635492
transform 1 0 11316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_115
timestamp 1624635492
transform 1 0 11684 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1624635492
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1624635492
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_135
timestamp 1624635492
transform 1 0 13524 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1624635492
transform 1 0 12420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1624635492
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_12
timestamp 1624635492
transform 1 0 2208 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1624635492
transform 1 0 1656 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 2208 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1624635492
transform -1 0 1656 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1624635492
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_36
timestamp 1624635492
transform 1 0 4416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_24
timestamp 1624635492
transform 1 0 3312 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_58
timestamp 1624635492
transform 1 0 6440 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_56
timestamp 1624635492
transform 1 0 6256 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1624635492
transform 1 0 5520 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1624635492
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_70
timestamp 1624635492
transform 1 0 7544 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_94
timestamp 1624635492
transform 1 0 9752 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_82
timestamp 1624635492
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_115
timestamp 1624635492
transform 1 0 11684 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1624635492
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1624635492
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1624635492
transform 1 0 12788 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1624635492
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1624635492
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1624635492
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1624635492
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_27
timestamp 1624635492
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1624635492
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1624635492
transform 1 0 6072 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1624635492
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_74
timestamp 1624635492
transform 1 0 7912 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_70
timestamp 1624635492
transform 1 0 7544 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_66
timestamp 1624635492
transform 1 0 7176 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _308_
timestamp 1624635492
transform -1 0 7912 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_99
timestamp 1624635492
transform 1 0 10212 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1624635492
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1624635492
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_111
timestamp 1624635492
transform 1 0 11316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_135
timestamp 1624635492
transform 1 0 13524 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_123
timestamp 1624635492
transform 1 0 12420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1624635492
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1624635492
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1624635492
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1624635492
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1624635492
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1624635492
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_51
timestamp 1624635492
transform 1 0 5796 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1624635492
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_70
timestamp 1624635492
transform 1 0 7544 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_94
timestamp 1624635492
transform 1 0 9752 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_82
timestamp 1624635492
transform 1 0 8648 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1624635492
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1624635492
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1624635492
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_135
timestamp 1624635492
transform 1 0 13524 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_131
timestamp 1624635492
transform 1 0 13156 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1624635492
transform 1 0 12788 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _158_
timestamp 1624635492
transform 1 0 13248 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1624635492
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1624635492
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1624635492
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_30
timestamp 1624635492
transform 1 0 3864 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1624635492
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1624635492
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_54
timestamp 1624635492
transform 1 0 6072 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_42
timestamp 1624635492
transform 1 0 4968 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_78
timestamp 1624635492
transform 1 0 8280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_66
timestamp 1624635492
transform 1 0 7176 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_99
timestamp 1624635492
transform 1 0 10212 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_87
timestamp 1624635492
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1624635492
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1624635492
transform 1 0 11316 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_135
timestamp 1624635492
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_123
timestamp 1624635492
transform 1 0 12420 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_17
timestamp 1624635492
transform 1 0 2668 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1624635492
transform 1 0 2116 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1624635492
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output392_A
timestamp 1624635492
transform 1 0 2484 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output392
timestamp 1624635492
transform -1 0 2116 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1624635492
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_29
timestamp 1624635492
transform 1 0 3772 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_58
timestamp 1624635492
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_53
timestamp 1624635492
transform 1 0 5980 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_41
timestamp 1624635492
transform 1 0 4876 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1624635492
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_70
timestamp 1624635492
transform 1 0 7544 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1624635492
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_82
timestamp 1624635492
transform 1 0 8648 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_115
timestamp 1624635492
transform 1 0 11684 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_106
timestamp 1624635492
transform 1 0 10856 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1624635492
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_127
timestamp 1624635492
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1624635492
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1624635492
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output430
timestamp 1624635492
transform -1 0 2116 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1624635492
transform 1 0 1380 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1624635492
transform 1 0 1380 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _114_
timestamp 1624635492
transform 1 0 2484 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output430_A
timestamp 1624635492
transform 1 0 2116 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_11
timestamp 1624635492
transform 1 0 2116 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_13
timestamp 1624635492
transform 1 0 2300 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_18
timestamp 1624635492
transform 1 0 2760 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1624635492
transform 1 0 3864 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1624635492
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_25
timestamp 1624635492
transform 1 0 3404 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1624635492
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_58
timestamp 1624635492
transform 1 0 6440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_54
timestamp 1624635492
transform 1 0 6072 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1624635492
transform 1 0 4968 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_54
timestamp 1624635492
transform 1 0 6072 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1624635492
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1624635492
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_70
timestamp 1624635492
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_77
timestamp 1624635492
transform 1 0 8188 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1624635492
transform 1 0 7084 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _197_
timestamp 1624635492
transform 1 0 6808 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_94
timestamp 1624635492
transform 1 0 9752 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_82
timestamp 1624635492
transform 1 0 8648 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_99
timestamp 1624635492
transform 1 0 10212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_87
timestamp 1624635492
transform 1 0 9108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_85
timestamp 1624635492
transform 1 0 8924 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1624635492
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_115
timestamp 1624635492
transform 1 0 11684 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_106
timestamp 1624635492
transform 1 0 10856 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_111
timestamp 1624635492
transform 1 0 11316 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1624635492
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _307_
timestamp 1624635492
transform -1 0 12328 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_134
timestamp 1624635492
transform 1 0 13432 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_122
timestamp 1624635492
transform 1 0 12328 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_135
timestamp 1624635492
transform 1 0 13524 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_123
timestamp 1624635492
transform 1 0 12420 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1624635492
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1624635492
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1624635492
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_37
timestamp 1624635492
transform 1 0 4508 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_30
timestamp 1624635492
transform 1 0 3864 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_27
timestamp 1624635492
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1624635492
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _172_
timestamp 1624635492
transform 1 0 4232 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_49
timestamp 1624635492
transform 1 0 5612 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_77
timestamp 1624635492
transform 1 0 8188 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_73
timestamp 1624635492
transform 1 0 7820 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_61
timestamp 1624635492
transform 1 0 6716 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _213_
timestamp 1624635492
transform 1 0 7912 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_99
timestamp 1624635492
transform 1 0 10212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1624635492
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_85
timestamp 1624635492
transform 1 0 8924 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1624635492
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_111
timestamp 1624635492
transform 1 0 11316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_135
timestamp 1624635492
transform 1 0 13524 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_123
timestamp 1624635492
transform 1 0 12420 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1624635492
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1624635492
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1624635492
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1624635492
transform 1 0 18308 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _219_
timestamp 1624635492
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 18952 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_168
timestamp 1624635492
transform 1 0 16560 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1624635492
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_8  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 16836 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1624635492
transform 1 0 18308 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 18952 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1624635492
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1624635492
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1624635492
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_187
timestamp 1624635492
transform 1 0 18308 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_181
timestamp 1624635492
transform 1 0 17756 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_178
timestamp 1624635492
transform 1 0 17480 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__B
timestamp 1624635492
transform -1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1624635492
transform 1 0 18124 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 18952 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1624635492
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1624635492
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1624635492
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1624635492
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1624635492
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1624635492
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1624635492
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_190
timestamp 1624635492
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_184
timestamp 1624635492
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_188
timestamp 1624635492
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_180
timestamp 1624635492
transform 1 0 17664 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 18952 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 18952 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_146
timestamp 1624635492
transform 1 0 14536 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1624635492
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1624635492
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1624635492
transform 1 0 16744 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_158
timestamp 1624635492
transform 1 0 15640 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1624635492
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_175
timestamp 1624635492
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1624635492
transform 1 0 17112 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_204
timestamp 1624635492
transform 1 0 19872 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_199
timestamp 1624635492
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1624635492
transform 1 0 19780 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_216
timestamp 1624635492
transform 1 0 20976 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1624635492
transform 1 0 22540 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1624635492
transform 1 0 22080 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1624635492
transform 1 0 22448 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_257
timestamp 1624635492
transform 1 0 24748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_245
timestamp 1624635492
transform 1 0 23644 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1624635492
transform 1 0 25116 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_262
timestamp 1624635492
transform 1 0 25208 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1624635492
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1624635492
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1624635492
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1624635492
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1624635492
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1624635492
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1624635492
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1624635492
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1624635492
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1624635492
transform 1 0 23276 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_229
timestamp 1624635492
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1624635492
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1624635492
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1624635492
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1624635492
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1624635492
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1624635492
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_156
timestamp 1624635492
transform 1 0 15456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1624635492
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1624635492
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_192
timestamp 1624635492
transform 1 0 18768 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1624635492
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_225
timestamp 1624635492
transform 1 0 21804 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_213
timestamp 1624635492
transform 1 0 20700 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1624635492
transform 1 0 22908 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1624635492
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_249
timestamp 1624635492
transform 1 0 24012 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1624635492
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1624635492
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_143
timestamp 1624635492
transform 1 0 14260 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1624635492
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_167
timestamp 1624635492
transform 1 0 16468 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_155
timestamp 1624635492
transform 1 0 15364 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1624635492
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1624635492
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1624635492
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_220
timestamp 1624635492
transform 1 0 21344 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1624635492
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1624635492
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1624635492
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1624635492
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1624635492
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_265
timestamp 1624635492
transform 1 0 25484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_144
timestamp 1624635492
transform 1 0 14352 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1624635492
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _191_
timestamp 1624635492
transform 1 0 15088 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_167
timestamp 1624635492
transform 1 0 16468 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_155
timestamp 1624635492
transform 1 0 15364 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_179
timestamp 1624635492
transform 1 0 17572 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1624635492
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_199
timestamp 1624635492
transform 1 0 19412 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_191
timestamp 1624635492
transform 1 0 18676 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1624635492
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1624635492
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1624635492
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1624635492
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1624635492
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1624635492
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1624635492
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_270
timestamp 1624635492
transform 1 0 25944 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_144
timestamp 1624635492
transform 1 0 14352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_140
timestamp 1624635492
transform 1 0 13984 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_144
timestamp 1624635492
transform 1 0 14352 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1624635492
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1624635492
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1624635492
transform 1 0 15456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1624635492
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_168
timestamp 1624635492
transform 1 0 16560 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_156
timestamp 1624635492
transform 1 0 15456 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1624635492
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1624635492
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1624635492
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1624635492
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_192
timestamp 1624635492
transform 1 0 18768 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1624635492
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1624635492
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_225
timestamp 1624635492
transform 1 0 21804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1624635492
transform 1 0 20700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_220
timestamp 1624635492
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1624635492
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1624635492
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1624635492
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1624635492
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1624635492
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1624635492
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_249
timestamp 1624635492
transform 1 0 24012 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1624635492
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1624635492
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_270
timestamp 1624635492
transform 1 0 25944 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_265
timestamp 1624635492
transform 1 0 25484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_151
timestamp 1624635492
transform 1 0 14996 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_139
timestamp 1624635492
transform 1 0 13892 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1624635492
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_163
timestamp 1624635492
transform 1 0 16100 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1624635492
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1624635492
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1624635492
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1624635492
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1624635492
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1624635492
transform 1 0 23276 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_229
timestamp 1624635492
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1624635492
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1624635492
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1624635492
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1624635492
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1624635492
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_168
timestamp 1624635492
transform 1 0 16560 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1624635492
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1624635492
transform 1 0 17664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1624635492
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_192
timestamp 1624635492
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1624635492
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_213
timestamp 1624635492
transform 1 0 20700 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  _049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 23000 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_238
timestamp 1624635492
transform 1 0 23000 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__049__A
timestamp 1624635492
transform -1 0 23552 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1624635492
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_256
timestamp 1624635492
transform 1 0 24656 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_244
timestamp 1624635492
transform 1 0 23552 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1624635492
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1624635492
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1624635492
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1624635492
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1624635492
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_163
timestamp 1624635492
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1624635492
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1624635492
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1624635492
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1624635492
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1624635492
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1624635492
transform 1 0 23276 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1624635492
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1624635492
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1624635492
transform 1 0 24380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_265
timestamp 1624635492
transform 1 0 25484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1624635492
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1624635492
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1624635492
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1624635492
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1624635492
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1624635492
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_192
timestamp 1624635492
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1624635492
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1624635492
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1624635492
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1624635492
transform 1 0 22908 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1624635492
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_249
timestamp 1624635492
transform 1 0 24012 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1624635492
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1624635492
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_144
timestamp 1624635492
transform 1 0 14352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_151
timestamp 1624635492
transform 1 0 14996 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_139
timestamp 1624635492
transform 1 0 13892 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1624635492
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_168
timestamp 1624635492
transform 1 0 16560 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_156
timestamp 1624635492
transform 1 0 15456 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_172
timestamp 1624635492
transform 1 0 16928 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_163
timestamp 1624635492
transform 1 0 16100 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1624635492
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_180
timestamp 1624635492
transform 1 0 17664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1624635492
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1624635492
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_192
timestamp 1624635492
transform 1 0 18768 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1624635492
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1624635492
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_225
timestamp 1624635492
transform 1 0 21804 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_213
timestamp 1624635492
transform 1 0 20700 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_220
timestamp 1624635492
transform 1 0 21344 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1624635492
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_237
timestamp 1624635492
transform 1 0 22908 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1624635492
transform 1 0 23276 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_229
timestamp 1624635492
transform 1 0 22172 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1624635492
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1624635492
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_256
timestamp 1624635492
transform 1 0 24656 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_252
timestamp 1624635492
transform 1 0 24288 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1624635492
transform 1 0 24380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1624635492
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _265_
timestamp 1624635492
transform 1 0 24012 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1624635492
transform 1 0 25944 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_265
timestamp 1624635492
transform 1 0 25484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1624635492
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1624635492
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1624635492
transform 1 0 16928 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_163
timestamp 1624635492
transform 1 0 16100 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1624635492
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_187
timestamp 1624635492
transform 1 0 18308 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_184
timestamp 1624635492
transform 1 0 18032 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__D
timestamp 1624635492
transform -1 0 18308 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1624635492
transform 1 0 19964 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1624635492
transform 1 0 18860 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__CLK
timestamp 1624635492
transform 1 0 18676 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1624635492
transform 1 0 21804 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_217
timestamp 1624635492
transform 1 0 21068 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1624635492
transform 1 0 23276 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_229
timestamp 1624635492
transform 1 0 22172 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1624635492
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1624635492
transform 1 0 24380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1624635492
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_144
timestamp 1624635492
transform 1 0 14352 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1624635492
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_156
timestamp 1624635492
transform 1 0 15456 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _336_
timestamp 1624635492
transform -1 0 18124 0 -1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1624635492
transform 1 0 18124 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _171_
timestamp 1624635492
transform -1 0 18768 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_201
timestamp 1624635492
transform 1 0 19596 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_192
timestamp 1624635492
transform 1 0 18768 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1624635492
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1624635492
transform 1 0 21804 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1624635492
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1624635492
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1624635492
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_249
timestamp 1624635492
transform 1 0 24012 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1624635492
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1624635492
transform 1 0 25944 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1624635492
transform 1 0 14628 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_172
timestamp 1624635492
transform 1 0 16928 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_159
timestamp 1624635492
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1624635492
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_183
timestamp 1624635492
transform 1 0 17940 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _222_
timestamp 1624635492
transform 1 0 18492 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _164_
timestamp 1624635492
transform -1 0 17940 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_204
timestamp 1624635492
transform 1 0 19872 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_192
timestamp 1624635492
transform 1 0 18768 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_216
timestamp 1624635492
transform 1 0 20976 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_241
timestamp 1624635492
transform 1 0 23276 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_229
timestamp 1624635492
transform 1 0 22172 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1624635492
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1624635492
transform 1 0 24380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_265
timestamp 1624635492
transform 1 0 25484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_144
timestamp 1624635492
transform 1 0 14352 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1624635492
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_168
timestamp 1624635492
transform 1 0 16560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_156
timestamp 1624635492
transform 1 0 15456 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_180
timestamp 1624635492
transform 1 0 17664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_201
timestamp 1624635492
transform 1 0 19596 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_192
timestamp 1624635492
transform 1 0 18768 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1624635492
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_225
timestamp 1624635492
transform 1 0 21804 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_213
timestamp 1624635492
transform 1 0 20700 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_237
timestamp 1624635492
transform 1 0 22908 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_258
timestamp 1624635492
transform 1 0 24840 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_249
timestamp 1624635492
transform 1 0 24012 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1624635492
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_270
timestamp 1624635492
transform 1 0 25944 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_151
timestamp 1624635492
transform 1 0 14996 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_139
timestamp 1624635492
transform 1 0 13892 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1624635492
transform 1 0 16928 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_163
timestamp 1624635492
transform 1 0 16100 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1624635492
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1624635492
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1624635492
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_220
timestamp 1624635492
transform 1 0 21344 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1624635492
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_241
timestamp 1624635492
transform 1 0 23276 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1624635492
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1624635492
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1624635492
transform 1 0 24380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1624635492
transform 1 0 25484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_146
timestamp 1624635492
transform 1 0 14536 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_144
timestamp 1624635492
transform 1 0 14352 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1624635492
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_172
timestamp 1624635492
transform 1 0 16928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_170
timestamp 1624635492
transform 1 0 16744 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_158
timestamp 1624635492
transform 1 0 15640 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_168
timestamp 1624635492
transform 1 0 16560 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_156
timestamp 1624635492
transform 1 0 15456 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1624635492
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1624635492
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1624635492
transform 1 0 17664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1624635492
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_201
timestamp 1624635492
transform 1 0 19596 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_192
timestamp 1624635492
transform 1 0 18768 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1624635492
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_220
timestamp 1624635492
transform 1 0 21344 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1624635492
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_217
timestamp 1624635492
transform 1 0 21068 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1624635492
transform 1 0 20700 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _276_
timestamp 1624635492
transform 1 0 20792 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_241
timestamp 1624635492
transform 1 0 23276 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_229
timestamp 1624635492
transform 1 0 22172 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_241
timestamp 1624635492
transform 1 0 23276 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_229
timestamp 1624635492
transform 1 0 22172 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1624635492
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_253
timestamp 1624635492
transform 1 0 24380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_258
timestamp 1624635492
transform 1 0 24840 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1624635492
transform 1 0 24380 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1624635492
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1624635492
transform 1 0 25484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_270
timestamp 1624635492
transform 1 0 25944 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_144
timestamp 1624635492
transform 1 0 14352 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1624635492
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_168
timestamp 1624635492
transform 1 0 16560 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_156
timestamp 1624635492
transform 1 0 15456 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1624635492
transform 1 0 17664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_201
timestamp 1624635492
transform 1 0 19596 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_192
timestamp 1624635492
transform 1 0 18768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1624635492
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_225
timestamp 1624635492
transform 1 0 21804 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_213
timestamp 1624635492
transform 1 0 20700 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_237
timestamp 1624635492
transform 1 0 22908 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1624635492
transform 1 0 24840 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_249
timestamp 1624635492
transform 1 0 24012 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1624635492
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_271
timestamp 1624635492
transform 1 0 26036 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_265
timestamp 1624635492
transform 1 0 25484 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_wb_clk_i_A
timestamp 1624635492
transform -1 0 26036 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 25208 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_400
timestamp 1624635492
transform 1 0 37904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_294
timestamp 1624635492
transform 1 0 37628 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_400
timestamp 1624635492
transform 1 0 37904 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_296
timestamp 1624635492
transform 1 0 37628 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_400
timestamp 1624635492
transform 1 0 37904 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_298
timestamp 1624635492
transform 1 0 37628 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_400
timestamp 1624635492
transform 1 0 37904 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_400
timestamp 1624635492
transform 1 0 37904 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_302
timestamp 1624635492
transform 1 0 37628 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_300
timestamp 1624635492
transform 1 0 37628 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_291
timestamp 1624635492
transform 1 0 27876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1624635492
transform 1 0 27416 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_282
timestamp 1624635492
transform 1 0 27048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_274
timestamp 1624635492
transform 1 0 26312 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A1
timestamp 1624635492
transform -1 0 27416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1624635492
transform 1 0 27784 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1624635492
transform 1 0 29532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_296
timestamp 1624635492
transform 1 0 28336 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A2
timestamp 1624635492
transform 1 0 28152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_2  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 28704 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_325
timestamp 1624635492
transform 1 0 31004 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_320
timestamp 1624635492
transform 1 0 30544 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_315
timestamp 1624635492
transform 1 0 30084 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B1
timestamp 1624635492
transform -1 0 30084 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1624635492
transform -1 0 31004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1624635492
transform 1 0 30452 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 31924 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_349
timestamp 1624635492
transform 1 0 33212 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_347
timestamp 1624635492
transform 1 0 33028 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_335
timestamp 1624635492
transform 1 0 31924 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1624635492
transform 1 0 33120 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_372
timestamp 1624635492
transform 1 0 35328 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_360
timestamp 1624635492
transform 1 0 34224 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _167_
timestamp 1624635492
transform -1 0 34224 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_390
timestamp 1624635492
transform 1 0 36984 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_378
timestamp 1624635492
transform 1 0 35880 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_376
timestamp 1624635492
transform 1 0 35696 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1624635492
transform 1 0 35788 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_407
timestamp 1624635492
transform 1 0 38548 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1624635492
transform 1 0 38088 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1624635492
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1624635492
transform 1 0 27968 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_286
timestamp 1624635492
transform 1 0 27416 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_277
timestamp 1624635492
transform 1 0 26588 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__C1
timestamp 1624635492
transform 1 0 27784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1624635492
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_309
timestamp 1624635492
transform 1 0 29532 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_298
timestamp 1624635492
transform 1 0 28520 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A3
timestamp 1624635492
transform 1 0 28336 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _187_
timestamp 1624635492
transform -1 0 29532 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_330
timestamp 1624635492
transform 1 0 31464 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_318
timestamp 1624635492
transform 1 0 30360 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _289_
timestamp 1624635492
transform 1 0 30084 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1624635492
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1624635492
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1624635492
transform 1 0 34868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1624635492
transform 1 0 33764 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_391
timestamp 1624635492
transform 1 0 37076 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1624635492
transform 1 0 35972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_400
timestamp 1624635492
transform 1 0 37904 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1624635492
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_282
timestamp 1624635492
transform 1 0 27048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_306
timestamp 1624635492
transform 1 0 29256 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_294
timestamp 1624635492
transform 1 0 28152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_327
timestamp 1624635492
transform 1 0 31188 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_315
timestamp 1624635492
transform 1 0 30084 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1624635492
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_349
timestamp 1624635492
transform 1 0 33212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_345
timestamp 1624635492
transform 1 0 32844 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_339
timestamp 1624635492
transform 1 0 32292 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _253_
timestamp 1624635492
transform 1 0 32936 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_372
timestamp 1624635492
transform 1 0 35328 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_369
timestamp 1624635492
transform 1 0 35052 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_361
timestamp 1624635492
transform 1 0 34316 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1624635492
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_390
timestamp 1624635492
transform 1 0 36984 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_384
timestamp 1624635492
transform 1 0 36432 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _214_
timestamp 1624635492
transform 1 0 37076 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_406
timestamp 1624635492
transform 1 0 38456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_394
timestamp 1624635492
transform 1 0 37352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1624635492
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1624635492
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1624635492
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_310
timestamp 1624635492
transform 1 0 29624 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_298
timestamp 1624635492
transform 1 0 28520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_331
timestamp 1624635492
transform 1 0 31556 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_322
timestamp 1624635492
transform 1 0 30728 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _240_
timestamp 1624635492
transform 1 0 31280 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_343
timestamp 1624635492
transform 1 0 32660 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_339
timestamp 1624635492
transform 1 0 32292 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1624635492
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _205_
timestamp 1624635492
transform 1 0 33396 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_366
timestamp 1624635492
transform 1 0 34776 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_354
timestamp 1624635492
transform 1 0 33672 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_381
timestamp 1624635492
transform 1 0 36156 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _203_
timestamp 1624635492
transform 1 0 35880 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_400
timestamp 1624635492
transform 1 0 37904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_393
timestamp 1624635492
transform 1 0 37260 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1624635492
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_282
timestamp 1624635492
transform 1 0 27048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_306
timestamp 1624635492
transform 1 0 29256 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_294
timestamp 1624635492
transform 1 0 28152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_329
timestamp 1624635492
transform 1 0 31372 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_317
timestamp 1624635492
transform 1 0 30268 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A1
timestamp 1624635492
transform -1 0 30268 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1624635492
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_341
timestamp 1624635492
transform 1 0 32476 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_372
timestamp 1624635492
transform 1 0 35328 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_365
timestamp 1624635492
transform 1 0 34684 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_353
timestamp 1624635492
transform 1 0 33580 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1624635492
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_384
timestamp 1624635492
transform 1 0 36432 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_404
timestamp 1624635492
transform 1 0 38272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_396
timestamp 1624635492
transform 1 0 37536 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__D
timestamp 1624635492
transform -1 0 38272 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_282
timestamp 1624635492
transform 1 0 27048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1624635492
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_277
timestamp 1624635492
transform 1 0 26588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1624635492
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_306
timestamp 1624635492
transform 1 0 29256 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_294
timestamp 1624635492
transform 1 0 28152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_310
timestamp 1624635492
transform 1 0 29624 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1624635492
transform 1 0 28520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__B1
timestamp 1624635492
transform 1 0 29808 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_327
timestamp 1624635492
transform 1 0 31188 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_315
timestamp 1624635492
transform 1 0 30084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1624635492
transform 1 0 31648 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1624635492
transform 1 0 31096 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_314
timestamp 1624635492
transform 1 0 29992 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A2
timestamp 1624635492
transform 1 0 31464 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1624635492
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 31096 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1624635492
transform 1 0 33396 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1624635492
transform 1 0 32292 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_343
timestamp 1624635492
transform 1 0 32660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_338
timestamp 1624635492
transform 1 0 32200 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__B2
timestamp 1624635492
transform 1 0 32016 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1624635492
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_372
timestamp 1624635492
transform 1 0 35328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_363
timestamp 1624635492
transform 1 0 34500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1624635492
transform 1 0 34868 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_355
timestamp 1624635492
transform 1 0 33764 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1624635492
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_384
timestamp 1624635492
transform 1 0 36432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_391
timestamp 1624635492
transform 1 0 37076 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_379
timestamp 1624635492
transform 1 0 35972 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_402
timestamp 1624635492
transform 1 0 38088 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_396
timestamp 1624635492
transform 1 0 37536 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_400
timestamp 1624635492
transform 1 0 37904 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__CLK
timestamp 1624635492
transform 1 0 37904 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1624635492
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _348_
timestamp 1624635492
transform 1 0 38272 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_39_286
timestamp 1624635492
transform 1 0 27416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_277
timestamp 1624635492
transform 1 0 26588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1624635492
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_310
timestamp 1624635492
transform 1 0 29624 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_298
timestamp 1624635492
transform 1 0 28520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_322
timestamp 1624635492
transform 1 0 30728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1624635492
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_334
timestamp 1624635492
transform 1 0 31832 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1624635492
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1624635492
transform 1 0 34868 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1624635492
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_391
timestamp 1624635492
transform 1 0 37076 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1624635492
transform 1 0 35972 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_400
timestamp 1624635492
transform 1 0 37904 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1624635492
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1624635492
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_305
timestamp 1624635492
transform 1 0 29164 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_294
timestamp 1624635492
transform 1 0 28152 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _287_
timestamp 1624635492
transform 1 0 28888 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1624635492
transform 1 0 31188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1624635492
transform 1 0 30084 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1624635492
transform 1 0 29900 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1624635492
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_351
timestamp 1624635492
transform 1 0 33396 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1624635492
transform 1 0 32292 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _120_
timestamp 1624635492
transform 1 0 33488 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_372
timestamp 1624635492
transform 1 0 35328 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_367
timestamp 1624635492
transform 1 0 34868 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_355
timestamp 1624635492
transform 1 0 33764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1624635492
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_384
timestamp 1624635492
transform 1 0 36432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_408
timestamp 1624635492
transform 1 0 38640 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_396
timestamp 1624635492
transform 1 0 37536 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1624635492
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_277
timestamp 1624635492
transform 1 0 26588 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1624635492
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_310
timestamp 1624635492
transform 1 0 29624 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_298
timestamp 1624635492
transform 1 0 28520 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_322
timestamp 1624635492
transform 1 0 30728 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1624635492
transform 1 0 32660 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_334
timestamp 1624635492
transform 1 0 31832 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1624635492
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1624635492
transform 1 0 34868 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_355
timestamp 1624635492
transform 1 0 33764 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_392
timestamp 1624635492
transform 1 0 37168 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_387
timestamp 1624635492
transform 1 0 36708 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_379
timestamp 1624635492
transform 1 0 35972 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _174_
timestamp 1624635492
transform -1 0 37168 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_400
timestamp 1624635492
transform 1 0 37904 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_398
timestamp 1624635492
transform 1 0 37720 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1624635492
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1624635492
transform 1 0 27048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_306
timestamp 1624635492
transform 1 0 29256 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1624635492
transform 1 0 28152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_327
timestamp 1624635492
transform 1 0 31188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_315
timestamp 1624635492
transform 1 0 30084 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1624635492
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1624635492
transform 1 0 33396 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1624635492
transform 1 0 32292 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_372
timestamp 1624635492
transform 1 0 35328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_363
timestamp 1624635492
transform 1 0 34500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1624635492
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_384
timestamp 1624635492
transform 1 0 36432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_408
timestamp 1624635492
transform 1 0 38640 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_396
timestamp 1624635492
transform 1 0 37536 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _258_
timestamp 1624635492
transform 1 0 27140 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_277
timestamp 1624635492
transform 1 0 26588 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_282
timestamp 1624635492
transform 1 0 27048 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1624635492
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A2
timestamp 1624635492
transform -1 0 27876 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_286
timestamp 1624635492
transform 1 0 27416 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_286
timestamp 1624635492
transform 1 0 27416 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_290
timestamp 1624635492
transform 1 0 27784 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 29072 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_43_291
timestamp 1624635492
transform 1 0 27876 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_310
timestamp 1624635492
transform 1 0 29624 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1624635492
transform 1 0 29072 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_303
timestamp 1624635492
transform 1 0 28980 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A1
timestamp 1624635492
transform 1 0 29440 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_329
timestamp 1624635492
transform 1 0 31372 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_317
timestamp 1624635492
transform 1 0 30268 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_327
timestamp 1624635492
transform 1 0 31188 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_315
timestamp 1624635492
transform 1 0 30084 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__B1
timestamp 1624635492
transform 1 0 30084 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1624635492
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_341
timestamp 1624635492
transform 1 0 32476 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_343
timestamp 1624635492
transform 1 0 32660 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_339
timestamp 1624635492
transform 1 0 32292 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1624635492
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_372
timestamp 1624635492
transform 1 0 35328 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_365
timestamp 1624635492
transform 1 0 34684 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_353
timestamp 1624635492
transform 1 0 33580 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1624635492
transform 1 0 34868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_355
timestamp 1624635492
transform 1 0 33764 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1624635492
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_384
timestamp 1624635492
transform 1 0 36432 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_391
timestamp 1624635492
transform 1 0 37076 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1624635492
transform 1 0 35972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_404
timestamp 1624635492
transform 1 0 38272 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_400
timestamp 1624635492
transform 1 0 37904 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_396
timestamp 1624635492
transform 1 0 37536 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_400
timestamp 1624635492
transform 1 0 37904 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1624635492
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _163_
timestamp 1624635492
transform -1 0 38272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_286
timestamp 1624635492
transform 1 0 27416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1624635492
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1624635492
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_310
timestamp 1624635492
transform 1 0 29624 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1624635492
transform 1 0 28520 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_330
timestamp 1624635492
transform 1 0 31464 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_326
timestamp 1624635492
transform 1 0 31096 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_322
timestamp 1624635492
transform 1 0 30728 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _144_
timestamp 1624635492
transform 1 0 31188 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_343
timestamp 1624635492
transform 1 0 32660 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1624635492
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1624635492
transform 1 0 34868 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_355
timestamp 1624635492
transform 1 0 33764 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_391
timestamp 1624635492
transform 1 0 37076 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1624635492
transform 1 0 35972 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_400
timestamp 1624635492
transform 1 0 37904 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1624635492
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1624635492
transform 1 0 27048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_306
timestamp 1624635492
transform 1 0 29256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_294
timestamp 1624635492
transform 1 0 28152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_328
timestamp 1624635492
transform 1 0 31280 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_323
timestamp 1624635492
transform 1 0 30820 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_315
timestamp 1624635492
transform 1 0 30084 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A3
timestamp 1624635492
transform 1 0 31096 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1624635492
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_352
timestamp 1624635492
transform 1 0 33488 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_340
timestamp 1624635492
transform 1 0 32384 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_372
timestamp 1624635492
transform 1 0 35328 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_370
timestamp 1624635492
transform 1 0 35144 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_364
timestamp 1624635492
transform 1 0 34592 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1624635492
transform 1 0 35236 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_384
timestamp 1624635492
transform 1 0 36432 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_408
timestamp 1624635492
transform 1 0 38640 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_396
timestamp 1624635492
transform 1 0 37536 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1624635492
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1624635492
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1624635492
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_310
timestamp 1624635492
transform 1 0 29624 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_298
timestamp 1624635492
transform 1 0 28520 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_326
timestamp 1624635492
transform 1 0 31096 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_322
timestamp 1624635492
transform 1 0 30728 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A2
timestamp 1624635492
transform 1 0 30912 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_1  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 31464 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_351
timestamp 1624635492
transform 1 0 33396 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_345
timestamp 1624635492
transform 1 0 32844 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_338
timestamp 1624635492
transform 1 0 32200 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__C1
timestamp 1624635492
transform -1 0 33396 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B1
timestamp 1624635492
transform 1 0 32660 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1624635492
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_363
timestamp 1624635492
transform 1 0 34500 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_392
timestamp 1624635492
transform 1 0 37168 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_380
timestamp 1624635492
transform 1 0 36064 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_375
timestamp 1624635492
transform 1 0 35604 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _312_
timestamp 1624635492
transform -1 0 36064 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_400
timestamp 1624635492
transform 1 0 37904 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_398
timestamp 1624635492
transform 1 0 37720 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1624635492
transform 1 0 37812 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_282
timestamp 1624635492
transform 1 0 27048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_306
timestamp 1624635492
transform 1 0 29256 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_294
timestamp 1624635492
transform 1 0 28152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_326
timestamp 1624635492
transform 1 0 31096 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_323
timestamp 1624635492
transform 1 0 30820 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_315
timestamp 1624635492
transform 1 0 30084 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A1
timestamp 1624635492
transform 1 0 30912 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1624635492
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_350
timestamp 1624635492
transform 1 0 33304 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_338
timestamp 1624635492
transform 1 0 32200 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1624635492
transform 1 0 35328 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_370
timestamp 1624635492
transform 1 0 35144 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_362
timestamp 1624635492
transform 1 0 34408 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1624635492
transform 1 0 35236 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_384
timestamp 1624635492
transform 1 0 36432 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_408
timestamp 1624635492
transform 1 0 38640 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_396
timestamp 1624635492
transform 1 0 37536 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_290
timestamp 1624635492
transform 1 0 27784 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1624635492
transform 1 0 27416 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_277
timestamp 1624635492
transform 1 0 26588 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B1
timestamp 1624635492
transform 1 0 27876 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1624635492
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_307
timestamp 1624635492
transform 1 0 29348 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_301
timestamp 1624635492
transform 1 0 28796 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_293
timestamp 1624635492
transform 1 0 28060 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _301_
timestamp 1624635492
transform -1 0 29348 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_331
timestamp 1624635492
transform 1 0 31556 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_319
timestamp 1624635492
transform 1 0 30452 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_343
timestamp 1624635492
transform 1 0 32660 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_339
timestamp 1624635492
transform 1 0 32292 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1624635492
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1624635492
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_355
timestamp 1624635492
transform 1 0 33764 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_391
timestamp 1624635492
transform 1 0 37076 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1624635492
transform 1 0 35972 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_400
timestamp 1624635492
transform 1 0 37904 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1624635492
transform 1 0 37812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_286
timestamp 1624635492
transform 1 0 27416 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_277
timestamp 1624635492
transform 1 0 26588 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_287
timestamp 1624635492
transform 1 0 27508 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_276
timestamp 1624635492
transform 1 0 26496 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A3
timestamp 1624635492
transform 1 0 26312 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A1
timestamp 1624635492
transform 1 0 27876 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1624635492
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _184_
timestamp 1624635492
transform -1 0 28060 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _074_
timestamp 1624635492
transform -1 0 27508 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1624635492
transform 1 0 29164 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1624635492
transform 1 0 28060 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_311
timestamp 1624635492
transform 1 0 29716 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_299
timestamp 1624635492
transform 1 0 28612 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_293
timestamp 1624635492
transform 1 0 28060 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A2
timestamp 1624635492
transform 1 0 28428 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_329
timestamp 1624635492
transform 1 0 31372 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1624635492
transform 1 0 30268 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_327
timestamp 1624635492
transform 1 0 31188 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_315
timestamp 1624635492
transform 1 0 30084 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1624635492
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1624635492
transform 1 0 32660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_341
timestamp 1624635492
transform 1 0 32476 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1624635492
transform 1 0 33396 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1624635492
transform 1 0 32292 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1624635492
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1624635492
transform 1 0 34868 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1624635492
transform 1 0 33764 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_372
timestamp 1624635492
transform 1 0 35328 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_363
timestamp 1624635492
transform 1 0 34500 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1624635492
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1624635492
transform 1 0 35972 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_391
timestamp 1624635492
transform 1 0 37076 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_379
timestamp 1624635492
transform 1 0 35972 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A1
timestamp 1624635492
transform 1 0 37076 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _118_
timestamp 1624635492
transform 1 0 35696 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_408
timestamp 1624635492
transform 1 0 38640 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_400
timestamp 1624635492
transform 1 0 37904 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_393
timestamp 1624635492
transform 1 0 37260 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_403
timestamp 1624635492
transform 1 0 38180 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1624635492
transform 1 0 37812 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_283
timestamp 1624635492
transform 1 0 27140 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_307
timestamp 1624635492
transform 1 0 29348 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_295
timestamp 1624635492
transform 1 0 28244 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_327
timestamp 1624635492
transform 1 0 31188 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1624635492
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_313
timestamp 1624635492
transform 1 0 29900 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1624635492
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_351
timestamp 1624635492
transform 1 0 33396 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_339
timestamp 1624635492
transform 1 0 32292 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1624635492
transform 1 0 35328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_363
timestamp 1624635492
transform 1 0 34500 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1624635492
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_391
timestamp 1624635492
transform 1 0 37076 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_388
timestamp 1624635492
transform 1 0 36800 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_384
timestamp 1624635492
transform 1 0 36432 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__B1
timestamp 1624635492
transform 1 0 36892 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_409
timestamp 1624635492
transform 1 0 38732 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1624635492
transform 1 0 38180 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A2
timestamp 1624635492
transform 1 0 38548 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _057_
timestamp 1624635492
transform -1 0 38180 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_424
timestamp 1624635492
transform 1 0 40112 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_412
timestamp 1624635492
transform 1 0 39008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_436
timestamp 1624635492
transform 1 0 41216 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_455
timestamp 1624635492
transform 1 0 42964 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_448
timestamp 1624635492
transform 1 0 42320 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1682
timestamp 1624635492
transform 1 0 42872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_479
timestamp 1624635492
transform 1 0 45172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_467
timestamp 1624635492
transform 1 0 44068 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_491
timestamp 1624635492
transform 1 0 46276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_512
timestamp 1624635492
transform 1 0 48208 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_503
timestamp 1624635492
transform 1 0 47380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1683
timestamp 1624635492
transform 1 0 48116 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_524
timestamp 1624635492
transform 1 0 49312 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_536
timestamp 1624635492
transform 1 0 50416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_427
timestamp 1624635492
transform 1 0 40388 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_424
timestamp 1624635492
transform 1 0 40112 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_412
timestamp 1624635492
transform 1 0 39008 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1687
timestamp 1624635492
transform 1 0 40296 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_439
timestamp 1624635492
transform 1 0 41492 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_463
timestamp 1624635492
transform 1 0 43700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_451
timestamp 1624635492
transform 1 0 42596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_475
timestamp 1624635492
transform 1 0 44804 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_496
timestamp 1624635492
transform 1 0 46736 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_484
timestamp 1624635492
transform 1 0 45632 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1688
timestamp 1624635492
transform 1 0 45540 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_507
timestamp 1624635492
transform 1 0 47748 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _262_
timestamp 1624635492
transform 1 0 47472 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_531
timestamp 1624635492
transform 1 0 49956 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_519
timestamp 1624635492
transform 1 0 48852 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_541
timestamp 1624635492
transform 1 0 50876 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_539
timestamp 1624635492
transform 1 0 50692 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1689
timestamp 1624635492
transform 1 0 50784 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_424
timestamp 1624635492
transform 1 0 40112 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_412
timestamp 1624635492
transform 1 0 39008 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_436
timestamp 1624635492
transform 1 0 41216 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_455
timestamp 1624635492
transform 1 0 42964 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_448
timestamp 1624635492
transform 1 0 42320 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1693
timestamp 1624635492
transform 1 0 42872 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_479
timestamp 1624635492
transform 1 0 45172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_467
timestamp 1624635492
transform 1 0 44068 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_491
timestamp 1624635492
transform 1 0 46276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_512
timestamp 1624635492
transform 1 0 48208 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_503
timestamp 1624635492
transform 1 0 47380 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1694
timestamp 1624635492
transform 1 0 48116 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_524
timestamp 1624635492
transform 1 0 49312 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_536
timestamp 1624635492
transform 1 0 50416 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_424
timestamp 1624635492
transform 1 0 40112 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_412
timestamp 1624635492
transform 1 0 39008 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_427
timestamp 1624635492
transform 1 0 40388 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_424
timestamp 1624635492
transform 1 0 40112 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_412
timestamp 1624635492
transform 1 0 39008 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1698
timestamp 1624635492
transform 1 0 40296 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_436
timestamp 1624635492
transform 1 0 41216 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_439
timestamp 1624635492
transform 1 0 41492 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_455
timestamp 1624635492
transform 1 0 42964 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_448
timestamp 1624635492
transform 1 0 42320 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_463
timestamp 1624635492
transform 1 0 43700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_451
timestamp 1624635492
transform 1 0 42596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1704
timestamp 1624635492
transform 1 0 42872 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_479
timestamp 1624635492
transform 1 0 45172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_467
timestamp 1624635492
transform 1 0 44068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_475
timestamp 1624635492
transform 1 0 44804 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_491
timestamp 1624635492
transform 1 0 46276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_496
timestamp 1624635492
transform 1 0 46736 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_484
timestamp 1624635492
transform 1 0 45632 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1699
timestamp 1624635492
transform 1 0 45540 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_512
timestamp 1624635492
transform 1 0 48208 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_503
timestamp 1624635492
transform 1 0 47380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_508
timestamp 1624635492
transform 1 0 47840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1705
timestamp 1624635492
transform 1 0 48116 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1624635492
transform 1 0 49772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_524
timestamp 1624635492
transform 1 0 49312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_532
timestamp 1624635492
transform 1 0 50048 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_520
timestamp 1624635492
transform 1 0 48944 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _272_
timestamp 1624635492
transform 1 0 49496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1624635492
transform 1 0 50876 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_541
timestamp 1624635492
transform 1 0 50876 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1700
timestamp 1624635492
transform 1 0 50784 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _156_
timestamp 1624635492
transform -1 0 51520 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_419
timestamp 1624635492
transform 1 0 39652 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_436
timestamp 1624635492
transform 1 0 41216 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_431
timestamp 1624635492
transform 1 0 40756 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1624635492
transform 1 0 41124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_460
timestamp 1624635492
transform 1 0 43424 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_448
timestamp 1624635492
transform 1 0 42320 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1624635492
transform 1 0 44988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_465
timestamp 1624635492
transform 1 0 43884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1624635492
transform 1 0 43792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_494
timestamp 1624635492
transform 1 0 46552 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_489
timestamp 1624635492
transform 1 0 46092 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1624635492
transform 1 0 46460 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_506
timestamp 1624635492
transform 1 0 47656 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_523
timestamp 1624635492
transform 1 0 49220 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_518
timestamp 1624635492
transform 1 0 48760 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1624635492
transform 1 0 49128 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_539
timestamp 1624635492
transform 1 0 50692 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_535
timestamp 1624635492
transform 1 0 50324 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _226_
timestamp 1624635492
transform -1 0 50692 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_424
timestamp 1624635492
transform 1 0 40112 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_412
timestamp 1624635492
transform 1 0 39008 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_436
timestamp 1624635492
transform 1 0 41216 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_457
timestamp 1624635492
transform 1 0 43148 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_448
timestamp 1624635492
transform 1 0 42320 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1624635492
transform 1 0 43056 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_481
timestamp 1624635492
transform 1 0 45356 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_469
timestamp 1624635492
transform 1 0 44252 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_493
timestamp 1624635492
transform 1 0 46460 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_514
timestamp 1624635492
transform 1 0 48392 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1624635492
transform 1 0 47564 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1624635492
transform 1 0 48300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_526
timestamp 1624635492
transform 1 0 49496 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_538
timestamp 1624635492
transform 1 0 50600 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_426
timestamp 1624635492
transform 1 0 40296 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_418
timestamp 1624635492
transform 1 0 39560 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_441
timestamp 1624635492
transform 1 0 41676 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_429
timestamp 1624635492
transform 1 0 40572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1624635492
transform 1 0 40480 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_453
timestamp 1624635492
transform 1 0 42780 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_477
timestamp 1624635492
transform 1 0 44988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_465
timestamp 1624635492
transform 1 0 43884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_498
timestamp 1624635492
transform 1 0 46920 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_486
timestamp 1624635492
transform 1 0 45816 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1624635492
transform 1 0 45724 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_510
timestamp 1624635492
transform 1 0 48024 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_534
timestamp 1624635492
transform 1 0 50232 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_522
timestamp 1624635492
transform 1 0 49128 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_543
timestamp 1624635492
transform 1 0 51060 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1624635492
transform 1 0 50968 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_424
timestamp 1624635492
transform 1 0 40112 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_412
timestamp 1624635492
transform 1 0 39008 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_436
timestamp 1624635492
transform 1 0 41216 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_457
timestamp 1624635492
transform 1 0 43148 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_448
timestamp 1624635492
transform 1 0 42320 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1624635492
transform 1 0 43056 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_481
timestamp 1624635492
transform 1 0 45356 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_469
timestamp 1624635492
transform 1 0 44252 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_493
timestamp 1624635492
transform 1 0 46460 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_514
timestamp 1624635492
transform 1 0 48392 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1624635492
transform 1 0 47564 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1624635492
transform 1 0 48300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_526
timestamp 1624635492
transform 1 0 49496 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_538
timestamp 1624635492
transform 1 0 50600 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_416
timestamp 1624635492
transform 1 0 39376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_441
timestamp 1624635492
transform 1 0 41676 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_429
timestamp 1624635492
transform 1 0 40572 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1624635492
transform 1 0 40480 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_453
timestamp 1624635492
transform 1 0 42780 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_477
timestamp 1624635492
transform 1 0 44988 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_465
timestamp 1624635492
transform 1 0 43884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_498
timestamp 1624635492
transform 1 0 46920 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_486
timestamp 1624635492
transform 1 0 45816 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1624635492
transform 1 0 45724 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_510
timestamp 1624635492
transform 1 0 48024 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_534
timestamp 1624635492
transform 1 0 50232 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_522
timestamp 1624635492
transform 1 0 49128 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_543
timestamp 1624635492
transform 1 0 51060 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1624635492
transform 1 0 50968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_426
timestamp 1624635492
transform 1 0 40296 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_414
timestamp 1624635492
transform 1 0 39192 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_423
timestamp 1624635492
transform 1 0 40020 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_441
timestamp 1624635492
transform 1 0 41676 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_429
timestamp 1624635492
transform 1 0 40572 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_435
timestamp 1624635492
transform 1 0 41124 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1624635492
transform 1 0 40480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_453
timestamp 1624635492
transform 1 0 42780 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_457
timestamp 1624635492
transform 1 0 43148 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_455
timestamp 1624635492
transform 1 0 42964 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_447
timestamp 1624635492
transform 1 0 42228 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1624635492
transform 1 0 43056 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1624635492
transform 1 0 44988 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_465
timestamp 1624635492
transform 1 0 43884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_481
timestamp 1624635492
transform 1 0 45356 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_469
timestamp 1624635492
transform 1 0 44252 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_498
timestamp 1624635492
transform 1 0 46920 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_486
timestamp 1624635492
transform 1 0 45816 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_495
timestamp 1624635492
transform 1 0 46644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_489
timestamp 1624635492
transform 1 0 46092 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1624635492
transform 1 0 45724 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _212_
timestamp 1624635492
transform -1 0 46644 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_510
timestamp 1624635492
transform 1 0 48024 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_514
timestamp 1624635492
transform 1 0 48392 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_507
timestamp 1624635492
transform 1 0 47748 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1624635492
transform 1 0 48300 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_534
timestamp 1624635492
transform 1 0 50232 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_522
timestamp 1624635492
transform 1 0 49128 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_526
timestamp 1624635492
transform 1 0 49496 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_543
timestamp 1624635492
transform 1 0 51060 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_538
timestamp 1624635492
transform 1 0 50600 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1624635492
transform 1 0 50968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_424
timestamp 1624635492
transform 1 0 40112 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_412
timestamp 1624635492
transform 1 0 39008 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_436
timestamp 1624635492
transform 1 0 41216 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_457
timestamp 1624635492
transform 1 0 43148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_448
timestamp 1624635492
transform 1 0 42320 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1624635492
transform 1 0 43056 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_481
timestamp 1624635492
transform 1 0 45356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_469
timestamp 1624635492
transform 1 0 44252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_493
timestamp 1624635492
transform 1 0 46460 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_514
timestamp 1624635492
transform 1 0 48392 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1624635492
transform 1 0 47564 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1624635492
transform 1 0 48300 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_526
timestamp 1624635492
transform 1 0 49496 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_538
timestamp 1624635492
transform 1 0 50600 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_420
timestamp 1624635492
transform 1 0 39744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_441
timestamp 1624635492
transform 1 0 41676 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_429
timestamp 1624635492
transform 1 0 40572 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1624635492
transform 1 0 40480 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_453
timestamp 1624635492
transform 1 0 42780 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_477
timestamp 1624635492
transform 1 0 44988 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_465
timestamp 1624635492
transform 1 0 43884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_498
timestamp 1624635492
transform 1 0 46920 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_486
timestamp 1624635492
transform 1 0 45816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1624635492
transform 1 0 45724 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_510
timestamp 1624635492
transform 1 0 48024 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_534
timestamp 1624635492
transform 1 0 50232 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_522
timestamp 1624635492
transform 1 0 49128 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_543
timestamp 1624635492
transform 1 0 51060 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1624635492
transform 1 0 50968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_424
timestamp 1624635492
transform 1 0 40112 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_412
timestamp 1624635492
transform 1 0 39008 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_436
timestamp 1624635492
transform 1 0 41216 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_457
timestamp 1624635492
transform 1 0 43148 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_448
timestamp 1624635492
transform 1 0 42320 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1624635492
transform 1 0 43056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_481
timestamp 1624635492
transform 1 0 45356 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_469
timestamp 1624635492
transform 1 0 44252 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_493
timestamp 1624635492
transform 1 0 46460 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_514
timestamp 1624635492
transform 1 0 48392 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1624635492
transform 1 0 47564 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1624635492
transform 1 0 48300 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_526
timestamp 1624635492
transform 1 0 49496 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_538
timestamp 1624635492
transform 1 0 50600 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_420
timestamp 1624635492
transform 1 0 39744 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_441
timestamp 1624635492
transform 1 0 41676 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_429
timestamp 1624635492
transform 1 0 40572 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1624635492
transform 1 0 40480 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_453
timestamp 1624635492
transform 1 0 42780 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_477
timestamp 1624635492
transform 1 0 44988 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_465
timestamp 1624635492
transform 1 0 43884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_498
timestamp 1624635492
transform 1 0 46920 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_486
timestamp 1624635492
transform 1 0 45816 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1624635492
transform 1 0 45724 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_510
timestamp 1624635492
transform 1 0 48024 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_534
timestamp 1624635492
transform 1 0 50232 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_522
timestamp 1624635492
transform 1 0 49128 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_543
timestamp 1624635492
transform 1 0 51060 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1624635492
transform 1 0 50968 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_416
timestamp 1624635492
transform 1 0 39376 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_424
timestamp 1624635492
transform 1 0 40112 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_412
timestamp 1624635492
transform 1 0 39008 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_441
timestamp 1624635492
transform 1 0 41676 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_429
timestamp 1624635492
transform 1 0 40572 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_436
timestamp 1624635492
transform 1 0 41216 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1624635492
transform 1 0 40480 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_458
timestamp 1624635492
transform 1 0 43240 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_452
timestamp 1624635492
transform 1 0 42688 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_457
timestamp 1624635492
transform 1 0 43148 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_448
timestamp 1624635492
transform 1 0 42320 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1624635492
transform 1 0 43056 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1624635492
transform 1 0 43056 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 1624635492
transform -1 0 42688 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_470
timestamp 1624635492
transform 1 0 44344 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_481
timestamp 1624635492
transform 1 0 45356 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_469
timestamp 1624635492
transform 1 0 44252 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_498
timestamp 1624635492
transform 1 0 46920 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_486
timestamp 1624635492
transform 1 0 45816 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_482
timestamp 1624635492
transform 1 0 45448 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_493
timestamp 1624635492
transform 1 0 46460 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1624635492
transform 1 0 45724 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A1
timestamp 1624635492
transform -1 0 47472 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A2
timestamp 1624635492
transform 1 0 47656 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_505
timestamp 1624635492
transform 1 0 47564 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_504
timestamp 1624635492
transform 1 0 47472 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1624635492
transform 1 0 48300 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A3
timestamp 1624635492
transform 1 0 47840 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__C1
timestamp 1624635492
transform 1 0 48392 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_508
timestamp 1624635492
transform 1 0 47840 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_512
timestamp 1624635492
transform 1 0 48208 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_510
timestamp 1624635492
transform 1 0 48024 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_4  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 48392 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_43_516
timestamp 1624635492
transform 1 0 48576 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_531
timestamp 1624635492
transform 1 0 49956 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_528
timestamp 1624635492
transform 1 0 49680 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_543
timestamp 1624635492
transform 1 0 51060 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_541
timestamp 1624635492
transform 1 0 50876 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_537
timestamp 1624635492
transform 1 0 50508 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_540
timestamp 1624635492
transform 1 0 50784 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__B1
timestamp 1624635492
transform -1 0 50508 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1624635492
transform 1 0 50968 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_424
timestamp 1624635492
transform 1 0 40112 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_412
timestamp 1624635492
transform 1 0 39008 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_436
timestamp 1624635492
transform 1 0 41216 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_457
timestamp 1624635492
transform 1 0 43148 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_448
timestamp 1624635492
transform 1 0 42320 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1624635492
transform 1 0 43056 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_481
timestamp 1624635492
transform 1 0 45356 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_469
timestamp 1624635492
transform 1 0 44252 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_493
timestamp 1624635492
transform 1 0 46460 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_514
timestamp 1624635492
transform 1 0 48392 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1624635492
transform 1 0 47564 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1624635492
transform 1 0 48300 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_526
timestamp 1624635492
transform 1 0 49496 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_538
timestamp 1624635492
transform 1 0 50600 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_420
timestamp 1624635492
transform 1 0 39744 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_441
timestamp 1624635492
transform 1 0 41676 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_429
timestamp 1624635492
transform 1 0 40572 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1624635492
transform 1 0 40480 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_453
timestamp 1624635492
transform 1 0 42780 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_477
timestamp 1624635492
transform 1 0 44988 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_465
timestamp 1624635492
transform 1 0 43884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_498
timestamp 1624635492
transform 1 0 46920 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_486
timestamp 1624635492
transform 1 0 45816 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1624635492
transform 1 0 45724 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_510
timestamp 1624635492
transform 1 0 48024 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_534
timestamp 1624635492
transform 1 0 50232 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_522
timestamp 1624635492
transform 1 0 49128 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_543
timestamp 1624635492
transform 1 0 51060 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1624635492
transform 1 0 50968 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_424
timestamp 1624635492
transform 1 0 40112 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_412
timestamp 1624635492
transform 1 0 39008 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_436
timestamp 1624635492
transform 1 0 41216 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_457
timestamp 1624635492
transform 1 0 43148 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_448
timestamp 1624635492
transform 1 0 42320 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1624635492
transform 1 0 43056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_481
timestamp 1624635492
transform 1 0 45356 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_469
timestamp 1624635492
transform 1 0 44252 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_493
timestamp 1624635492
transform 1 0 46460 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_514
timestamp 1624635492
transform 1 0 48392 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1624635492
transform 1 0 47564 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1624635492
transform 1 0 48300 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_526
timestamp 1624635492
transform 1 0 49496 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_538
timestamp 1624635492
transform 1 0 50600 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_420
timestamp 1624635492
transform 1 0 39744 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_441
timestamp 1624635492
transform 1 0 41676 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_429
timestamp 1624635492
transform 1 0 40572 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1624635492
transform 1 0 40480 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_453
timestamp 1624635492
transform 1 0 42780 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_477
timestamp 1624635492
transform 1 0 44988 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_465
timestamp 1624635492
transform 1 0 43884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_498
timestamp 1624635492
transform 1 0 46920 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_486
timestamp 1624635492
transform 1 0 45816 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1624635492
transform 1 0 45724 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_510
timestamp 1624635492
transform 1 0 48024 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_534
timestamp 1624635492
transform 1 0 50232 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_522
timestamp 1624635492
transform 1 0 49128 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_543
timestamp 1624635492
transform 1 0 51060 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1624635492
transform 1 0 50968 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_424
timestamp 1624635492
transform 1 0 40112 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_412
timestamp 1624635492
transform 1 0 39008 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_436
timestamp 1624635492
transform 1 0 41216 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_457
timestamp 1624635492
transform 1 0 43148 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_448
timestamp 1624635492
transform 1 0 42320 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1624635492
transform 1 0 43056 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_481
timestamp 1624635492
transform 1 0 45356 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_469
timestamp 1624635492
transform 1 0 44252 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_493
timestamp 1624635492
transform 1 0 46460 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_514
timestamp 1624635492
transform 1 0 48392 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1624635492
transform 1 0 47564 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1624635492
transform 1 0 48300 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_526
timestamp 1624635492
transform 1 0 49496 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_538
timestamp 1624635492
transform 1 0 50600 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_426
timestamp 1624635492
transform 1 0 40296 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_414
timestamp 1624635492
transform 1 0 39192 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_427
timestamp 1624635492
transform 1 0 40388 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_415
timestamp 1624635492
transform 1 0 39284 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _175_
timestamp 1624635492
transform -1 0 39192 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_438
timestamp 1624635492
transform 1 0 41400 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_441
timestamp 1624635492
transform 1 0 41676 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_429
timestamp 1624635492
transform 1 0 40572 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1624635492
transform 1 0 40480 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_457
timestamp 1624635492
transform 1 0 43148 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_450
timestamp 1624635492
transform 1 0 42504 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_453
timestamp 1624635492
transform 1 0 42780 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1624635492
transform 1 0 43056 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_481
timestamp 1624635492
transform 1 0 45356 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_469
timestamp 1624635492
transform 1 0 44252 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_477
timestamp 1624635492
transform 1 0 44988 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_465
timestamp 1624635492
transform 1 0 43884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_493
timestamp 1624635492
transform 1 0 46460 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_498
timestamp 1624635492
transform 1 0 46920 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_486
timestamp 1624635492
transform 1 0 45816 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1624635492
transform 1 0 45724 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_514
timestamp 1624635492
transform 1 0 48392 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1624635492
transform 1 0 47564 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_510
timestamp 1624635492
transform 1 0 48024 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__A
timestamp 1624635492
transform 1 0 48484 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1624635492
transform 1 0 48300 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_534
timestamp 1624635492
transform 1 0 50232 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_517
timestamp 1624635492
transform 1 0 48668 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_534
timestamp 1624635492
transform 1 0 50232 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_522
timestamp 1624635492
transform 1 0 49128 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  _051_
timestamp 1624635492
transform 1 0 49036 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_51_546
timestamp 1624635492
transform 1 0 51336 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_543
timestamp 1624635492
transform 1 0 51060 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1624635492
transform 1 0 50968 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_427
timestamp 1624635492
transform 1 0 40388 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_415
timestamp 1624635492
transform 1 0 39284 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__B2
timestamp 1624635492
transform 1 0 39100 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_441
timestamp 1624635492
transform 1 0 41676 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_429
timestamp 1624635492
transform 1 0 40572 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1624635492
transform 1 0 40480 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_453
timestamp 1624635492
transform 1 0 42780 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_477
timestamp 1624635492
transform 1 0 44988 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_465
timestamp 1624635492
transform 1 0 43884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_498
timestamp 1624635492
transform 1 0 46920 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_486
timestamp 1624635492
transform 1 0 45816 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1624635492
transform 1 0 45724 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_510
timestamp 1624635492
transform 1 0 48024 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_534
timestamp 1624635492
transform 1 0 50232 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_522
timestamp 1624635492
transform 1 0 49128 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_543
timestamp 1624635492
transform 1 0 51060 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1624635492
transform 1 0 50968 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_560
timestamp 1624635492
transform 1 0 52624 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_548
timestamp 1624635492
transform 1 0 51520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1684
timestamp 1624635492
transform 1 0 53360 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_581
timestamp 1624635492
transform 1 0 54556 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_569
timestamp 1624635492
transform 1 0 53452 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_609
timestamp 1624635492
transform 1 0 57132 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1624635492
transform 1 0 56028 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_593
timestamp 1624635492
transform 1 0 55660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _207_
timestamp 1624635492
transform -1 0 56028 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_626
timestamp 1624635492
transform 1 0 58696 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1624635492
transform 1 0 58236 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1685
timestamp 1624635492
transform 1 0 58604 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_650
timestamp 1624635492
transform 1 0 60904 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_638
timestamp 1624635492
transform 1 0 59800 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_672
timestamp 1624635492
transform 1 0 62928 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_660
timestamp 1624635492
transform 1 0 61824 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_656
timestamp 1624635492
transform 1 0 61456 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _250_
timestamp 1624635492
transform -1 0 61824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_680
timestamp 1624635492
transform 1 0 63664 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1686
timestamp 1624635492
transform 1 0 63848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_565
timestamp 1624635492
transform 1 0 53084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_553
timestamp 1624635492
transform 1 0 51980 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_589
timestamp 1624635492
transform 1 0 55292 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_577
timestamp 1624635492
transform 1 0 54188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_610
timestamp 1624635492
transform 1 0 57224 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_598
timestamp 1624635492
transform 1 0 56120 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1690
timestamp 1624635492
transform 1 0 56028 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_622
timestamp 1624635492
transform 1 0 58328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_655
timestamp 1624635492
transform 1 0 61364 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_646
timestamp 1624635492
transform 1 0 60536 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_634
timestamp 1624635492
transform 1 0 59432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1691
timestamp 1624635492
transform 1 0 61272 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_667
timestamp 1624635492
transform 1 0 62468 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_679
timestamp 1624635492
transform 1 0 63572 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_560
timestamp 1624635492
transform 1 0 52624 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_548
timestamp 1624635492
transform 1 0 51520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1695
timestamp 1624635492
transform 1 0 53360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_581
timestamp 1624635492
transform 1 0 54556 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_569
timestamp 1624635492
transform 1 0 53452 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_605
timestamp 1624635492
transform 1 0 56764 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_593
timestamp 1624635492
transform 1 0 55660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_626
timestamp 1624635492
transform 1 0 58696 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1624635492
transform 1 0 57868 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1696
timestamp 1624635492
transform 1 0 58604 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_650
timestamp 1624635492
transform 1 0 60904 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_638
timestamp 1624635492
transform 1 0 59800 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_671
timestamp 1624635492
transform 1 0 62836 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_659
timestamp 1624635492
transform 1 0 61732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _161_
timestamp 1624635492
transform -1 0 61732 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_679
timestamp 1624635492
transform 1 0 63572 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1697
timestamp 1624635492
transform 1 0 63848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_565
timestamp 1624635492
transform 1 0 53084 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_553
timestamp 1624635492
transform 1 0 51980 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_560
timestamp 1624635492
transform 1 0 52624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_548
timestamp 1624635492
transform 1 0 51520 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1706
timestamp 1624635492
transform 1 0 53360 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_581
timestamp 1624635492
transform 1 0 54556 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_569
timestamp 1624635492
transform 1 0 53452 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_584
timestamp 1624635492
transform 1 0 54832 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_572
timestamp 1624635492
transform 1 0 53728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_605
timestamp 1624635492
transform 1 0 56764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_593
timestamp 1624635492
transform 1 0 55660 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_610
timestamp 1624635492
transform 1 0 57224 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_598
timestamp 1624635492
transform 1 0 56120 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_596
timestamp 1624635492
transform 1 0 55936 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1701
timestamp 1624635492
transform 1 0 56028 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_626
timestamp 1624635492
transform 1 0 58696 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1624635492
transform 1 0 57868 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_622
timestamp 1624635492
transform 1 0 58328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1707
timestamp 1624635492
transform 1 0 58604 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_650
timestamp 1624635492
transform 1 0 60904 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_638
timestamp 1624635492
transform 1 0 59800 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_655
timestamp 1624635492
transform 1 0 61364 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_646
timestamp 1624635492
transform 1 0 60536 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_634
timestamp 1624635492
transform 1 0 59432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1702
timestamp 1624635492
transform 1 0 61272 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_674
timestamp 1624635492
transform 1 0 63112 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_662
timestamp 1624635492
transform 1 0 62008 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_667
timestamp 1624635492
transform 1 0 62468 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_679
timestamp 1624635492
transform 1 0 63572 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1708
timestamp 1624635492
transform 1 0 63848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_564
timestamp 1624635492
transform 1 0 52992 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_552
timestamp 1624635492
transform 1 0 51888 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1624635492
transform 1 0 51796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _215_
timestamp 1624635492
transform -1 0 53544 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_581
timestamp 1624635492
transform 1 0 54556 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_578
timestamp 1624635492
transform 1 0 54280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_570
timestamp 1624635492
transform 1 0 53544 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1624635492
transform 1 0 54464 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_610
timestamp 1624635492
transform 1 0 57224 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_605
timestamp 1624635492
transform 1 0 56764 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_593
timestamp 1624635492
transform 1 0 55660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1624635492
transform 1 0 57132 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_622
timestamp 1624635492
transform 1 0 58328 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_651
timestamp 1624635492
transform 1 0 60996 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_639
timestamp 1624635492
transform 1 0 59892 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_634
timestamp 1624635492
transform 1 0 59432 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1624635492
transform 1 0 59800 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_668
timestamp 1624635492
transform 1 0 62560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_663
timestamp 1624635492
transform 1 0 62100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1624635492
transform 1 0 62468 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_680
timestamp 1624635492
transform 1 0 63664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_562
timestamp 1624635492
transform 1 0 52808 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_550
timestamp 1624635492
transform 1 0 51704 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_583
timestamp 1624635492
transform 1 0 54740 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_571
timestamp 1624635492
transform 1 0 53636 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1624635492
transform 1 0 53544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_607
timestamp 1624635492
transform 1 0 56948 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_595
timestamp 1624635492
transform 1 0 55844 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_628
timestamp 1624635492
transform 1 0 58880 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_619
timestamp 1624635492
transform 1 0 58052 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1624635492
transform 1 0 58788 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_652
timestamp 1624635492
transform 1 0 61088 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_640
timestamp 1624635492
transform 1 0 59984 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_676
timestamp 1624635492
transform 1 0 63296 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_664
timestamp 1624635492
transform 1 0 62192 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_567
timestamp 1624635492
transform 1 0 53268 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_555
timestamp 1624635492
transform 1 0 52164 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_579
timestamp 1624635492
transform 1 0 54372 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_600
timestamp 1624635492
transform 1 0 56304 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_591
timestamp 1624635492
transform 1 0 55476 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1624635492
transform 1 0 56212 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_624
timestamp 1624635492
transform 1 0 58512 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_612
timestamp 1624635492
transform 1 0 57408 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_648
timestamp 1624635492
transform 1 0 60720 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_636
timestamp 1624635492
transform 1 0 59616 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_669
timestamp 1624635492
transform 1 0 62652 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_657
timestamp 1624635492
transform 1 0 61548 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1624635492
transform 1 0 61456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_681
timestamp 1624635492
transform 1 0 63756 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_562
timestamp 1624635492
transform 1 0 52808 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_550
timestamp 1624635492
transform 1 0 51704 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_583
timestamp 1624635492
transform 1 0 54740 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_571
timestamp 1624635492
transform 1 0 53636 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1624635492
transform 1 0 53544 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_607
timestamp 1624635492
transform 1 0 56948 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_595
timestamp 1624635492
transform 1 0 55844 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_628
timestamp 1624635492
transform 1 0 58880 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_619
timestamp 1624635492
transform 1 0 58052 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1624635492
transform 1 0 58788 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_652
timestamp 1624635492
transform 1 0 61088 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_640
timestamp 1624635492
transform 1 0 59984 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_676
timestamp 1624635492
transform 1 0 63296 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_664
timestamp 1624635492
transform 1 0 62192 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_567
timestamp 1624635492
transform 1 0 53268 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_555
timestamp 1624635492
transform 1 0 52164 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_579
timestamp 1624635492
transform 1 0 54372 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_600
timestamp 1624635492
transform 1 0 56304 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_591
timestamp 1624635492
transform 1 0 55476 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1624635492
transform 1 0 56212 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_624
timestamp 1624635492
transform 1 0 58512 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_612
timestamp 1624635492
transform 1 0 57408 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_648
timestamp 1624635492
transform 1 0 60720 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_636
timestamp 1624635492
transform 1 0 59616 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_669
timestamp 1624635492
transform 1 0 62652 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_657
timestamp 1624635492
transform 1 0 61548 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1624635492
transform 1 0 61456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_681
timestamp 1624635492
transform 1 0 63756 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_567
timestamp 1624635492
transform 1 0 53268 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_555
timestamp 1624635492
transform 1 0 52164 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_562
timestamp 1624635492
transform 1 0 52808 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_550
timestamp 1624635492
transform 1 0 51704 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_588
timestamp 1624635492
transform 1 0 55200 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_576
timestamp 1624635492
transform 1 0 54096 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_573
timestamp 1624635492
transform 1 0 53820 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_583
timestamp 1624635492
transform 1 0 54740 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_571
timestamp 1624635492
transform 1 0 53636 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__B
timestamp 1624635492
transform 1 0 53912 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1624635492
transform 1 0 53544 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1624635492
transform 1 0 56212 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__RESET_B
timestamp 1624635492
transform 1 0 55660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_595
timestamp 1624635492
transform 1 0 55844 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_592
timestamp 1624635492
transform 1 0 55568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_595
timestamp 1624635492
transform 1 0 55844 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_600
timestamp 1624635492
transform 1 0 56304 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__D
timestamp 1624635492
transform -1 0 56672 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_601
timestamp 1624635492
transform 1 0 56396 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 56672 0 -1 23392
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_37_604
timestamp 1624635492
transform 1 0 56672 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_625
timestamp 1624635492
transform 1 0 58604 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_628
timestamp 1624635492
transform 1 0 58880 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_624
timestamp 1624635492
transform 1 0 58512 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_616
timestamp 1624635492
transform 1 0 57776 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1624635492
transform 1 0 58788 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_655
timestamp 1624635492
transform 1 0 61364 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_649
timestamp 1624635492
transform 1 0 60812 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_637
timestamp 1624635492
transform 1 0 59708 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_652
timestamp 1624635492
transform 1 0 61088 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_640
timestamp 1624635492
transform 1 0 59984 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_669
timestamp 1624635492
transform 1 0 62652 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_657
timestamp 1624635492
transform 1 0 61548 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_675
timestamp 1624635492
transform 1 0 63204 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_663
timestamp 1624635492
transform 1 0 62100 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1624635492
transform 1 0 61456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _154_
timestamp 1624635492
transform 1 0 61824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_681
timestamp 1624635492
transform 1 0 63756 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_566
timestamp 1624635492
transform 1 0 53176 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_562
timestamp 1624635492
transform 1 0 52808 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_550
timestamp 1624635492
transform 1 0 51704 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__C
timestamp 1624635492
transform 1 0 52992 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_587
timestamp 1624635492
transform 1 0 55108 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_574
timestamp 1624635492
transform 1 0 53912 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_571
timestamp 1624635492
transform 1 0 53636 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1624635492
transform 1 0 53728 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1624635492
transform 1 0 53544 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 54280 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_39_610
timestamp 1624635492
transform 1 0 57224 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_602
timestamp 1624635492
transform 1 0 56488 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_599
timestamp 1624635492
transform 1 0 56212 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__CLK
timestamp 1624635492
transform 1 0 56304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _135_
timestamp 1624635492
transform -1 0 57592 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_628
timestamp 1624635492
transform 1 0 58880 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_626
timestamp 1624635492
transform 1 0 58696 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_614
timestamp 1624635492
transform 1 0 57592 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1624635492
transform 1 0 58788 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_652
timestamp 1624635492
transform 1 0 61088 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_640
timestamp 1624635492
transform 1 0 59984 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_676
timestamp 1624635492
transform 1 0 63296 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_664
timestamp 1624635492
transform 1 0 62192 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_567
timestamp 1624635492
transform 1 0 53268 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_555
timestamp 1624635492
transform 1 0 52164 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_579
timestamp 1624635492
transform 1 0 54372 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_575
timestamp 1624635492
transform 1 0 54004 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _306_
timestamp 1624635492
transform -1 0 54372 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_600
timestamp 1624635492
transform 1 0 56304 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_591
timestamp 1624635492
transform 1 0 55476 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1624635492
transform 1 0 56212 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_624
timestamp 1624635492
transform 1 0 58512 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_612
timestamp 1624635492
transform 1 0 57408 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_648
timestamp 1624635492
transform 1 0 60720 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_636
timestamp 1624635492
transform 1 0 59616 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1624635492
transform 1 0 62652 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1624635492
transform 1 0 61548 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1624635492
transform 1 0 61456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1624635492
transform 1 0 63756 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_562
timestamp 1624635492
transform 1 0 52808 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_550
timestamp 1624635492
transform 1 0 51704 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_583
timestamp 1624635492
transform 1 0 54740 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_571
timestamp 1624635492
transform 1 0 53636 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1624635492
transform 1 0 53544 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_607
timestamp 1624635492
transform 1 0 56948 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_595
timestamp 1624635492
transform 1 0 55844 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_628
timestamp 1624635492
transform 1 0 58880 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_619
timestamp 1624635492
transform 1 0 58052 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1624635492
transform 1 0 58788 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_652
timestamp 1624635492
transform 1 0 61088 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_640
timestamp 1624635492
transform 1 0 59984 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_676
timestamp 1624635492
transform 1 0 63296 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_664
timestamp 1624635492
transform 1 0 62192 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_567
timestamp 1624635492
transform 1 0 53268 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_555
timestamp 1624635492
transform 1 0 52164 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_579
timestamp 1624635492
transform 1 0 54372 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_600
timestamp 1624635492
transform 1 0 56304 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_591
timestamp 1624635492
transform 1 0 55476 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1624635492
transform 1 0 56212 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_624
timestamp 1624635492
transform 1 0 58512 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_612
timestamp 1624635492
transform 1 0 57408 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_648
timestamp 1624635492
transform 1 0 60720 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_636
timestamp 1624635492
transform 1 0 59616 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1624635492
transform 1 0 62652 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1624635492
transform 1 0 61548 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1624635492
transform 1 0 61456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1624635492
transform 1 0 63756 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_567
timestamp 1624635492
transform 1 0 53268 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_555
timestamp 1624635492
transform 1 0 52164 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_564
timestamp 1624635492
transform 1 0 52992 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_552
timestamp 1624635492
transform 1 0 51888 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_579
timestamp 1624635492
transform 1 0 54372 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_589
timestamp 1624635492
transform 1 0 55292 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_583
timestamp 1624635492
transform 1 0 54740 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_571
timestamp 1624635492
transform 1 0 53636 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1624635492
transform 1 0 53544 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_600
timestamp 1624635492
transform 1 0 56304 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_591
timestamp 1624635492
transform 1 0 55476 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_608
timestamp 1624635492
transform 1 0 57040 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_596
timestamp 1624635492
transform 1 0 55936 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1624635492
transform 1 0 56212 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 55936 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_624
timestamp 1624635492
transform 1 0 58512 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_612
timestamp 1624635492
transform 1 0 57408 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_628
timestamp 1624635492
transform 1 0 58880 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_626
timestamp 1624635492
transform 1 0 58696 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_620
timestamp 1624635492
transform 1 0 58144 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1624635492
transform 1 0 58788 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_648
timestamp 1624635492
transform 1 0 60720 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_636
timestamp 1624635492
transform 1 0 59616 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_652
timestamp 1624635492
transform 1 0 61088 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_640
timestamp 1624635492
transform 1 0 59984 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_672
timestamp 1624635492
transform 1 0 62928 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1624635492
transform 1 0 61548 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_676
timestamp 1624635492
transform 1 0 63296 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_664
timestamp 1624635492
transform 1 0 62192 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1624635492
transform 1 0 61456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _317_
timestamp 1624635492
transform -1 0 62928 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_562
timestamp 1624635492
transform 1 0 52808 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_550
timestamp 1624635492
transform 1 0 51704 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_583
timestamp 1624635492
transform 1 0 54740 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_571
timestamp 1624635492
transform 1 0 53636 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1624635492
transform 1 0 53544 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_607
timestamp 1624635492
transform 1 0 56948 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_595
timestamp 1624635492
transform 1 0 55844 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_628
timestamp 1624635492
transform 1 0 58880 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_619
timestamp 1624635492
transform 1 0 58052 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1624635492
transform 1 0 58788 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_652
timestamp 1624635492
transform 1 0 61088 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_640
timestamp 1624635492
transform 1 0 59984 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_676
timestamp 1624635492
transform 1 0 63296 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_664
timestamp 1624635492
transform 1 0 62192 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_567
timestamp 1624635492
transform 1 0 53268 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_555
timestamp 1624635492
transform 1 0 52164 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_579
timestamp 1624635492
transform 1 0 54372 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_600
timestamp 1624635492
transform 1 0 56304 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_591
timestamp 1624635492
transform 1 0 55476 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1624635492
transform 1 0 56212 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_624
timestamp 1624635492
transform 1 0 58512 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_612
timestamp 1624635492
transform 1 0 57408 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_648
timestamp 1624635492
transform 1 0 60720 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_636
timestamp 1624635492
transform 1 0 59616 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_669
timestamp 1624635492
transform 1 0 62652 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_657
timestamp 1624635492
transform 1 0 61548 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1624635492
transform 1 0 61456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_681
timestamp 1624635492
transform 1 0 63756 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_562
timestamp 1624635492
transform 1 0 52808 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_550
timestamp 1624635492
transform 1 0 51704 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_583
timestamp 1624635492
transform 1 0 54740 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_571
timestamp 1624635492
transform 1 0 53636 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1624635492
transform 1 0 53544 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_607
timestamp 1624635492
transform 1 0 56948 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_595
timestamp 1624635492
transform 1 0 55844 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_628
timestamp 1624635492
transform 1 0 58880 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_619
timestamp 1624635492
transform 1 0 58052 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1624635492
transform 1 0 58788 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_648
timestamp 1624635492
transform 1 0 60720 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_644
timestamp 1624635492
transform 1 0 60352 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_640
timestamp 1624635492
transform 1 0 59984 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _246_
timestamp 1624635492
transform -1 0 60720 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_672
timestamp 1624635492
transform 1 0 62928 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_660
timestamp 1624635492
transform 1 0 61824 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_567
timestamp 1624635492
transform 1 0 53268 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_555
timestamp 1624635492
transform 1 0 52164 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_586
timestamp 1624635492
transform 1 0 55016 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_579
timestamp 1624635492
transform 1 0 54372 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _101_
timestamp 1624635492
transform -1 0 55016 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_600
timestamp 1624635492
transform 1 0 56304 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_598
timestamp 1624635492
transform 1 0 56120 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1624635492
transform 1 0 56212 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_624
timestamp 1624635492
transform 1 0 58512 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_612
timestamp 1624635492
transform 1 0 57408 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_648
timestamp 1624635492
transform 1 0 60720 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_636
timestamp 1624635492
transform 1 0 59616 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_669
timestamp 1624635492
transform 1 0 62652 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_657
timestamp 1624635492
transform 1 0 61548 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1624635492
transform 1 0 61456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_681
timestamp 1624635492
transform 1 0 63756 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_562
timestamp 1624635492
transform 1 0 52808 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_550
timestamp 1624635492
transform 1 0 51704 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_583
timestamp 1624635492
transform 1 0 54740 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_571
timestamp 1624635492
transform 1 0 53636 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1624635492
transform 1 0 53544 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_607
timestamp 1624635492
transform 1 0 56948 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_595
timestamp 1624635492
transform 1 0 55844 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_628
timestamp 1624635492
transform 1 0 58880 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_619
timestamp 1624635492
transform 1 0 58052 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1624635492
transform 1 0 58788 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _304_
timestamp 1624635492
transform -1 0 59524 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_647
timestamp 1624635492
transform 1 0 60628 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_635
timestamp 1624635492
transform 1 0 59524 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_671
timestamp 1624635492
transform 1 0 62836 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_659
timestamp 1624635492
transform 1 0 61732 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_558
timestamp 1624635492
transform 1 0 52440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_567
timestamp 1624635492
transform 1 0 53268 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_555
timestamp 1624635492
transform 1 0 52164 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_583
timestamp 1624635492
transform 1 0 54740 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_571
timestamp 1624635492
transform 1 0 53636 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_579
timestamp 1624635492
transform 1 0 54372 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1624635492
transform 1 0 53544 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_607
timestamp 1624635492
transform 1 0 56948 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_595
timestamp 1624635492
transform 1 0 55844 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_600
timestamp 1624635492
transform 1 0 56304 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_591
timestamp 1624635492
transform 1 0 55476 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1624635492
transform 1 0 56212 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_628
timestamp 1624635492
transform 1 0 58880 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_619
timestamp 1624635492
transform 1 0 58052 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_624
timestamp 1624635492
transform 1 0 58512 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_612
timestamp 1624635492
transform 1 0 57408 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1624635492
transform 1 0 58788 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_652
timestamp 1624635492
transform 1 0 61088 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_640
timestamp 1624635492
transform 1 0 59984 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_648
timestamp 1624635492
transform 1 0 60720 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_636
timestamp 1624635492
transform 1 0 59616 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_676
timestamp 1624635492
transform 1 0 63296 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_664
timestamp 1624635492
transform 1 0 62192 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_669
timestamp 1624635492
transform 1 0 62652 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_657
timestamp 1624635492
transform 1 0 61548 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1624635492
transform 1 0 61456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_681
timestamp 1624635492
transform 1 0 63756 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_567
timestamp 1624635492
transform 1 0 53268 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_555
timestamp 1624635492
transform 1 0 52164 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_579
timestamp 1624635492
transform 1 0 54372 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_600
timestamp 1624635492
transform 1 0 56304 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_591
timestamp 1624635492
transform 1 0 55476 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1624635492
transform 1 0 56212 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_624
timestamp 1624635492
transform 1 0 58512 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_612
timestamp 1624635492
transform 1 0 57408 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_648
timestamp 1624635492
transform 1 0 60720 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_636
timestamp 1624635492
transform 1 0 59616 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_669
timestamp 1624635492
transform 1 0 62652 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_657
timestamp 1624635492
transform 1 0 61548 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1624635492
transform 1 0 61456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_681
timestamp 1624635492
transform 1 0 63756 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_695
timestamp 1624635492
transform 1 0 65044 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_683
timestamp 1624635492
transform 1 0 63940 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_707
timestamp 1624635492
transform 1 0 66148 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_719
timestamp 1624635492
transform 1 0 67252 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_731
timestamp 1624635492
transform 1 0 68356 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_295
timestamp 1624635492
transform -1 0 68816 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_695
timestamp 1624635492
transform 1 0 65044 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_683
timestamp 1624635492
transform 1 0 63940 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_691
timestamp 1624635492
transform 1 0 64676 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_707
timestamp 1624635492
transform 1 0 66148 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_703
timestamp 1624635492
transform 1 0 65780 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_719
timestamp 1624635492
transform 1 0 67252 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_721
timestamp 1624635492
transform 1 0 67436 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_718
timestamp 1624635492
transform 1 0 67160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_712
timestamp 1624635492
transform 1 0 66608 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output438_A
timestamp 1624635492
transform -1 0 67436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1692
timestamp 1624635492
transform 1 0 66516 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_731
timestamp 1624635492
transform 1 0 68356 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_729
timestamp 1624635492
transform 1 0 68172 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output438
timestamp 1624635492
transform 1 0 67804 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_299
timestamp 1624635492
transform -1 0 68816 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_297
timestamp 1624635492
transform -1 0 68816 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_691
timestamp 1624635492
transform 1 0 64676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_703
timestamp 1624635492
transform 1 0 65780 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_712
timestamp 1624635492
transform 1 0 66608 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1703
timestamp 1624635492
transform 1 0 66516 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_732
timestamp 1624635492
transform 1 0 68448 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_724
timestamp 1624635492
transform 1 0 67712 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_301
timestamp 1624635492
transform -1 0 68816 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_695
timestamp 1624635492
transform 1 0 65044 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_683
timestamp 1624635492
transform 1 0 63940 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_707
timestamp 1624635492
transform 1 0 66148 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_721
timestamp 1624635492
transform 1 0 67436 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output400_A
timestamp 1624635492
transform -1 0 67436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1624635492
transform 1 0 68172 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output400
timestamp 1624635492
transform 1 0 67804 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_303
timestamp 1624635492
transform -1 0 68816 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_685
timestamp 1624635492
transform 1 0 64124 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_692
timestamp 1624635492
transform 1 0 64768 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1624635492
transform 1 0 64032 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_697
timestamp 1624635492
transform 1 0 65228 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_697
timestamp 1624635492
transform 1 0 65228 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1624635492
transform 1 0 65136 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_717
timestamp 1624635492
transform 1 0 67068 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_709
timestamp 1624635492
transform 1 0 66332 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_721
timestamp 1624635492
transform 1 0 67436 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_709
timestamp 1624635492
transform 1 0 66332 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 67528 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1624635492
transform 1 0 68172 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_722
timestamp 1624635492
transform 1 0 67528 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_732
timestamp 1624635492
transform 1 0 68448 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_726
timestamp 1624635492
transform 1 0 67896 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1624635492
transform -1 0 68172 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1624635492
transform 1 0 67804 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 68816 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 68816 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_693
timestamp 1624635492
transform 1 0 64860 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_705
timestamp 1624635492
transform 1 0 65964 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_714
timestamp 1624635492
transform 1 0 66792 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1624635492
transform 1 0 66700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_732
timestamp 1624635492
transform 1 0 68448 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_726
timestamp 1624635492
transform 1 0 67896 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 68816 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_693
timestamp 1624635492
transform 1 0 64860 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_685
timestamp 1624635492
transform 1 0 64124 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1624635492
transform 1 0 64032 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_705
timestamp 1624635492
transform 1 0 65964 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_697
timestamp 1624635492
transform 1 0 65228 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_714
timestamp 1624635492
transform 1 0 66792 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_721
timestamp 1624635492
transform 1 0 67436 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_717
timestamp 1624635492
transform 1 0 67068 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_709
timestamp 1624635492
transform 1 0 66332 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output439_A
timestamp 1624635492
transform 1 0 67252 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1624635492
transform 1 0 66700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_732
timestamp 1624635492
transform 1 0 68448 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_726
timestamp 1624635492
transform 1 0 67896 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1624635492
transform 1 0 68172 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output439
timestamp 1624635492
transform 1 0 67804 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1624635492
transform -1 0 68816 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1624635492
transform -1 0 68816 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_685
timestamp 1624635492
transform 1 0 64124 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_683
timestamp 1624635492
transform 1 0 63940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1624635492
transform 1 0 64032 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_697
timestamp 1624635492
transform 1 0 65228 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_721
timestamp 1624635492
transform 1 0 67436 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_709
timestamp 1624635492
transform 1 0 66332 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1624635492
transform -1 0 68816 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_693
timestamp 1624635492
transform 1 0 64860 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_705
timestamp 1624635492
transform 1 0 65964 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_721
timestamp 1624635492
transform 1 0 67436 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_718
timestamp 1624635492
transform 1 0 67160 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_714
timestamp 1624635492
transform 1 0 66792 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output401_A
timestamp 1624635492
transform -1 0 67436 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1624635492
transform 1 0 66700 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_729
timestamp 1624635492
transform 1 0 68172 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output401
timestamp 1624635492
transform 1 0 67804 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1624635492
transform -1 0 68816 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_693
timestamp 1624635492
transform 1 0 64860 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1624635492
transform 1 0 64124 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1624635492
transform 1 0 64032 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_705
timestamp 1624635492
transform 1 0 65964 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_697
timestamp 1624635492
transform 1 0 65228 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_714
timestamp 1624635492
transform 1 0 66792 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_721
timestamp 1624635492
transform 1 0 67436 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_709
timestamp 1624635492
transform 1 0 66332 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1624635492
transform 1 0 66700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_729
timestamp 1624635492
transform 1 0 68172 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1624635492
transform -1 0 68816 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1624635492
transform -1 0 68816 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _127_
timestamp 1624635492
transform -1 0 68172 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_692
timestamp 1624635492
transform 1 0 64768 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_685
timestamp 1624635492
transform 1 0 64124 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1624635492
transform 1 0 64032 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _318_
timestamp 1624635492
transform -1 0 64768 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_704
timestamp 1624635492
transform 1 0 65872 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_716
timestamp 1624635492
transform 1 0 66976 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 67528 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1624635492
transform 1 0 68172 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_722
timestamp 1624635492
transform 1 0 67528 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1624635492
transform -1 0 68172 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1624635492
transform -1 0 68816 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1624635492
transform 1 0 64124 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_693
timestamp 1624635492
transform 1 0 64860 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1624635492
transform 1 0 64032 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_697
timestamp 1624635492
transform 1 0 65228 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_708
timestamp 1624635492
transform 1 0 66240 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _102_
timestamp 1624635492
transform -1 0 66240 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_721
timestamp 1624635492
transform 1 0 67436 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_717
timestamp 1624635492
transform 1 0 67068 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_709
timestamp 1624635492
transform 1 0 66332 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_714
timestamp 1624635492
transform 1 0 66792 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_712
timestamp 1624635492
transform 1 0 66608 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output440_A
timestamp 1624635492
transform 1 0 67252 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1624635492
transform 1 0 66700 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1624635492
transform 1 0 68172 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_732
timestamp 1624635492
transform 1 0 68448 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_726
timestamp 1624635492
transform 1 0 67896 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output440
timestamp 1624635492
transform 1 0 67804 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1624635492
transform -1 0 68816 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1624635492
transform -1 0 68816 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_684
timestamp 1624635492
transform 1 0 64032 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_708
timestamp 1624635492
transform 1 0 66240 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_696
timestamp 1624635492
transform 1 0 65136 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_714
timestamp 1624635492
transform 1 0 66792 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_712
timestamp 1624635492
transform 1 0 66608 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1624635492
transform 1 0 66700 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_732
timestamp 1624635492
transform 1 0 68448 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_726
timestamp 1624635492
transform 1 0 67896 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1624635492
transform -1 0 68816 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1624635492
transform 1 0 64124 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1624635492
transform 1 0 64032 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1624635492
transform 1 0 65228 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_721
timestamp 1624635492
transform 1 0 67436 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_717
timestamp 1624635492
transform 1 0 67068 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_709
timestamp 1624635492
transform 1 0 66332 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output402_A
timestamp 1624635492
transform 1 0 67252 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1624635492
transform 1 0 68172 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output402
timestamp 1624635492
transform 1 0 67804 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1624635492
transform -1 0 68816 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1624635492
transform 1 0 64124 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_693
timestamp 1624635492
transform 1 0 64860 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1624635492
transform 1 0 64032 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _267_
timestamp 1624635492
transform -1 0 65228 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1624635492
transform 1 0 65228 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_697
timestamp 1624635492
transform 1 0 65228 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_721
timestamp 1624635492
transform 1 0 67436 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1624635492
transform 1 0 66332 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_714
timestamp 1624635492
transform 1 0 66792 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_709
timestamp 1624635492
transform 1 0 66332 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1624635492
transform 1 0 66700 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_732
timestamp 1624635492
transform 1 0 68448 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_726
timestamp 1624635492
transform 1 0 67896 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1624635492
transform -1 0 68816 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1624635492
transform -1 0 68816 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_693
timestamp 1624635492
transform 1 0 64860 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_705
timestamp 1624635492
transform 1 0 65964 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_714
timestamp 1624635492
transform 1 0 66792 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1624635492
transform 1 0 66700 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_732
timestamp 1624635492
transform 1 0 68448 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_726
timestamp 1624635492
transform 1 0 67896 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1624635492
transform -1 0 68816 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_693
timestamp 1624635492
transform 1 0 64860 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1624635492
transform 1 0 64124 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_683
timestamp 1624635492
transform 1 0 63940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1624635492
transform 1 0 64032 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_705
timestamp 1624635492
transform 1 0 65964 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1624635492
transform 1 0 65228 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_714
timestamp 1624635492
transform 1 0 66792 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_721
timestamp 1624635492
transform 1 0 67436 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1624635492
transform 1 0 66332 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 67528 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1624635492
transform 1 0 66700 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_729
timestamp 1624635492
transform 1 0 68172 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_722
timestamp 1624635492
transform 1 0 67528 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1624635492
transform -1 0 68172 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1624635492
transform -1 0 68816 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1624635492
transform -1 0 68816 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1624635492
transform 1 0 64124 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1624635492
transform 1 0 64032 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1624635492
transform 1 0 65228 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_721
timestamp 1624635492
transform 1 0 67436 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1624635492
transform 1 0 66332 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1624635492
transform -1 0 68816 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_693
timestamp 1624635492
transform 1 0 64860 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_705
timestamp 1624635492
transform 1 0 65964 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_714
timestamp 1624635492
transform 1 0 66792 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1624635492
transform 1 0 66700 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_729
timestamp 1624635492
transform 1 0 68172 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_722
timestamp 1624635492
transform 1 0 67528 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output441
timestamp 1624635492
transform 1 0 67804 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1624635492
transform -1 0 68816 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_12
timestamp 1624635492
transform 1 0 2208 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_6
timestamp 1624635492
transform 1 0 1656 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1624635492
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1624635492
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 2208 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1624635492
transform -1 0 1656 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1624635492
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1624635492
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1624635492
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_28
timestamp 1624635492
transform 1 0 3680 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1624635492
transform 1 0 3312 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1624635492
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1624635492
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1624635492
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_54
timestamp 1624635492
transform 1 0 6072 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1624635492
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_58
timestamp 1624635492
transform 1 0 6440 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_51
timestamp 1624635492
transform 1 0 5796 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1624635492
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_78
timestamp 1624635492
transform 1 0 8280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_66
timestamp 1624635492
transform 1 0 7176 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_70
timestamp 1624635492
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_99
timestamp 1624635492
transform 1 0 10212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_87
timestamp 1624635492
transform 1 0 9108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_94
timestamp 1624635492
transform 1 0 9752 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_82
timestamp 1624635492
transform 1 0 8648 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1624635492
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_111
timestamp 1624635492
transform 1 0 11316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_115
timestamp 1624635492
transform 1 0 11684 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_106
timestamp 1624635492
transform 1 0 10856 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1624635492
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_135
timestamp 1624635492
transform 1 0 13524 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_123
timestamp 1624635492
transform 1 0 12420 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_127
timestamp 1624635492
transform 1 0 12788 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1624635492
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1624635492
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1624635492
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1624635492
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1624635492
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_58
timestamp 1624635492
transform 1 0 6440 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_51
timestamp 1624635492
transform 1 0 5796 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1624635492
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_77
timestamp 1624635492
transform 1 0 8188 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_65
timestamp 1624635492
transform 1 0 7084 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _180_
timestamp 1624635492
transform 1 0 6808 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_89
timestamp 1624635492
transform 1 0 9292 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_115
timestamp 1624635492
transform 1 0 11684 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1624635492
transform 1 0 11500 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_101
timestamp 1624635492
transform 1 0 10396 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1624635492
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_127
timestamp 1624635492
transform 1 0 12788 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1624635492
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1624635492
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1624635492
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1624635492
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1624635492
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1624635492
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_54
timestamp 1624635492
transform 1 0 6072 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1624635492
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_78
timestamp 1624635492
transform 1 0 8280 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_66
timestamp 1624635492
transform 1 0 7176 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1624635492
transform 1 0 10212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1624635492
transform 1 0 9108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1624635492
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_111
timestamp 1624635492
transform 1 0 11316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_135
timestamp 1624635492
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_123
timestamp 1624635492
transform 1 0 12420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1624635492
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1624635492
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1624635492
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1624635492
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1624635492
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_58
timestamp 1624635492
transform 1 0 6440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_51
timestamp 1624635492
transform 1 0 5796 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1624635492
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_70
timestamp 1624635492
transform 1 0 7544 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1624635492
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_82
timestamp 1624635492
transform 1 0 8648 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_115
timestamp 1624635492
transform 1 0 11684 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_106
timestamp 1624635492
transform 1 0 10856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1624635492
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_127
timestamp 1624635492
transform 1 0 12788 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_17
timestamp 1624635492
transform 1 0 2668 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_11
timestamp 1624635492
transform 1 0 2116 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1624635492
transform 1 0 1380 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output391_A
timestamp 1624635492
transform 1 0 2484 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output391
timestamp 1624635492
transform -1 0 2116 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1624635492
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1624635492
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1624635492
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1624635492
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1624635492
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1624635492
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1624635492
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_99
timestamp 1624635492
transform 1 0 10212 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_95
timestamp 1624635492
transform 1 0 9844 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_87
timestamp 1624635492
transform 1 0 9108 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1624635492
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _155_
timestamp 1624635492
transform 1 0 9936 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_111
timestamp 1624635492
transform 1 0 11316 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_135
timestamp 1624635492
transform 1 0 13524 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_123
timestamp 1624635492
transform 1 0 12420 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1624635492
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1624635492
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1624635492
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1624635492
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1624635492
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1624635492
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1624635492
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1624635492
transform 1 0 3588 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1624635492
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1624635492
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1624635492
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1624635492
transform 1 0 6072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1624635492
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_58
timestamp 1624635492
transform 1 0 6440 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_51
timestamp 1624635492
transform 1 0 5796 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1624635492
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_78
timestamp 1624635492
transform 1 0 8280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1624635492
transform 1 0 7176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _347_
timestamp 1624635492
transform 1 0 6808 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_60_99
timestamp 1624635492
transform 1 0 10212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_87
timestamp 1624635492
transform 1 0 9108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1624635492
transform 1 0 9660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_87
timestamp 1624635492
transform 1 0 9108 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_81
timestamp 1624635492
transform 1 0 8556 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__CLK
timestamp 1624635492
transform -1 0 9660 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__D
timestamp 1624635492
transform -1 0 9108 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1624635492
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_111
timestamp 1624635492
transform 1 0 11316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_115
timestamp 1624635492
transform 1 0 11684 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_113
timestamp 1624635492
transform 1 0 11500 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_105
timestamp 1624635492
transform 1 0 10764 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1624635492
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1624635492
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1624635492
transform 1 0 12420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_127
timestamp 1624635492
transform 1 0 12788 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_17
timestamp 1624635492
transform 1 0 2668 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_11
timestamp 1624635492
transform 1 0 2116 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1624635492
transform 1 0 1380 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output429_A
timestamp 1624635492
transform -1 0 2668 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output429
timestamp 1624635492
transform -1 0 2116 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1624635492
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_29
timestamp 1624635492
transform 1 0 3772 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_58
timestamp 1624635492
transform 1 0 6440 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_53
timestamp 1624635492
transform 1 0 5980 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_41
timestamp 1624635492
transform 1 0 4876 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1624635492
transform 1 0 6348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_79
timestamp 1624635492
transform 1 0 8372 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_67
timestamp 1624635492
transform 1 0 7268 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _199_
timestamp 1624635492
transform 1 0 6992 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_91
timestamp 1624635492
transform 1 0 9476 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_115
timestamp 1624635492
transform 1 0 11684 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_111
timestamp 1624635492
transform 1 0 11316 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_103
timestamp 1624635492
transform 1 0 10580 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1624635492
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_127
timestamp 1624635492
transform 1 0 12788 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_15
timestamp 1624635492
transform 1 0 2484 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1624635492
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1624635492
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _279_
timestamp 1624635492
transform 1 0 2668 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1624635492
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_28
timestamp 1624635492
transform 1 0 3680 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1624635492
transform 1 0 2944 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1624635492
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_49
timestamp 1624635492
transform 1 0 5612 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_42
timestamp 1624635492
transform 1 0 4968 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _268_
timestamp 1624635492
transform 1 0 5336 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_73
timestamp 1624635492
transform 1 0 7820 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_61
timestamp 1624635492
transform 1 0 6716 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1624635492
transform 1 0 10212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_87
timestamp 1624635492
transform 1 0 9108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_85
timestamp 1624635492
transform 1 0 8924 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1624635492
transform 1 0 9016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_111
timestamp 1624635492
transform 1 0 11316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_135
timestamp 1624635492
transform 1 0 13524 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_123
timestamp 1624635492
transform 1 0 12420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_12
timestamp 1624635492
transform 1 0 2208 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_6
timestamp 1624635492
transform 1 0 1656 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 2208 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1624635492
transform -1 0 1656 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1624635492
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_36
timestamp 1624635492
transform 1 0 4416 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_24
timestamp 1624635492
transform 1 0 3312 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_58
timestamp 1624635492
transform 1 0 6440 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_56
timestamp 1624635492
transform 1 0 6256 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1624635492
transform 1 0 5520 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1624635492
transform 1 0 6348 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_70
timestamp 1624635492
transform 1 0 7544 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1624635492
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_82
timestamp 1624635492
transform 1 0 8648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_115
timestamp 1624635492
transform 1 0 11684 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_106
timestamp 1624635492
transform 1 0 10856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1624635492
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_127
timestamp 1624635492
transform 1 0 12788 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1624635492
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1624635492
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1624635492
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_30
timestamp 1624635492
transform 1 0 3864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_27
timestamp 1624635492
transform 1 0 3588 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1624635492
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_54
timestamp 1624635492
transform 1 0 6072 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_42
timestamp 1624635492
transform 1 0 4968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_78
timestamp 1624635492
transform 1 0 8280 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_66
timestamp 1624635492
transform 1 0 7176 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_99
timestamp 1624635492
transform 1 0 10212 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_87
timestamp 1624635492
transform 1 0 9108 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1624635492
transform 1 0 9016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_111
timestamp 1624635492
transform 1 0 11316 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_135
timestamp 1624635492
transform 1 0 13524 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_123
timestamp 1624635492
transform 1 0 12420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1624635492
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1624635492
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1624635492
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1624635492
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1624635492
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_58
timestamp 1624635492
transform 1 0 6440 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_51
timestamp 1624635492
transform 1 0 5796 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1624635492
transform 1 0 6348 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_70
timestamp 1624635492
transform 1 0 7544 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_94
timestamp 1624635492
transform 1 0 9752 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_82
timestamp 1624635492
transform 1 0 8648 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_115
timestamp 1624635492
transform 1 0 11684 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_106
timestamp 1624635492
transform 1 0 10856 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1624635492
transform 1 0 11592 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_127
timestamp 1624635492
transform 1 0 12788 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1624635492
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1624635492
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1624635492
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1624635492
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1624635492
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1624635492
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1624635492
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1624635492
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_30
timestamp 1624635492
transform 1 0 3864 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_27
timestamp 1624635492
transform 1 0 3588 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1624635492
transform 1 0 3772 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_58
timestamp 1624635492
transform 1 0 6440 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_51
timestamp 1624635492
transform 1 0 5796 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_54
timestamp 1624635492
transform 1 0 6072 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_42
timestamp 1624635492
transform 1 0 4968 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1624635492
transform 1 0 6348 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_70
timestamp 1624635492
transform 1 0 7544 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_78
timestamp 1624635492
transform 1 0 8280 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_66
timestamp 1624635492
transform 1 0 7176 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_94
timestamp 1624635492
transform 1 0 9752 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_82
timestamp 1624635492
transform 1 0 8648 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_99
timestamp 1624635492
transform 1 0 10212 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_87
timestamp 1624635492
transform 1 0 9108 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1624635492
transform 1 0 9016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_115
timestamp 1624635492
transform 1 0 11684 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_106
timestamp 1624635492
transform 1 0 10856 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_111
timestamp 1624635492
transform 1 0 11316 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1624635492
transform 1 0 11592 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_127
timestamp 1624635492
transform 1 0 12788 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_135
timestamp 1624635492
transform 1 0 13524 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_123
timestamp 1624635492
transform 1 0 12420 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_17
timestamp 1624635492
transform 1 0 2668 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_11
timestamp 1624635492
transform 1 0 2116 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1624635492
transform 1 0 1380 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output389_A
timestamp 1624635492
transform -1 0 2668 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output389
timestamp 1624635492
transform -1 0 2116 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1624635492
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_30
timestamp 1624635492
transform 1 0 3864 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1624635492
transform 1 0 3772 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_54
timestamp 1624635492
transform 1 0 6072 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_42
timestamp 1624635492
transform 1 0 4968 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_78
timestamp 1624635492
transform 1 0 8280 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_66
timestamp 1624635492
transform 1 0 7176 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_99
timestamp 1624635492
transform 1 0 10212 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_87
timestamp 1624635492
transform 1 0 9108 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1624635492
transform 1 0 9016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_111
timestamp 1624635492
transform 1 0 11316 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_135
timestamp 1624635492
transform 1 0 13524 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_123
timestamp 1624635492
transform 1 0 12420 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1624635492
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1624635492
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1624635492
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1624635492
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1624635492
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_58
timestamp 1624635492
transform 1 0 6440 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_51
timestamp 1624635492
transform 1 0 5796 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1624635492
transform 1 0 6348 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_70
timestamp 1624635492
transform 1 0 7544 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_94
timestamp 1624635492
transform 1 0 9752 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_82
timestamp 1624635492
transform 1 0 8648 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_115
timestamp 1624635492
transform 1 0 11684 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_106
timestamp 1624635492
transform 1 0 10856 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1624635492
transform 1 0 11592 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_127
timestamp 1624635492
transform 1 0 12788 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_17
timestamp 1624635492
transform 1 0 2668 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_11
timestamp 1624635492
transform 1 0 2116 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1624635492
transform 1 0 1380 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output427_A
timestamp 1624635492
transform 1 0 2484 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output427
timestamp 1624635492
transform -1 0 2116 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1624635492
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_30
timestamp 1624635492
transform 1 0 3864 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1624635492
transform 1 0 3772 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_54
timestamp 1624635492
transform 1 0 6072 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_42
timestamp 1624635492
transform 1 0 4968 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_78
timestamp 1624635492
transform 1 0 8280 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_66
timestamp 1624635492
transform 1 0 7176 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_99
timestamp 1624635492
transform 1 0 10212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_87
timestamp 1624635492
transform 1 0 9108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1624635492
transform 1 0 9016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_111
timestamp 1624635492
transform 1 0 11316 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_135
timestamp 1624635492
transform 1 0 13524 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_123
timestamp 1624635492
transform 1 0 12420 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1624635492
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1624635492
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1624635492
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1624635492
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1624635492
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_58
timestamp 1624635492
transform 1 0 6440 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_51
timestamp 1624635492
transform 1 0 5796 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1624635492
transform 1 0 6348 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_70
timestamp 1624635492
transform 1 0 7544 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_94
timestamp 1624635492
transform 1 0 9752 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_82
timestamp 1624635492
transform 1 0 8648 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_115
timestamp 1624635492
transform 1 0 11684 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_106
timestamp 1624635492
transform 1 0 10856 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1624635492
transform 1 0 11592 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_127
timestamp 1624635492
transform 1 0 12788 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_12
timestamp 1624635492
transform 1 0 2208 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_6
timestamp 1624635492
transform 1 0 1656 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1624635492
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1624635492
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 2208 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform -1 0 1656 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1624635492
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1624635492
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_36
timestamp 1624635492
transform 1 0 4416 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_24
timestamp 1624635492
transform 1 0 3312 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_30
timestamp 1624635492
transform 1 0 3864 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_27
timestamp 1624635492
transform 1 0 3588 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1624635492
transform 1 0 3772 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_58
timestamp 1624635492
transform 1 0 6440 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_56
timestamp 1624635492
transform 1 0 6256 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_48
timestamp 1624635492
transform 1 0 5520 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_54
timestamp 1624635492
transform 1 0 6072 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_42
timestamp 1624635492
transform 1 0 4968 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1624635492
transform 1 0 6348 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_70
timestamp 1624635492
transform 1 0 7544 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_78
timestamp 1624635492
transform 1 0 8280 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_66
timestamp 1624635492
transform 1 0 7176 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_94
timestamp 1624635492
transform 1 0 9752 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_82
timestamp 1624635492
transform 1 0 8648 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_99
timestamp 1624635492
transform 1 0 10212 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_87
timestamp 1624635492
transform 1 0 9108 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1624635492
transform 1 0 9016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_115
timestamp 1624635492
transform 1 0 11684 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_106
timestamp 1624635492
transform 1 0 10856 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_111
timestamp 1624635492
transform 1 0 11316 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1624635492
transform 1 0 11592 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_127
timestamp 1624635492
transform 1 0 12788 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_135
timestamp 1624635492
transform 1 0 13524 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_123
timestamp 1624635492
transform 1 0 12420 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1624635492
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1624635492
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1624635492
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_30
timestamp 1624635492
transform 1 0 3864 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_27
timestamp 1624635492
transform 1 0 3588 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1624635492
transform 1 0 3772 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_54
timestamp 1624635492
transform 1 0 6072 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_42
timestamp 1624635492
transform 1 0 4968 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_78
timestamp 1624635492
transform 1 0 8280 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_66
timestamp 1624635492
transform 1 0 7176 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_99
timestamp 1624635492
transform 1 0 10212 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_87
timestamp 1624635492
transform 1 0 9108 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1624635492
transform 1 0 9016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_118
timestamp 1624635492
transform 1 0 11960 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_111
timestamp 1624635492
transform 1 0 11316 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _311_
timestamp 1624635492
transform -1 0 11960 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_128
timestamp 1624635492
transform 1 0 12880 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_124
timestamp 1624635492
transform 1 0 12512 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _239_
timestamp 1624635492
transform 1 0 12604 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1624635492
transform 1 0 1380 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1624635492
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _345_
timestamp 1624635492
transform -1 0 3312 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_36
timestamp 1624635492
transform 1 0 4416 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_30
timestamp 1624635492
transform 1 0 3864 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_24
timestamp 1624635492
transform 1 0 3312 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__CLK
timestamp 1624635492
transform 1 0 4232 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__D
timestamp 1624635492
transform 1 0 3680 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_58
timestamp 1624635492
transform 1 0 6440 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_56
timestamp 1624635492
transform 1 0 6256 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_48
timestamp 1624635492
transform 1 0 5520 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1624635492
transform 1 0 6348 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_70
timestamp 1624635492
transform 1 0 7544 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_94
timestamp 1624635492
transform 1 0 9752 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_82
timestamp 1624635492
transform 1 0 8648 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_115
timestamp 1624635492
transform 1 0 11684 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_106
timestamp 1624635492
transform 1 0 10856 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1624635492
transform 1 0 11592 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_132
timestamp 1624635492
transform 1 0 13248 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_127
timestamp 1624635492
transform 1 0 12788 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1624635492
transform 1 0 13616 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1624635492
transform 1 0 12972 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1624635492
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1624635492
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1624635492
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_30
timestamp 1624635492
transform 1 0 3864 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_27
timestamp 1624635492
transform 1 0 3588 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1624635492
transform 1 0 3772 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_54
timestamp 1624635492
transform 1 0 6072 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_42
timestamp 1624635492
transform 1 0 4968 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_78
timestamp 1624635492
transform 1 0 8280 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_66
timestamp 1624635492
transform 1 0 7176 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_99
timestamp 1624635492
transform 1 0 10212 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_87
timestamp 1624635492
transform 1 0 9108 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1624635492
transform 1 0 9016 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_111
timestamp 1624635492
transform 1 0 11316 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_135
timestamp 1624635492
transform 1 0 13524 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_123
timestamp 1624635492
transform 1 0 12420 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1624635492
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1624635492
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1624635492
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1624635492
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1624635492
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_58
timestamp 1624635492
transform 1 0 6440 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_51
timestamp 1624635492
transform 1 0 5796 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1624635492
transform 1 0 6348 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_70
timestamp 1624635492
transform 1 0 7544 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_94
timestamp 1624635492
transform 1 0 9752 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_82
timestamp 1624635492
transform 1 0 8648 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_115
timestamp 1624635492
transform 1 0 11684 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_113
timestamp 1624635492
transform 1 0 11500 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_107
timestamp 1624635492
transform 1 0 10948 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_102
timestamp 1624635492
transform 1 0 10488 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1624635492
transform 1 0 11592 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _316_
timestamp 1624635492
transform -1 0 10948 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_127
timestamp 1624635492
transform 1 0 12788 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_17
timestamp 1624635492
transform 1 0 2668 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_11
timestamp 1624635492
transform 1 0 2116 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1624635492
transform 1 0 1380 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output388_A
timestamp 1624635492
transform -1 0 2668 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output388
timestamp 1624635492
transform -1 0 2116 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1624635492
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_30
timestamp 1624635492
transform 1 0 3864 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1624635492
transform 1 0 3772 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_54
timestamp 1624635492
transform 1 0 6072 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_42
timestamp 1624635492
transform 1 0 4968 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_78
timestamp 1624635492
transform 1 0 8280 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_66
timestamp 1624635492
transform 1 0 7176 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_99
timestamp 1624635492
transform 1 0 10212 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_87
timestamp 1624635492
transform 1 0 9108 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1624635492
transform 1 0 9016 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_111
timestamp 1624635492
transform 1 0 11316 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_135
timestamp 1624635492
transform 1 0 13524 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_123
timestamp 1624635492
transform 1 0 12420 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1624635492
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1624635492
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1624635492
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1624635492
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1624635492
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_58
timestamp 1624635492
transform 1 0 6440 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_51
timestamp 1624635492
transform 1 0 5796 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1624635492
transform 1 0 6348 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_70
timestamp 1624635492
transform 1 0 7544 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_94
timestamp 1624635492
transform 1 0 9752 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_82
timestamp 1624635492
transform 1 0 8648 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_115
timestamp 1624635492
transform 1 0 11684 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_106
timestamp 1624635492
transform 1 0 10856 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1624635492
transform 1 0 11592 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_130
timestamp 1624635492
transform 1 0 13064 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _152_
timestamp 1624635492
transform 1 0 12788 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1624635492
transform 1 0 14352 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1624635492
transform 1 0 14996 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_139
timestamp 1624635492
transform 1 0 13892 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1624635492
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_168
timestamp 1624635492
transform 1 0 16560 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_156
timestamp 1624635492
transform 1 0 15456 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1624635492
transform 1 0 16928 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_163
timestamp 1624635492
transform 1 0 16100 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1624635492
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_180
timestamp 1624635492
transform 1 0 17664 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1624635492
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_201
timestamp 1624635492
transform 1 0 19596 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_192
timestamp 1624635492
transform 1 0 18768 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1624635492
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1624635492
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_225
timestamp 1624635492
transform 1 0 21804 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_213
timestamp 1624635492
transform 1 0 20700 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_220
timestamp 1624635492
transform 1 0 21344 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1624635492
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_237
timestamp 1624635492
transform 1 0 22908 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_241
timestamp 1624635492
transform 1 0 23276 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_229
timestamp 1624635492
transform 1 0 22172 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1624635492
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_258
timestamp 1624635492
transform 1 0 24840 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_249
timestamp 1624635492
transform 1 0 24012 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_253
timestamp 1624635492
transform 1 0 24380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1624635492
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_270
timestamp 1624635492
transform 1 0 25944 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1624635492
transform 1 0 25484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_151
timestamp 1624635492
transform 1 0 14996 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_139
timestamp 1624635492
transform 1 0 13892 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1624635492
transform 1 0 16928 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_163
timestamp 1624635492
transform 1 0 16100 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1624635492
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1624635492
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1624635492
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_220
timestamp 1624635492
transform 1 0 21344 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1624635492
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_241
timestamp 1624635492
transform 1 0 23276 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_229
timestamp 1624635492
transform 1 0 22172 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1624635492
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_253
timestamp 1624635492
transform 1 0 24380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_265
timestamp 1624635492
transform 1 0 25484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_144
timestamp 1624635492
transform 1 0 14352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1624635492
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1624635492
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_156
timestamp 1624635492
transform 1 0 15456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1624635492
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_201
timestamp 1624635492
transform 1 0 19596 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_192
timestamp 1624635492
transform 1 0 18768 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1624635492
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_225
timestamp 1624635492
transform 1 0 21804 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_213
timestamp 1624635492
transform 1 0 20700 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_237
timestamp 1624635492
transform 1 0 22908 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1624635492
transform 1 0 24840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_249
timestamp 1624635492
transform 1 0 24012 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1624635492
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1624635492
transform 1 0 25944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1624635492
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_139
timestamp 1624635492
transform 1 0 13892 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1624635492
transform 1 0 16928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_163
timestamp 1624635492
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1624635492
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1624635492
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1624635492
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_220
timestamp 1624635492
transform 1 0 21344 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1624635492
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_241
timestamp 1624635492
transform 1 0 23276 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_229
timestamp 1624635492
transform 1 0 22172 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1624635492
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_253
timestamp 1624635492
transform 1 0 24380 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _264_
timestamp 1624635492
transform 1 0 24932 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_262
timestamp 1624635492
transform 1 0 25208 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1624635492
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1624635492
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1624635492
transform 1 0 16560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1624635492
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_180
timestamp 1624635492
transform 1 0 17664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1624635492
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_192
timestamp 1624635492
transform 1 0 18768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1624635492
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_225
timestamp 1624635492
transform 1 0 21804 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_213
timestamp 1624635492
transform 1 0 20700 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_237
timestamp 1624635492
transform 1 0 22908 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1624635492
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_249
timestamp 1624635492
transform 1 0 24012 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1624635492
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1624635492
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_144
timestamp 1624635492
transform 1 0 14352 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1624635492
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_139
timestamp 1624635492
transform 1 0 13892 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1624635492
transform 1 0 14260 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_168
timestamp 1624635492
transform 1 0 16560 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_156
timestamp 1624635492
transform 1 0 15456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1624635492
transform 1 0 16928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_163
timestamp 1624635492
transform 1 0 16100 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1624635492
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_180
timestamp 1624635492
transform 1 0 17664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1624635492
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_201
timestamp 1624635492
transform 1 0 19596 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_192
timestamp 1624635492
transform 1 0 18768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1624635492
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1624635492
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_225
timestamp 1624635492
transform 1 0 21804 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_213
timestamp 1624635492
transform 1 0 20700 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_220
timestamp 1624635492
transform 1 0 21344 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1624635492
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_237
timestamp 1624635492
transform 1 0 22908 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_241
timestamp 1624635492
transform 1 0 23276 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_229
timestamp 1624635492
transform 1 0 22172 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1624635492
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1624635492
transform 1 0 24840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_249
timestamp 1624635492
transform 1 0 24012 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_253
timestamp 1624635492
transform 1 0 24380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1624635492
transform 1 0 24748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_270
timestamp 1624635492
transform 1 0 25944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_265
timestamp 1624635492
transform 1 0 25484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_151
timestamp 1624635492
transform 1 0 14996 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_139
timestamp 1624635492
transform 1 0 13892 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_172
timestamp 1624635492
transform 1 0 16928 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_163
timestamp 1624635492
transform 1 0 16100 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1624635492
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1624635492
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1624635492
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_220
timestamp 1624635492
transform 1 0 21344 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1624635492
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_241
timestamp 1624635492
transform 1 0 23276 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_229
timestamp 1624635492
transform 1 0 22172 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1624635492
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_253
timestamp 1624635492
transform 1 0 24380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_265
timestamp 1624635492
transform 1 0 25484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1624635492
transform 1 0 14352 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1624635492
transform 1 0 14260 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1624635492
transform 1 0 16560 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_156
timestamp 1624635492
transform 1 0 15456 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_180
timestamp 1624635492
transform 1 0 17664 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1624635492
transform 1 0 19596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_192
timestamp 1624635492
transform 1 0 18768 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1624635492
transform 1 0 19504 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1624635492
transform 1 0 21804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_213
timestamp 1624635492
transform 1 0 20700 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1624635492
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1624635492
transform 1 0 24840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1624635492
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1624635492
transform 1 0 24748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_270
timestamp 1624635492
transform 1 0 25944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_151
timestamp 1624635492
transform 1 0 14996 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_139
timestamp 1624635492
transform 1 0 13892 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_172
timestamp 1624635492
transform 1 0 16928 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_163
timestamp 1624635492
transform 1 0 16100 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1624635492
transform 1 0 16836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1624635492
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1624635492
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_220
timestamp 1624635492
transform 1 0 21344 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1624635492
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1624635492
transform 1 0 23276 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1624635492
transform 1 0 22172 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1624635492
transform 1 0 22080 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1624635492
transform 1 0 24380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_265
timestamp 1624635492
transform 1 0 25484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_144
timestamp 1624635492
transform 1 0 14352 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1624635492
transform 1 0 14260 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_168
timestamp 1624635492
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_156
timestamp 1624635492
transform 1 0 15456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_180
timestamp 1624635492
transform 1 0 17664 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_201
timestamp 1624635492
transform 1 0 19596 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_192
timestamp 1624635492
transform 1 0 18768 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1624635492
transform 1 0 19504 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1624635492
transform 1 0 21804 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_213
timestamp 1624635492
transform 1 0 20700 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_237
timestamp 1624635492
transform 1 0 22908 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_258
timestamp 1624635492
transform 1 0 24840 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_249
timestamp 1624635492
transform 1 0 24012 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1624635492
transform 1 0 24748 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_270
timestamp 1624635492
transform 1 0 25944 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_151
timestamp 1624635492
transform 1 0 14996 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_139
timestamp 1624635492
transform 1 0 13892 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_172
timestamp 1624635492
transform 1 0 16928 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_163
timestamp 1624635492
transform 1 0 16100 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1624635492
transform 1 0 16836 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1624635492
transform 1 0 18032 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_196
timestamp 1624635492
transform 1 0 19136 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_220
timestamp 1624635492
transform 1 0 21344 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_208
timestamp 1624635492
transform 1 0 20240 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_241
timestamp 1624635492
transform 1 0 23276 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_229
timestamp 1624635492
transform 1 0 22172 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1624635492
transform 1 0 22080 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_253
timestamp 1624635492
transform 1 0 24380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_265
timestamp 1624635492
transform 1 0 25484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_151
timestamp 1624635492
transform 1 0 14996 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_139
timestamp 1624635492
transform 1 0 13892 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_144
timestamp 1624635492
transform 1 0 14352 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1624635492
transform 1 0 14260 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_172
timestamp 1624635492
transform 1 0 16928 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_163
timestamp 1624635492
transform 1 0 16100 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_168
timestamp 1624635492
transform 1 0 16560 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_156
timestamp 1624635492
transform 1 0 15456 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1624635492
transform 1 0 16836 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1624635492
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_180
timestamp 1624635492
transform 1 0 17664 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_196
timestamp 1624635492
transform 1 0 19136 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_201
timestamp 1624635492
transform 1 0 19596 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_192
timestamp 1624635492
transform 1 0 18768 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1624635492
transform 1 0 19504 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_220
timestamp 1624635492
transform 1 0 21344 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_208
timestamp 1624635492
transform 1 0 20240 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_225
timestamp 1624635492
transform 1 0 21804 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_213
timestamp 1624635492
transform 1 0 20700 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_241
timestamp 1624635492
transform 1 0 23276 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_229
timestamp 1624635492
transform 1 0 22172 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_237
timestamp 1624635492
transform 1 0 22908 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1624635492
transform 1 0 22080 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_253
timestamp 1624635492
transform 1 0 24380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_258
timestamp 1624635492
transform 1 0 24840 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_249
timestamp 1624635492
transform 1 0 24012 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1624635492
transform 1 0 24748 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_265
timestamp 1624635492
transform 1 0 25484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_270
timestamp 1624635492
transform 1 0 25944 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_144
timestamp 1624635492
transform 1 0 14352 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1624635492
transform 1 0 14260 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_168
timestamp 1624635492
transform 1 0 16560 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_156
timestamp 1624635492
transform 1 0 15456 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_180
timestamp 1624635492
transform 1 0 17664 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_201
timestamp 1624635492
transform 1 0 19596 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_192
timestamp 1624635492
transform 1 0 18768 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1624635492
transform 1 0 19504 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_225
timestamp 1624635492
transform 1 0 21804 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_213
timestamp 1624635492
transform 1 0 20700 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_237
timestamp 1624635492
transform 1 0 22908 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_258
timestamp 1624635492
transform 1 0 24840 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_249
timestamp 1624635492
transform 1 0 24012 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1624635492
transform 1 0 24748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_270
timestamp 1624635492
transform 1 0 25944 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_151
timestamp 1624635492
transform 1 0 14996 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_139
timestamp 1624635492
transform 1 0 13892 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_172
timestamp 1624635492
transform 1 0 16928 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_163
timestamp 1624635492
transform 1 0 16100 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1624635492
transform 1 0 16836 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_184
timestamp 1624635492
transform 1 0 18032 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_196
timestamp 1624635492
transform 1 0 19136 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_220
timestamp 1624635492
transform 1 0 21344 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_208
timestamp 1624635492
transform 1 0 20240 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_241
timestamp 1624635492
transform 1 0 23276 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_229
timestamp 1624635492
transform 1 0 22172 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1624635492
transform 1 0 22080 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_253
timestamp 1624635492
transform 1 0 24380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_265
timestamp 1624635492
transform 1 0 25484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_144
timestamp 1624635492
transform 1 0 14352 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1624635492
transform 1 0 14260 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_168
timestamp 1624635492
transform 1 0 16560 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_156
timestamp 1624635492
transform 1 0 15456 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_180
timestamp 1624635492
transform 1 0 17664 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_201
timestamp 1624635492
transform 1 0 19596 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_192
timestamp 1624635492
transform 1 0 18768 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1624635492
transform 1 0 19504 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_225
timestamp 1624635492
transform 1 0 21804 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_213
timestamp 1624635492
transform 1 0 20700 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_240
timestamp 1624635492
transform 1 0 23184 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1624635492
transform 1 0 22908 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_258
timestamp 1624635492
transform 1 0 24840 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_254
timestamp 1624635492
transform 1 0 24472 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_246
timestamp 1624635492
transform 1 0 23736 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1624635492
transform 1 0 23552 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1624635492
transform 1 0 24748 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_270
timestamp 1624635492
transform 1 0 25944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_151
timestamp 1624635492
transform 1 0 14996 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_139
timestamp 1624635492
transform 1 0 13892 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_172
timestamp 1624635492
transform 1 0 16928 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_163
timestamp 1624635492
transform 1 0 16100 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1624635492
transform 1 0 16836 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_187
timestamp 1624635492
transform 1 0 18308 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_179
timestamp 1624635492
transform 1 0 17572 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_176
timestamp 1624635492
transform 1 0 17296 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__A1
timestamp 1624635492
transform 1 0 17388 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__B2
timestamp 1624635492
transform 1 0 18492 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_203
timestamp 1624635492
transform 1 0 19780 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_191
timestamp 1624635492
transform 1 0 18676 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_215
timestamp 1624635492
transform 1 0 20884 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_241
timestamp 1624635492
transform 1 0 23276 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_229
timestamp 1624635492
transform 1 0 22172 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_227
timestamp 1624635492
transform 1 0 21988 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1624635492
transform 1 0 22080 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_253
timestamp 1624635492
transform 1 0 24380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_265
timestamp 1624635492
transform 1 0 25484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_151
timestamp 1624635492
transform 1 0 14996 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_139
timestamp 1624635492
transform 1 0 13892 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_144
timestamp 1624635492
transform 1 0 14352 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1624635492
transform 1 0 14260 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_172
timestamp 1624635492
transform 1 0 16928 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_163
timestamp 1624635492
transform 1 0 16100 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_72_172
timestamp 1624635492
transform 1 0 16928 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_163
timestamp 1624635492
transform 1 0 16100 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_156
timestamp 1624635492
transform 1 0 15456 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1624635492
transform 1 0 16836 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _320_
timestamp 1624635492
transform -1 0 16928 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _255_
timestamp 1624635492
transform 1 0 15824 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_190
timestamp 1624635492
transform 1 0 18584 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_184
timestamp 1624635492
transform 1 0 18032 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_187
timestamp 1624635492
transform 1 0 18308 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_178
timestamp 1624635492
transform 1 0 17480 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _055_
timestamp 1624635492
transform -1 0 18308 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1624635492
transform 1 0 19964 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1624635492
transform 1 0 18860 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_201
timestamp 1624635492
transform 1 0 19596 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_199
timestamp 1624635492
transform 1 0 19412 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_193
timestamp 1624635492
transform 1 0 18860 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__B1
timestamp 1624635492
transform 1 0 18676 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__A2
timestamp 1624635492
transform 1 0 18676 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1624635492
transform 1 0 19504 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_225
timestamp 1624635492
transform 1 0 21804 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_217
timestamp 1624635492
transform 1 0 21068 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_225
timestamp 1624635492
transform 1 0 21804 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_213
timestamp 1624635492
transform 1 0 20700 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_241
timestamp 1624635492
transform 1 0 23276 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_229
timestamp 1624635492
transform 1 0 22172 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_237
timestamp 1624635492
transform 1 0 22908 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1624635492
transform 1 0 22080 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_253
timestamp 1624635492
transform 1 0 24380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_258
timestamp 1624635492
transform 1 0 24840 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_249
timestamp 1624635492
transform 1 0 24012 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1624635492
transform 1 0 24748 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_273
timestamp 1624635492
transform 1 0 26220 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_265
timestamp 1624635492
transform 1 0 25484 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_270
timestamp 1624635492
transform 1 0 25944 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_144
timestamp 1624635492
transform 1 0 14352 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_140
timestamp 1624635492
transform 1 0 13984 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1624635492
transform 1 0 14260 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_168
timestamp 1624635492
transform 1 0 16560 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_156
timestamp 1624635492
transform 1 0 15456 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_180
timestamp 1624635492
transform 1 0 17664 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_201
timestamp 1624635492
transform 1 0 19596 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_192
timestamp 1624635492
transform 1 0 18768 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1624635492
transform 1 0 19504 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _275_
timestamp 1624635492
transform 1 0 19964 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_220
timestamp 1624635492
transform 1 0 21344 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_208
timestamp 1624635492
transform 1 0 20240 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_232
timestamp 1624635492
transform 1 0 22448 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_258
timestamp 1624635492
transform 1 0 24840 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_256
timestamp 1624635492
transform 1 0 24656 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_244
timestamp 1624635492
transform 1 0 23552 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1624635492
transform 1 0 24748 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_270
timestamp 1624635492
transform 1 0 25944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_150
timestamp 1624635492
transform 1 0 14904 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_138
timestamp 1624635492
transform 1 0 13800 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_172
timestamp 1624635492
transform 1 0 16928 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_170
timestamp 1624635492
transform 1 0 16744 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_162
timestamp 1624635492
transform 1 0 16008 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1624635492
transform 1 0 16836 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_184
timestamp 1624635492
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_196
timestamp 1624635492
transform 1 0 19136 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_220
timestamp 1624635492
transform 1 0 21344 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_208
timestamp 1624635492
transform 1 0 20240 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_241
timestamp 1624635492
transform 1 0 23276 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_229
timestamp 1624635492
transform 1 0 22172 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1624635492
transform 1 0 22080 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_253
timestamp 1624635492
transform 1 0 24380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_265
timestamp 1624635492
transform 1 0 25484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_144
timestamp 1624635492
transform 1 0 14352 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1624635492
transform 1 0 14260 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_168
timestamp 1624635492
transform 1 0 16560 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_156
timestamp 1624635492
transform 1 0 15456 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_180
timestamp 1624635492
transform 1 0 17664 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_201
timestamp 1624635492
transform 1 0 19596 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_192
timestamp 1624635492
transform 1 0 18768 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1624635492
transform 1 0 19504 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_225
timestamp 1624635492
transform 1 0 21804 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_213
timestamp 1624635492
transform 1 0 20700 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_237
timestamp 1624635492
transform 1 0 22908 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_258
timestamp 1624635492
transform 1 0 24840 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_249
timestamp 1624635492
transform 1 0 24012 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1624635492
transform 1 0 24748 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_270
timestamp 1624635492
transform 1 0 25944 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_151
timestamp 1624635492
transform 1 0 14996 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_139
timestamp 1624635492
transform 1 0 13892 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_172
timestamp 1624635492
transform 1 0 16928 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_163
timestamp 1624635492
transform 1 0 16100 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1624635492
transform 1 0 16836 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_184
timestamp 1624635492
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_196
timestamp 1624635492
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_220
timestamp 1624635492
transform 1 0 21344 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_208
timestamp 1624635492
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_241
timestamp 1624635492
transform 1 0 23276 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_229
timestamp 1624635492
transform 1 0 22172 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1624635492
transform 1 0 22080 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_253
timestamp 1624635492
transform 1 0 24380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_265
timestamp 1624635492
transform 1 0 25484 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_152
timestamp 1624635492
transform 1 0 15088 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_144
timestamp 1624635492
transform 1 0 14352 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__D
timestamp 1624635492
transform 1 0 15272 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1624635492
transform 1 0 14260 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_156
timestamp 1624635492
transform 1 0 15456 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _342_
timestamp 1624635492
transform -1 0 17388 0 -1 45152
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_78_183
timestamp 1624635492
transform 1 0 17940 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_177
timestamp 1624635492
transform 1 0 17388 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__CLK
timestamp 1624635492
transform 1 0 17756 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_201
timestamp 1624635492
transform 1 0 19596 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_199
timestamp 1624635492
transform 1 0 19412 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_195
timestamp 1624635492
transform 1 0 19044 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1624635492
transform 1 0 19504 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_225
timestamp 1624635492
transform 1 0 21804 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_213
timestamp 1624635492
transform 1 0 20700 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_237
timestamp 1624635492
transform 1 0 22908 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_258
timestamp 1624635492
transform 1 0 24840 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_249
timestamp 1624635492
transform 1 0 24012 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1624635492
transform 1 0 24748 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_270
timestamp 1624635492
transform 1 0 25944 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_154
timestamp 1624635492
transform 1 0 15272 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_142
timestamp 1624635492
transform 1 0 14168 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_172
timestamp 1624635492
transform 1 0 16928 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_170
timestamp 1624635492
transform 1 0 16744 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_166
timestamp 1624635492
transform 1 0 16376 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1624635492
transform 1 0 16836 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_184
timestamp 1624635492
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_196
timestamp 1624635492
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_220
timestamp 1624635492
transform 1 0 21344 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_208
timestamp 1624635492
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_241
timestamp 1624635492
transform 1 0 23276 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_229
timestamp 1624635492
transform 1 0 22172 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1624635492
transform 1 0 22080 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_253
timestamp 1624635492
transform 1 0 24380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_265
timestamp 1624635492
transform 1 0 25484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_288
timestamp 1624635492
transform 1 0 27600 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_281
timestamp 1624635492
transform 1 0 26956 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_286
timestamp 1624635492
transform 1 0 27416 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1624635492
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1624635492
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _190_
timestamp 1624635492
transform 1 0 27324 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _117_
timestamp 1624635492
transform 1 0 26680 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_312
timestamp 1624635492
transform 1 0 29808 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_300
timestamp 1624635492
transform 1 0 28704 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_310
timestamp 1624635492
transform 1 0 29624 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_298
timestamp 1624635492
transform 1 0 28520 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1624635492
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_327
timestamp 1624635492
transform 1 0 31188 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1624635492
transform 1 0 30084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_334
timestamp 1624635492
transform 1 0 31832 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_322
timestamp 1624635492
transform 1 0 30728 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_351
timestamp 1624635492
transform 1 0 33396 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_339
timestamp 1624635492
transform 1 0 32292 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1624635492
transform 1 0 33764 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1624635492
transform 1 0 32660 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1624635492
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_372
timestamp 1624635492
transform 1 0 35328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_363
timestamp 1624635492
transform 1 0 34500 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1624635492
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1624635492
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_388
timestamp 1624635492
transform 1 0 36800 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_384
timestamp 1624635492
transform 1 0 36432 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_398
timestamp 1624635492
transform 1 0 37720 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_390
timestamp 1624635492
transform 1 0 36984 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_387
timestamp 1624635492
transform 1 0 36708 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_379
timestamp 1624635492
transform 1 0 35972 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A3
timestamp 1624635492
transform 1 0 36800 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A2
timestamp 1624635492
transform 1 0 36616 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_2  _087_
timestamp 1624635492
transform 1 0 37168 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_54_407
timestamp 1624635492
transform 1 0 38548 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_401
timestamp 1624635492
transform 1 0 37996 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_400
timestamp 1624635492
transform 1 0 37904 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B1
timestamp 1624635492
transform 1 0 38364 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1624635492
transform 1 0 37812 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1624635492
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_277
timestamp 1624635492
transform 1 0 26588 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1624635492
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_310
timestamp 1624635492
transform 1 0 29624 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_298
timestamp 1624635492
transform 1 0 28520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_334
timestamp 1624635492
transform 1 0 31832 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1624635492
transform 1 0 30728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1624635492
transform 1 0 33764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1624635492
transform 1 0 32660 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1624635492
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1624635492
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_391
timestamp 1624635492
transform 1 0 37076 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1624635492
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_400
timestamp 1624635492
transform 1 0 37904 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1624635492
transform 1 0 37812 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1624635492
transform 1 0 27048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_306
timestamp 1624635492
transform 1 0 29256 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1624635492
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1624635492
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1624635492
transform 1 0 31188 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1624635492
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_351
timestamp 1624635492
transform 1 0 33396 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_339
timestamp 1624635492
transform 1 0 32292 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_372
timestamp 1624635492
transform 1 0 35328 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_363
timestamp 1624635492
transform 1 0 34500 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1624635492
transform 1 0 35236 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_396
timestamp 1624635492
transform 1 0 37536 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1624635492
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_408
timestamp 1624635492
transform 1 0 38640 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_286
timestamp 1624635492
transform 1 0 27416 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_282
timestamp 1624635492
transform 1 0 27048 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_274
timestamp 1624635492
transform 1 0 26312 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1624635492
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_310
timestamp 1624635492
transform 1 0 29624 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_298
timestamp 1624635492
transform 1 0 28520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_334
timestamp 1624635492
transform 1 0 31832 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1624635492
transform 1 0 30728 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_355
timestamp 1624635492
transform 1 0 33764 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1624635492
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1624635492
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1624635492
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_398
timestamp 1624635492
transform 1 0 37720 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_390
timestamp 1624635492
transform 1 0 36984 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_379
timestamp 1624635492
transform 1 0 35972 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _149_
timestamp 1624635492
transform 1 0 36708 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_400
timestamp 1624635492
transform 1 0 37904 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1624635492
transform 1 0 37812 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_282
timestamp 1624635492
transform 1 0 27048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_306
timestamp 1624635492
transform 1 0 29256 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1624635492
transform 1 0 28152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1624635492
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1624635492
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1624635492
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_347
timestamp 1624635492
transform 1 0 33028 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_341
timestamp 1624635492
transform 1 0 32476 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A1
timestamp 1624635492
transform -1 0 32476 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A2
timestamp 1624635492
transform 1 0 32844 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_372
timestamp 1624635492
transform 1 0 35328 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_359
timestamp 1624635492
transform 1 0 34132 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1624635492
transform 1 0 35236 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_396
timestamp 1624635492
transform 1 0 37536 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_384
timestamp 1624635492
transform 1 0 36432 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_408
timestamp 1624635492
transform 1 0 38640 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_282
timestamp 1624635492
transform 1 0 27048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1624635492
transform 1 0 27416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_277
timestamp 1624635492
transform 1 0 26588 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1624635492
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_306
timestamp 1624635492
transform 1 0 29256 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1624635492
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_314
timestamp 1624635492
transform 1 0 29992 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_310
timestamp 1624635492
transform 1 0 29624 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_298
timestamp 1624635492
transform 1 0 28520 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1624635492
transform 1 0 29992 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_326
timestamp 1624635492
transform 1 0 31096 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_323
timestamp 1624635492
transform 1 0 30820 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_315
timestamp 1624635492
transform 1 0 30084 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_330
timestamp 1624635492
transform 1 0 31464 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_318
timestamp 1624635492
transform 1 0 30360 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1624635492
transform 1 0 30912 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 31464 0 -1 35360
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _110_
timestamp 1624635492
transform 1 0 30084 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_350
timestamp 1624635492
transform 1 0 33304 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_356
timestamp 1624635492
transform 1 0 33856 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_343
timestamp 1624635492
transform 1 0 32660 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_338
timestamp 1624635492
transform 1 0 32200 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A3
timestamp 1624635492
transform 1 0 32016 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1624635492
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_2  _084_
timestamp 1624635492
transform 1 0 33028 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1624635492
transform 1 0 35328 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_370
timestamp 1624635492
transform 1 0 35144 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_362
timestamp 1624635492
transform 1 0 34408 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_368
timestamp 1624635492
transform 1 0 34960 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_362
timestamp 1624635492
transform 1 0 34408 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__C1
timestamp 1624635492
transform 1 0 34776 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B1
timestamp 1624635492
transform 1 0 34224 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1624635492
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_396
timestamp 1624635492
transform 1 0 37536 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_384
timestamp 1624635492
transform 1 0 36432 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_398
timestamp 1624635492
transform 1 0 37720 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_392
timestamp 1624635492
transform 1 0 37168 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_380
timestamp 1624635492
transform 1 0 36064 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_408
timestamp 1624635492
transform 1 0 38640 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_400
timestamp 1624635492
transform 1 0 37904 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1624635492
transform 1 0 37812 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1624635492
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_277
timestamp 1624635492
transform 1 0 26588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1624635492
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_310
timestamp 1624635492
transform 1 0 29624 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_298
timestamp 1624635492
transform 1 0 28520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_334
timestamp 1624635492
transform 1 0 31832 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_322
timestamp 1624635492
transform 1 0 30728 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_355
timestamp 1624635492
transform 1 0 33764 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_343
timestamp 1624635492
transform 1 0 32660 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1624635492
transform 1 0 32568 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1624635492
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_391
timestamp 1624635492
transform 1 0 37076 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1624635492
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_400
timestamp 1624635492
transform 1 0 37904 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1624635492
transform 1 0 37812 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_282
timestamp 1624635492
transform 1 0 27048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_306
timestamp 1624635492
transform 1 0 29256 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_294
timestamp 1624635492
transform 1 0 28152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1624635492
transform 1 0 29992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1624635492
transform 1 0 31188 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1624635492
transform 1 0 30084 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1624635492
transform 1 0 33396 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1624635492
transform 1 0 32292 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_372
timestamp 1624635492
transform 1 0 35328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_363
timestamp 1624635492
transform 1 0 34500 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1624635492
transform 1 0 35236 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_396
timestamp 1624635492
transform 1 0 37536 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_384
timestamp 1624635492
transform 1 0 36432 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_408
timestamp 1624635492
transform 1 0 38640 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_286
timestamp 1624635492
transform 1 0 27416 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_277
timestamp 1624635492
transform 1 0 26588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1624635492
transform 1 0 27324 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_310
timestamp 1624635492
transform 1 0 29624 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_298
timestamp 1624635492
transform 1 0 28520 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_334
timestamp 1624635492
transform 1 0 31832 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_322
timestamp 1624635492
transform 1 0 30728 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_355
timestamp 1624635492
transform 1 0 33764 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_343
timestamp 1624635492
transform 1 0 32660 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1624635492
transform 1 0 32568 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1624635492
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_391
timestamp 1624635492
transform 1 0 37076 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1624635492
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_400
timestamp 1624635492
transform 1 0 37904 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1624635492
transform 1 0 37812 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_282
timestamp 1624635492
transform 1 0 27048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_306
timestamp 1624635492
transform 1 0 29256 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_294
timestamp 1624635492
transform 1 0 28152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1624635492
transform 1 0 29992 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_327
timestamp 1624635492
transform 1 0 31188 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_315
timestamp 1624635492
transform 1 0 30084 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_351
timestamp 1624635492
transform 1 0 33396 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_339
timestamp 1624635492
transform 1 0 32292 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_372
timestamp 1624635492
transform 1 0 35328 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_363
timestamp 1624635492
transform 1 0 34500 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1624635492
transform 1 0 35236 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_396
timestamp 1624635492
transform 1 0 37536 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_384
timestamp 1624635492
transform 1 0 36432 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_408
timestamp 1624635492
transform 1 0 38640 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_286
timestamp 1624635492
transform 1 0 27416 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_277
timestamp 1624635492
transform 1 0 26588 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1624635492
transform 1 0 27324 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_310
timestamp 1624635492
transform 1 0 29624 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_298
timestamp 1624635492
transform 1 0 28520 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_334
timestamp 1624635492
transform 1 0 31832 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_322
timestamp 1624635492
transform 1 0 30728 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_355
timestamp 1624635492
transform 1 0 33764 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_343
timestamp 1624635492
transform 1 0 32660 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1624635492
transform 1 0 32568 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_377
timestamp 1624635492
transform 1 0 35788 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_373
timestamp 1624635492
transform 1 0 35420 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_367
timestamp 1624635492
transform 1 0 34868 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _278_
timestamp 1624635492
transform 1 0 35512 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_397
timestamp 1624635492
transform 1 0 37628 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_389
timestamp 1624635492
transform 1 0 36892 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_400
timestamp 1624635492
transform 1 0 37904 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1624635492
transform 1 0 37812 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_286
timestamp 1624635492
transform 1 0 27416 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_277
timestamp 1624635492
transform 1 0 26588 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_282
timestamp 1624635492
transform 1 0 27048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1624635492
transform 1 0 27324 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_310
timestamp 1624635492
transform 1 0 29624 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_298
timestamp 1624635492
transform 1 0 28520 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_306
timestamp 1624635492
transform 1 0 29256 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_294
timestamp 1624635492
transform 1 0 28152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1624635492
transform 1 0 29992 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_334
timestamp 1624635492
transform 1 0 31832 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_322
timestamp 1624635492
transform 1 0 30728 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_327
timestamp 1624635492
transform 1 0 31188 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_315
timestamp 1624635492
transform 1 0 30084 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_353
timestamp 1624635492
transform 1 0 33580 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_343
timestamp 1624635492
transform 1 0 32660 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_355
timestamp 1624635492
transform 1 0 33764 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_351
timestamp 1624635492
transform 1 0 33396 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_339
timestamp 1624635492
transform 1 0 32292 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__B
timestamp 1624635492
transform 1 0 33580 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__D
timestamp 1624635492
transform -1 0 33580 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1624635492
transform 1 0 32568 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_372
timestamp 1624635492
transform 1 0 35328 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_366
timestamp 1624635492
transform 1 0 34776 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_372
timestamp 1624635492
transform 1 0 35328 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_367
timestamp 1624635492
transform 1 0 34868 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__C
timestamp 1624635492
transform 1 0 35144 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1624635492
transform 1 0 35236 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _097_
timestamp 1624635492
transform 1 0 33948 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_67_396
timestamp 1624635492
transform 1 0 37536 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_384
timestamp 1624635492
transform 1 0 36432 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_396
timestamp 1624635492
transform 1 0 37536 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_384
timestamp 1624635492
transform 1 0 36432 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_400
timestamp 1624635492
transform 1 0 37904 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_408
timestamp 1624635492
transform 1 0 38640 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1624635492
transform 1 0 37812 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_282
timestamp 1624635492
transform 1 0 27048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_310
timestamp 1624635492
transform 1 0 29624 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_306
timestamp 1624635492
transform 1 0 29256 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_294
timestamp 1624635492
transform 1 0 28152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1624635492
transform 1 0 29992 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _321_
timestamp 1624635492
transform -1 0 29624 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_327
timestamp 1624635492
transform 1 0 31188 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_315
timestamp 1624635492
transform 1 0 30084 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_353
timestamp 1624635492
transform 1 0 33580 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_339
timestamp 1624635492
transform 1 0 32292 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1624635492
transform 1 0 33396 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_372
timestamp 1624635492
transform 1 0 35328 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_365
timestamp 1624635492
transform 1 0 34684 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1624635492
transform 1 0 35236 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_396
timestamp 1624635492
transform 1 0 37536 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_384
timestamp 1624635492
transform 1 0 36432 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_408
timestamp 1624635492
transform 1 0 38640 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_286
timestamp 1624635492
transform 1 0 27416 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_277
timestamp 1624635492
transform 1 0 26588 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1624635492
transform 1 0 27324 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_310
timestamp 1624635492
transform 1 0 29624 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_298
timestamp 1624635492
transform 1 0 28520 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_334
timestamp 1624635492
transform 1 0 31832 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_322
timestamp 1624635492
transform 1 0 30728 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_355
timestamp 1624635492
transform 1 0 33764 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_343
timestamp 1624635492
transform 1 0 32660 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1624635492
transform 1 0 32568 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_367
timestamp 1624635492
transform 1 0 34868 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_391
timestamp 1624635492
transform 1 0 37076 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1624635492
transform 1 0 35972 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_400
timestamp 1624635492
transform 1 0 37904 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1624635492
transform 1 0 37812 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_282
timestamp 1624635492
transform 1 0 27048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_306
timestamp 1624635492
transform 1 0 29256 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_294
timestamp 1624635492
transform 1 0 28152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1624635492
transform 1 0 29992 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_327
timestamp 1624635492
transform 1 0 31188 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_315
timestamp 1624635492
transform 1 0 30084 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_351
timestamp 1624635492
transform 1 0 33396 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_339
timestamp 1624635492
transform 1 0 32292 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_372
timestamp 1624635492
transform 1 0 35328 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_363
timestamp 1624635492
transform 1 0 34500 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1624635492
transform 1 0 35236 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_396
timestamp 1624635492
transform 1 0 37536 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_384
timestamp 1624635492
transform 1 0 36432 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_408
timestamp 1624635492
transform 1 0 38640 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_286
timestamp 1624635492
transform 1 0 27416 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_277
timestamp 1624635492
transform 1 0 26588 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1624635492
transform 1 0 27324 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_310
timestamp 1624635492
transform 1 0 29624 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_298
timestamp 1624635492
transform 1 0 28520 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_334
timestamp 1624635492
transform 1 0 31832 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_322
timestamp 1624635492
transform 1 0 30728 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_355
timestamp 1624635492
transform 1 0 33764 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_343
timestamp 1624635492
transform 1 0 32660 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1624635492
transform 1 0 32568 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1624635492
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_391
timestamp 1624635492
transform 1 0 37076 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1624635492
transform 1 0 35972 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_400
timestamp 1624635492
transform 1 0 37904 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1624635492
transform 1 0 37812 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_286
timestamp 1624635492
transform 1 0 27416 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_284
timestamp 1624635492
transform 1 0 27232 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_278
timestamp 1624635492
transform 1 0 26680 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_282
timestamp 1624635492
transform 1 0 27048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1624635492
transform 1 0 27324 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _285_
timestamp 1624635492
transform 1 0 26404 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_310
timestamp 1624635492
transform 1 0 29624 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_298
timestamp 1624635492
transform 1 0 28520 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_306
timestamp 1624635492
transform 1 0 29256 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_294
timestamp 1624635492
transform 1 0 28152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1624635492
transform 1 0 29992 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_334
timestamp 1624635492
transform 1 0 31832 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_322
timestamp 1624635492
transform 1 0 30728 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_324
timestamp 1624635492
transform 1 0 30912 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_321
timestamp 1624635492
transform 1 0 30636 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_315
timestamp 1624635492
transform 1 0 30084 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__CLK
timestamp 1624635492
transform 1 0 30728 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _343_
timestamp 1624635492
transform -1 0 33028 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_73_355
timestamp 1624635492
transform 1 0 33764 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_343
timestamp 1624635492
transform 1 0 32660 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_353
timestamp 1624635492
transform 1 0 33580 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_347
timestamp 1624635492
transform 1 0 33028 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__D
timestamp 1624635492
transform 1 0 33396 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1624635492
transform 1 0 32568 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1624635492
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_372
timestamp 1624635492
transform 1 0 35328 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_365
timestamp 1624635492
transform 1 0 34684 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1624635492
transform 1 0 35236 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _292_
timestamp 1624635492
transform 1 0 35696 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_391
timestamp 1624635492
transform 1 0 37076 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_379
timestamp 1624635492
transform 1 0 35972 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_391
timestamp 1624635492
transform 1 0 37076 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_379
timestamp 1624635492
transform 1 0 35972 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_400
timestamp 1624635492
transform 1 0 37904 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_403
timestamp 1624635492
transform 1 0 38180 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1624635492
transform 1 0 37812 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_282
timestamp 1624635492
transform 1 0 27048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_306
timestamp 1624635492
transform 1 0 29256 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_294
timestamp 1624635492
transform 1 0 28152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1624635492
transform 1 0 29992 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_327
timestamp 1624635492
transform 1 0 31188 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_315
timestamp 1624635492
transform 1 0 30084 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_351
timestamp 1624635492
transform 1 0 33396 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_339
timestamp 1624635492
transform 1 0 32292 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_372
timestamp 1624635492
transform 1 0 35328 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_363
timestamp 1624635492
transform 1 0 34500 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1624635492
transform 1 0 35236 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_396
timestamp 1624635492
transform 1 0 37536 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_384
timestamp 1624635492
transform 1 0 36432 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_408
timestamp 1624635492
transform 1 0 38640 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_286
timestamp 1624635492
transform 1 0 27416 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_277
timestamp 1624635492
transform 1 0 26588 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1624635492
transform 1 0 27324 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_310
timestamp 1624635492
transform 1 0 29624 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_298
timestamp 1624635492
transform 1 0 28520 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_334
timestamp 1624635492
transform 1 0 31832 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_322
timestamp 1624635492
transform 1 0 30728 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_355
timestamp 1624635492
transform 1 0 33764 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_343
timestamp 1624635492
transform 1 0 32660 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1624635492
transform 1 0 32568 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1624635492
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_391
timestamp 1624635492
transform 1 0 37076 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_379
timestamp 1624635492
transform 1 0 35972 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_400
timestamp 1624635492
transform 1 0 37904 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1624635492
transform 1 0 37812 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_282
timestamp 1624635492
transform 1 0 27048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_306
timestamp 1624635492
transform 1 0 29256 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_294
timestamp 1624635492
transform 1 0 28152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1624635492
transform 1 0 29992 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_328
timestamp 1624635492
transform 1 0 31280 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_322
timestamp 1624635492
transform 1 0 30728 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_315
timestamp 1624635492
transform 1 0 30084 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_wb_clk_i_A
timestamp 1624635492
transform 1 0 31096 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1624635492
transform -1 0 30728 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_352
timestamp 1624635492
transform 1 0 33488 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_340
timestamp 1624635492
transform 1 0 32384 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_372
timestamp 1624635492
transform 1 0 35328 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_370
timestamp 1624635492
transform 1 0 35144 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_364
timestamp 1624635492
transform 1 0 34592 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1624635492
transform 1 0 35236 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _169_
timestamp 1624635492
transform -1 0 35972 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_391
timestamp 1624635492
transform 1 0 37076 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_379
timestamp 1624635492
transform 1 0 35972 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_403
timestamp 1624635492
transform 1 0 38180 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_286
timestamp 1624635492
transform 1 0 27416 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_277
timestamp 1624635492
transform 1 0 26588 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1624635492
transform 1 0 27324 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_310
timestamp 1624635492
transform 1 0 29624 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_298
timestamp 1624635492
transform 1 0 28520 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_334
timestamp 1624635492
transform 1 0 31832 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_322
timestamp 1624635492
transform 1 0 30728 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_355
timestamp 1624635492
transform 1 0 33764 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_343
timestamp 1624635492
transform 1 0 32660 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1624635492
transform 1 0 32568 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_367
timestamp 1624635492
transform 1 0 34868 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_391
timestamp 1624635492
transform 1 0 37076 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_379
timestamp 1624635492
transform 1 0 35972 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_400
timestamp 1624635492
transform 1 0 37904 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1624635492
transform 1 0 37812 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_282
timestamp 1624635492
transform 1 0 27048 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_306
timestamp 1624635492
transform 1 0 29256 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_294
timestamp 1624635492
transform 1 0 28152 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1624635492
transform 1 0 29992 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_327
timestamp 1624635492
transform 1 0 31188 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_315
timestamp 1624635492
transform 1 0 30084 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_351
timestamp 1624635492
transform 1 0 33396 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_339
timestamp 1624635492
transform 1 0 32292 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_372
timestamp 1624635492
transform 1 0 35328 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_363
timestamp 1624635492
transform 1 0 34500 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1624635492
transform 1 0 35236 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_396
timestamp 1624635492
transform 1 0 37536 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_384
timestamp 1624635492
transform 1 0 36432 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_408
timestamp 1624635492
transform 1 0 38640 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_286
timestamp 1624635492
transform 1 0 27416 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_277
timestamp 1624635492
transform 1 0 26588 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1624635492
transform 1 0 27324 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_310
timestamp 1624635492
transform 1 0 29624 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_298
timestamp 1624635492
transform 1 0 28520 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_334
timestamp 1624635492
transform 1 0 31832 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_322
timestamp 1624635492
transform 1 0 30728 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_355
timestamp 1624635492
transform 1 0 33764 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_343
timestamp 1624635492
transform 1 0 32660 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1624635492
transform 1 0 32568 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_367
timestamp 1624635492
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_391
timestamp 1624635492
transform 1 0 37076 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_379
timestamp 1624635492
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_400
timestamp 1624635492
transform 1 0 37904 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1624635492
transform 1 0 37812 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_429
timestamp 1624635492
transform 1 0 40572 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_425
timestamp 1624635492
transform 1 0 40204 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_413
timestamp 1624635492
transform 1 0 39100 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_424
timestamp 1624635492
transform 1 0 40112 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_412
timestamp 1624635492
transform 1 0 39008 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__C1
timestamp 1624635492
transform -1 0 39100 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1624635492
transform 1 0 40480 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_441
timestamp 1624635492
transform 1 0 41676 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_448
timestamp 1624635492
transform 1 0 42320 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_436
timestamp 1624635492
transform 1 0 41216 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _273_
timestamp 1624635492
transform 1 0 42228 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_462
timestamp 1624635492
transform 1 0 43608 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_450
timestamp 1624635492
transform 1 0 42504 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_469
timestamp 1624635492
transform 1 0 44252 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_457
timestamp 1624635492
transform 1 0 43148 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1624635492
transform 1 0 43056 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_486
timestamp 1624635492
transform 1 0 45816 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_482
timestamp 1624635492
transform 1 0 45448 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_474
timestamp 1624635492
transform 1 0 44712 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_481
timestamp 1624635492
transform 1 0 45356 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1624635492
transform 1 0 45724 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_498
timestamp 1624635492
transform 1 0 46920 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1624635492
transform 1 0 47564 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_493
timestamp 1624635492
transform 1 0 46460 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_522
timestamp 1624635492
transform 1 0 49128 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_510
timestamp 1624635492
transform 1 0 48024 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_526
timestamp 1624635492
transform 1 0 49496 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_514
timestamp 1624635492
transform 1 0 48392 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1624635492
transform 1 0 48300 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_543
timestamp 1624635492
transform 1 0 51060 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_534
timestamp 1624635492
transform 1 0 50232 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_538
timestamp 1624635492
transform 1 0 50600 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1624635492
transform 1 0 50968 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_424
timestamp 1624635492
transform 1 0 40112 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_412
timestamp 1624635492
transform 1 0 39008 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_448
timestamp 1624635492
transform 1 0 42320 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_436
timestamp 1624635492
transform 1 0 41216 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_469
timestamp 1624635492
transform 1 0 44252 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_457
timestamp 1624635492
transform 1 0 43148 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1624635492
transform 1 0 43056 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_481
timestamp 1624635492
transform 1 0 45356 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1624635492
transform 1 0 47564 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_493
timestamp 1624635492
transform 1 0 46460 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_526
timestamp 1624635492
transform 1 0 49496 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_514
timestamp 1624635492
transform 1 0 48392 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1624635492
transform 1 0 48300 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_538
timestamp 1624635492
transform 1 0 50600 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_429
timestamp 1624635492
transform 1 0 40572 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_420
timestamp 1624635492
transform 1 0 39744 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1624635492
transform 1 0 40480 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_441
timestamp 1624635492
transform 1 0 41676 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_465
timestamp 1624635492
transform 1 0 43884 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_453
timestamp 1624635492
transform 1 0 42780 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_486
timestamp 1624635492
transform 1 0 45816 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_477
timestamp 1624635492
transform 1 0 44988 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1624635492
transform 1 0 45724 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_498
timestamp 1624635492
transform 1 0 46920 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_522
timestamp 1624635492
transform 1 0 49128 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_510
timestamp 1624635492
transform 1 0 48024 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_543
timestamp 1624635492
transform 1 0 51060 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_534
timestamp 1624635492
transform 1 0 50232 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1624635492
transform 1 0 50968 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_428
timestamp 1624635492
transform 1 0 40480 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_416
timestamp 1624635492
transform 1 0 39376 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_412
timestamp 1624635492
transform 1 0 39008 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _280_
timestamp 1624635492
transform 1 0 39100 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_440
timestamp 1624635492
transform 1 0 41584 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_469
timestamp 1624635492
transform 1 0 44252 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_457
timestamp 1624635492
transform 1 0 43148 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_452
timestamp 1624635492
transform 1 0 42688 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1624635492
transform 1 0 43056 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_481
timestamp 1624635492
transform 1 0 45356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1624635492
transform 1 0 47564 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_493
timestamp 1624635492
transform 1 0 46460 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_526
timestamp 1624635492
transform 1 0 49496 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_514
timestamp 1624635492
transform 1 0 48392 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1624635492
transform 1 0 48300 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_538
timestamp 1624635492
transform 1 0 50600 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_429
timestamp 1624635492
transform 1 0 40572 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_420
timestamp 1624635492
transform 1 0 39744 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1624635492
transform 1 0 40480 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_441
timestamp 1624635492
transform 1 0 41676 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_465
timestamp 1624635492
transform 1 0 43884 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_453
timestamp 1624635492
transform 1 0 42780 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_486
timestamp 1624635492
transform 1 0 45816 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_477
timestamp 1624635492
transform 1 0 44988 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1624635492
transform 1 0 45724 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_498
timestamp 1624635492
transform 1 0 46920 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_522
timestamp 1624635492
transform 1 0 49128 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_510
timestamp 1624635492
transform 1 0 48024 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_543
timestamp 1624635492
transform 1 0 51060 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_534
timestamp 1624635492
transform 1 0 50232 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1624635492
transform 1 0 50968 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_429
timestamp 1624635492
transform 1 0 40572 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_420
timestamp 1624635492
transform 1 0 39744 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_424
timestamp 1624635492
transform 1 0 40112 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_412
timestamp 1624635492
transform 1 0 39008 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1624635492
transform 1 0 40480 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_441
timestamp 1624635492
transform 1 0 41676 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_448
timestamp 1624635492
transform 1 0 42320 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_436
timestamp 1624635492
transform 1 0 41216 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_465
timestamp 1624635492
transform 1 0 43884 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_453
timestamp 1624635492
transform 1 0 42780 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_469
timestamp 1624635492
transform 1 0 44252 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_457
timestamp 1624635492
transform 1 0 43148 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1624635492
transform 1 0 43056 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_486
timestamp 1624635492
transform 1 0 45816 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_477
timestamp 1624635492
transform 1 0 44988 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_481
timestamp 1624635492
transform 1 0 45356 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_474
timestamp 1624635492
transform 1 0 44712 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1624635492
transform 1 0 45724 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _309_
timestamp 1624635492
transform -1 0 45356 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _134_
timestamp 1624635492
transform -1 0 44712 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_498
timestamp 1624635492
transform 1 0 46920 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1624635492
transform 1 0 47564 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_493
timestamp 1624635492
transform 1 0 46460 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_522
timestamp 1624635492
transform 1 0 49128 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_510
timestamp 1624635492
transform 1 0 48024 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_526
timestamp 1624635492
transform 1 0 49496 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_514
timestamp 1624635492
transform 1 0 48392 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1624635492
transform 1 0 48300 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_543
timestamp 1624635492
transform 1 0 51060 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_534
timestamp 1624635492
transform 1 0 50232 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_538
timestamp 1624635492
transform 1 0 50600 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1624635492
transform 1 0 50968 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_424
timestamp 1624635492
transform 1 0 40112 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_412
timestamp 1624635492
transform 1 0 39008 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_440
timestamp 1624635492
transform 1 0 41584 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_436
timestamp 1624635492
transform 1 0 41216 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__CLK
timestamp 1624635492
transform 1 0 41400 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_457
timestamp 1624635492
transform 1 0 43148 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_452
timestamp 1624635492
transform 1 0 42688 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1624635492
transform 1 0 43056 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _248_
timestamp 1624635492
transform 1 0 44252 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_484
timestamp 1624635492
transform 1 0 45632 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_472
timestamp 1624635492
transform 1 0 44528 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_508
timestamp 1624635492
transform 1 0 47840 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_496
timestamp 1624635492
transform 1 0 46736 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_526
timestamp 1624635492
transform 1 0 49496 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_514
timestamp 1624635492
transform 1 0 48392 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_512
timestamp 1624635492
transform 1 0 48208 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1624635492
transform 1 0 48300 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_538
timestamp 1624635492
transform 1 0 50600 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_429
timestamp 1624635492
transform 1 0 40572 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_420
timestamp 1624635492
transform 1 0 39744 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1624635492
transform 1 0 40480 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_438
timestamp 1624635492
transform 1 0 41400 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_435
timestamp 1624635492
transform 1 0 41124 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__D
timestamp 1624635492
transform -1 0 41400 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _340_
timestamp 1624635492
transform 1 0 41768 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_461
timestamp 1624635492
transform 1 0 43516 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_486
timestamp 1624635492
transform 1 0 45816 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_473
timestamp 1624635492
transform 1 0 44620 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1624635492
transform 1 0 45724 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_498
timestamp 1624635492
transform 1 0 46920 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_522
timestamp 1624635492
transform 1 0 49128 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_510
timestamp 1624635492
transform 1 0 48024 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_543
timestamp 1624635492
transform 1 0 51060 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_534
timestamp 1624635492
transform 1 0 50232 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1624635492
transform 1 0 50968 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_424
timestamp 1624635492
transform 1 0 40112 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_412
timestamp 1624635492
transform 1 0 39008 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_448
timestamp 1624635492
transform 1 0 42320 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_436
timestamp 1624635492
transform 1 0 41216 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_469
timestamp 1624635492
transform 1 0 44252 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_457
timestamp 1624635492
transform 1 0 43148 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1624635492
transform 1 0 43056 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_481
timestamp 1624635492
transform 1 0 45356 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1624635492
transform 1 0 47564 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_493
timestamp 1624635492
transform 1 0 46460 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_526
timestamp 1624635492
transform 1 0 49496 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_514
timestamp 1624635492
transform 1 0 48392 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1624635492
transform 1 0 48300 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_538
timestamp 1624635492
transform 1 0 50600 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_429
timestamp 1624635492
transform 1 0 40572 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_420
timestamp 1624635492
transform 1 0 39744 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1624635492
transform 1 0 40480 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_441
timestamp 1624635492
transform 1 0 41676 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_465
timestamp 1624635492
transform 1 0 43884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_453
timestamp 1624635492
transform 1 0 42780 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_486
timestamp 1624635492
transform 1 0 45816 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_477
timestamp 1624635492
transform 1 0 44988 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1624635492
transform 1 0 45724 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_498
timestamp 1624635492
transform 1 0 46920 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_522
timestamp 1624635492
transform 1 0 49128 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_510
timestamp 1624635492
transform 1 0 48024 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_543
timestamp 1624635492
transform 1 0 51060 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_534
timestamp 1624635492
transform 1 0 50232 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1624635492
transform 1 0 50968 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_424
timestamp 1624635492
transform 1 0 40112 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_412
timestamp 1624635492
transform 1 0 39008 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_445
timestamp 1624635492
transform 1 0 42044 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_433
timestamp 1624635492
transform 1 0 40940 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _194_
timestamp 1624635492
transform -1 0 40940 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_469
timestamp 1624635492
transform 1 0 44252 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_457
timestamp 1624635492
transform 1 0 43148 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_453
timestamp 1624635492
transform 1 0 42780 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1624635492
transform 1 0 43056 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_481
timestamp 1624635492
transform 1 0 45356 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _138_
timestamp 1624635492
transform -1 0 46368 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_504
timestamp 1624635492
transform 1 0 47472 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_492
timestamp 1624635492
transform 1 0 46368 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_526
timestamp 1624635492
transform 1 0 49496 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_514
timestamp 1624635492
transform 1 0 48392 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_512
timestamp 1624635492
transform 1 0 48208 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1624635492
transform 1 0 48300 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_538
timestamp 1624635492
transform 1 0 50600 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_424
timestamp 1624635492
transform 1 0 40112 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_412
timestamp 1624635492
transform 1 0 39008 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_429
timestamp 1624635492
transform 1 0 40572 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_420
timestamp 1624635492
transform 1 0 39744 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1624635492
transform 1 0 40480 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_448
timestamp 1624635492
transform 1 0 42320 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_436
timestamp 1624635492
transform 1 0 41216 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_448
timestamp 1624635492
transform 1 0 42320 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_436
timestamp 1624635492
transform 1 0 41216 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _298_
timestamp 1624635492
transform -1 0 41216 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_469
timestamp 1624635492
transform 1 0 44252 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_457
timestamp 1624635492
transform 1 0 43148 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_460
timestamp 1624635492
transform 1 0 43424 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1624635492
transform 1 0 43056 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_481
timestamp 1624635492
transform 1 0 45356 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_486
timestamp 1624635492
transform 1 0 45816 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_484
timestamp 1624635492
transform 1 0 45632 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_472
timestamp 1624635492
transform 1 0 44528 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1624635492
transform 1 0 45724 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1624635492
transform 1 0 47564 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_493
timestamp 1624635492
transform 1 0 46460 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_498
timestamp 1624635492
transform 1 0 46920 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_521
timestamp 1624635492
transform 1 0 49036 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_514
timestamp 1624635492
transform 1 0 48392 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_522
timestamp 1624635492
transform 1 0 49128 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_510
timestamp 1624635492
transform 1 0 48024 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1624635492
transform 1 0 48300 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _291_
timestamp 1624635492
transform 1 0 48760 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_545
timestamp 1624635492
transform 1 0 51244 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_533
timestamp 1624635492
transform 1 0 50140 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_543
timestamp 1624635492
transform 1 0 51060 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_534
timestamp 1624635492
transform 1 0 50232 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1624635492
transform 1 0 50968 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_429
timestamp 1624635492
transform 1 0 40572 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_420
timestamp 1624635492
transform 1 0 39744 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1624635492
transform 1 0 40480 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_441
timestamp 1624635492
transform 1 0 41676 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_465
timestamp 1624635492
transform 1 0 43884 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_453
timestamp 1624635492
transform 1 0 42780 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_486
timestamp 1624635492
transform 1 0 45816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_477
timestamp 1624635492
transform 1 0 44988 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1624635492
transform 1 0 45724 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_498
timestamp 1624635492
transform 1 0 46920 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_522
timestamp 1624635492
transform 1 0 49128 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_510
timestamp 1624635492
transform 1 0 48024 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_543
timestamp 1624635492
transform 1 0 51060 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_534
timestamp 1624635492
transform 1 0 50232 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1624635492
transform 1 0 50968 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_424
timestamp 1624635492
transform 1 0 40112 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_412
timestamp 1624635492
transform 1 0 39008 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_448
timestamp 1624635492
transform 1 0 42320 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_436
timestamp 1624635492
transform 1 0 41216 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_469
timestamp 1624635492
transform 1 0 44252 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_457
timestamp 1624635492
transform 1 0 43148 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1624635492
transform 1 0 43056 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_481
timestamp 1624635492
transform 1 0 45356 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1624635492
transform 1 0 47564 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_493
timestamp 1624635492
transform 1 0 46460 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_526
timestamp 1624635492
transform 1 0 49496 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_514
timestamp 1624635492
transform 1 0 48392 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1624635492
transform 1 0 48300 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_538
timestamp 1624635492
transform 1 0 50600 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_429
timestamp 1624635492
transform 1 0 40572 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_420
timestamp 1624635492
transform 1 0 39744 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1624635492
transform 1 0 40480 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_441
timestamp 1624635492
transform 1 0 41676 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_465
timestamp 1624635492
transform 1 0 43884 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_453
timestamp 1624635492
transform 1 0 42780 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_486
timestamp 1624635492
transform 1 0 45816 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_477
timestamp 1624635492
transform 1 0 44988 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1624635492
transform 1 0 45724 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_498
timestamp 1624635492
transform 1 0 46920 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_522
timestamp 1624635492
transform 1 0 49128 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_510
timestamp 1624635492
transform 1 0 48024 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_543
timestamp 1624635492
transform 1 0 51060 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_534
timestamp 1624635492
transform 1 0 50232 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1624635492
transform 1 0 50968 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_424
timestamp 1624635492
transform 1 0 40112 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_412
timestamp 1624635492
transform 1 0 39008 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_448
timestamp 1624635492
transform 1 0 42320 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_436
timestamp 1624635492
transform 1 0 41216 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_464
timestamp 1624635492
transform 1 0 43792 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_457
timestamp 1624635492
transform 1 0 43148 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1624635492
transform 1 0 43056 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _181_
timestamp 1624635492
transform -1 0 43792 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_488
timestamp 1624635492
transform 1 0 46000 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_476
timestamp 1624635492
transform 1 0 44896 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_502
timestamp 1624635492
transform 1 0 47288 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_496
timestamp 1624635492
transform 1 0 46736 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _210_
timestamp 1624635492
transform -1 0 47288 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_526
timestamp 1624635492
transform 1 0 49496 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_514
timestamp 1624635492
transform 1 0 48392 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_510
timestamp 1624635492
transform 1 0 48024 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1624635492
transform 1 0 48300 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_538
timestamp 1624635492
transform 1 0 50600 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_424
timestamp 1624635492
transform 1 0 40112 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_412
timestamp 1624635492
transform 1 0 39008 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_429
timestamp 1624635492
transform 1 0 40572 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_427
timestamp 1624635492
transform 1 0 40388 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_415
timestamp 1624635492
transform 1 0 39284 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1624635492
transform 1 0 40480 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_448
timestamp 1624635492
transform 1 0 42320 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_436
timestamp 1624635492
transform 1 0 41216 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_441
timestamp 1624635492
transform 1 0 41676 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_469
timestamp 1624635492
transform 1 0 44252 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_457
timestamp 1624635492
transform 1 0 43148 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_465
timestamp 1624635492
transform 1 0 43884 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_453
timestamp 1624635492
transform 1 0 42780 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1624635492
transform 1 0 43056 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_481
timestamp 1624635492
transform 1 0 45356 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_486
timestamp 1624635492
transform 1 0 45816 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_477
timestamp 1624635492
transform 1 0 44988 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1624635492
transform 1 0 45724 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1624635492
transform 1 0 47564 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_493
timestamp 1624635492
transform 1 0 46460 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_498
timestamp 1624635492
transform 1 0 46920 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_526
timestamp 1624635492
transform 1 0 49496 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_514
timestamp 1624635492
transform 1 0 48392 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_522
timestamp 1624635492
transform 1 0 49128 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_510
timestamp 1624635492
transform 1 0 48024 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1624635492
transform 1 0 48300 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_538
timestamp 1624635492
transform 1 0 50600 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_543
timestamp 1624635492
transform 1 0 51060 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_534
timestamp 1624635492
transform 1 0 50232 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1624635492
transform 1 0 50968 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _227_
timestamp 1624635492
transform -1 0 51612 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_429
timestamp 1624635492
transform 1 0 40572 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_420
timestamp 1624635492
transform 1 0 39744 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1624635492
transform 1 0 40480 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_441
timestamp 1624635492
transform 1 0 41676 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_465
timestamp 1624635492
transform 1 0 43884 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_453
timestamp 1624635492
transform 1 0 42780 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_486
timestamp 1624635492
transform 1 0 45816 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_477
timestamp 1624635492
transform 1 0 44988 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1624635492
transform 1 0 45724 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_498
timestamp 1624635492
transform 1 0 46920 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_521
timestamp 1624635492
transform 1 0 49036 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_518
timestamp 1624635492
transform 1 0 48760 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_510
timestamp 1624635492
transform 1 0 48024 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1624635492
transform 1 0 48852 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 49404 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_543
timestamp 1624635492
transform 1 0 51060 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_541
timestamp 1624635492
transform 1 0 50876 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_537
timestamp 1624635492
transform 1 0 50508 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1624635492
transform 1 0 50968 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_424
timestamp 1624635492
transform 1 0 40112 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_412
timestamp 1624635492
transform 1 0 39008 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_448
timestamp 1624635492
transform 1 0 42320 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_436
timestamp 1624635492
transform 1 0 41216 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_469
timestamp 1624635492
transform 1 0 44252 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_457
timestamp 1624635492
transform 1 0 43148 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1624635492
transform 1 0 43056 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_481
timestamp 1624635492
transform 1 0 45356 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1624635492
transform 1 0 47564 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_493
timestamp 1624635492
transform 1 0 46460 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_526
timestamp 1624635492
transform 1 0 49496 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_514
timestamp 1624635492
transform 1 0 48392 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1624635492
transform 1 0 48300 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_545
timestamp 1624635492
transform 1 0 51244 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_533
timestamp 1624635492
transform 1 0 50140 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _293_
timestamp 1624635492
transform 1 0 49864 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_429
timestamp 1624635492
transform 1 0 40572 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_427
timestamp 1624635492
transform 1 0 40388 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_415
timestamp 1624635492
transform 1 0 39284 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1624635492
transform 1 0 40480 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_441
timestamp 1624635492
transform 1 0 41676 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_465
timestamp 1624635492
transform 1 0 43884 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_453
timestamp 1624635492
transform 1 0 42780 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_486
timestamp 1624635492
transform 1 0 45816 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_477
timestamp 1624635492
transform 1 0 44988 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1624635492
transform 1 0 45724 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_498
timestamp 1624635492
transform 1 0 46920 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_522
timestamp 1624635492
transform 1 0 49128 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_510
timestamp 1624635492
transform 1 0 48024 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_543
timestamp 1624635492
transform 1 0 51060 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_534
timestamp 1624635492
transform 1 0 50232 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1624635492
transform 1 0 50968 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_424
timestamp 1624635492
transform 1 0 40112 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_412
timestamp 1624635492
transform 1 0 39008 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_448
timestamp 1624635492
transform 1 0 42320 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_436
timestamp 1624635492
transform 1 0 41216 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_469
timestamp 1624635492
transform 1 0 44252 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_457
timestamp 1624635492
transform 1 0 43148 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1624635492
transform 1 0 43056 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_481
timestamp 1624635492
transform 1 0 45356 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1624635492
transform 1 0 47564 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_493
timestamp 1624635492
transform 1 0 46460 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_526
timestamp 1624635492
transform 1 0 49496 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_514
timestamp 1624635492
transform 1 0 48392 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1624635492
transform 1 0 48300 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_538
timestamp 1624635492
transform 1 0 50600 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_429
timestamp 1624635492
transform 1 0 40572 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_427
timestamp 1624635492
transform 1 0 40388 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_419
timestamp 1624635492
transform 1 0 39652 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_416
timestamp 1624635492
transform 1 0 39376 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__B1
timestamp 1624635492
transform 1 0 39468 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1624635492
transform 1 0 40480 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_441
timestamp 1624635492
transform 1 0 41676 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_465
timestamp 1624635492
transform 1 0 43884 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_453
timestamp 1624635492
transform 1 0 42780 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_486
timestamp 1624635492
transform 1 0 45816 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_477
timestamp 1624635492
transform 1 0 44988 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1624635492
transform 1 0 45724 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_498
timestamp 1624635492
transform 1 0 46920 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_522
timestamp 1624635492
transform 1 0 49128 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_510
timestamp 1624635492
transform 1 0 48024 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_543
timestamp 1624635492
transform 1 0 51060 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_534
timestamp 1624635492
transform 1 0 50232 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1624635492
transform 1 0 50968 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_429
timestamp 1624635492
transform 1 0 40572 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_417
timestamp 1624635492
transform 1 0 39468 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_412
timestamp 1624635492
transform 1 0 39008 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A2
timestamp 1624635492
transform 1 0 39284 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _056_
timestamp 1624635492
transform -1 0 40572 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_447
timestamp 1624635492
transform 1 0 42228 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_435
timestamp 1624635492
transform 1 0 41124 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__B2
timestamp 1624635492
transform 1 0 40940 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_469
timestamp 1624635492
transform 1 0 44252 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_457
timestamp 1624635492
transform 1 0 43148 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_455
timestamp 1624635492
transform 1 0 42964 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1624635492
transform 1 0 43056 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_481
timestamp 1624635492
transform 1 0 45356 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1624635492
transform 1 0 47564 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_493
timestamp 1624635492
transform 1 0 46460 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_526
timestamp 1624635492
transform 1 0 49496 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_514
timestamp 1624635492
transform 1 0 48392 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1624635492
transform 1 0 48300 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_538
timestamp 1624635492
transform 1 0 50600 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_555
timestamp 1624635492
transform 1 0 52164 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_562
timestamp 1624635492
transform 1 0 52808 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_550
timestamp 1624635492
transform 1 0 51704 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_583
timestamp 1624635492
transform 1 0 54740 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_579
timestamp 1624635492
transform 1 0 54372 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_567
timestamp 1624635492
transform 1 0 53268 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_583
timestamp 1624635492
transform 1 0 54740 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_571
timestamp 1624635492
transform 1 0 53636 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__B
timestamp 1624635492
transform 1 0 54832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1624635492
transform 1 0 53544 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_602
timestamp 1624635492
transform 1 0 56488 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_595
timestamp 1624635492
transform 1 0 55844 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_586
timestamp 1624635492
transform 1 0 55016 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_595
timestamp 1624635492
transform 1 0 55844 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1624635492
transform 1 0 56304 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1624635492
transform 1 0 56212 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 55384 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_54_614
timestamp 1624635492
transform 1 0 57592 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_619
timestamp 1624635492
transform 1 0 58052 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_607
timestamp 1624635492
transform 1 0 56948 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_638
timestamp 1624635492
transform 1 0 59800 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_626
timestamp 1624635492
transform 1 0 58696 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_640
timestamp 1624635492
transform 1 0 59984 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_628
timestamp 1624635492
transform 1 0 58880 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1624635492
transform 1 0 58788 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1624635492
transform 1 0 61548 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_650
timestamp 1624635492
transform 1 0 60904 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_664
timestamp 1624635492
transform 1 0 62192 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_652
timestamp 1624635492
transform 1 0 61088 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1624635492
transform 1 0 61456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_681
timestamp 1624635492
transform 1 0 63756 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_669
timestamp 1624635492
transform 1 0 62652 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_676
timestamp 1624635492
transform 1 0 63296 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_562
timestamp 1624635492
transform 1 0 52808 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_550
timestamp 1624635492
transform 1 0 51704 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_583
timestamp 1624635492
transform 1 0 54740 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_571
timestamp 1624635492
transform 1 0 53636 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1624635492
transform 1 0 53544 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_595
timestamp 1624635492
transform 1 0 55844 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_619
timestamp 1624635492
transform 1 0 58052 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_607
timestamp 1624635492
transform 1 0 56948 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_640
timestamp 1624635492
transform 1 0 59984 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_628
timestamp 1624635492
transform 1 0 58880 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1624635492
transform 1 0 58788 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_664
timestamp 1624635492
transform 1 0 62192 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_652
timestamp 1624635492
transform 1 0 61088 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_676
timestamp 1624635492
transform 1 0 63296 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_555
timestamp 1624635492
transform 1 0 52164 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_579
timestamp 1624635492
transform 1 0 54372 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_567
timestamp 1624635492
transform 1 0 53268 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_600
timestamp 1624635492
transform 1 0 56304 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_591
timestamp 1624635492
transform 1 0 55476 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1624635492
transform 1 0 56212 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_624
timestamp 1624635492
transform 1 0 58512 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_612
timestamp 1624635492
transform 1 0 57408 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_636
timestamp 1624635492
transform 1 0 59616 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1624635492
transform 1 0 61548 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_648
timestamp 1624635492
transform 1 0 60720 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1624635492
transform 1 0 61456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1624635492
transform 1 0 63756 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1624635492
transform 1 0 62652 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_562
timestamp 1624635492
transform 1 0 52808 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_550
timestamp 1624635492
transform 1 0 51704 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_583
timestamp 1624635492
transform 1 0 54740 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_571
timestamp 1624635492
transform 1 0 53636 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1624635492
transform 1 0 53544 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_595
timestamp 1624635492
transform 1 0 55844 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_619
timestamp 1624635492
transform 1 0 58052 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_607
timestamp 1624635492
transform 1 0 56948 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_640
timestamp 1624635492
transform 1 0 59984 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_628
timestamp 1624635492
transform 1 0 58880 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1624635492
transform 1 0 58788 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_664
timestamp 1624635492
transform 1 0 62192 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_652
timestamp 1624635492
transform 1 0 61088 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_675
timestamp 1624635492
transform 1 0 63204 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _183_
timestamp 1624635492
transform -1 0 63204 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_555
timestamp 1624635492
transform 1 0 52164 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_579
timestamp 1624635492
transform 1 0 54372 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_567
timestamp 1624635492
transform 1 0 53268 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_600
timestamp 1624635492
transform 1 0 56304 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_598
timestamp 1624635492
transform 1 0 56120 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_592
timestamp 1624635492
transform 1 0 55568 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_587
timestamp 1624635492
transform 1 0 55108 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1624635492
transform 1 0 56212 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _204_
timestamp 1624635492
transform -1 0 55568 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_624
timestamp 1624635492
transform 1 0 58512 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_612
timestamp 1624635492
transform 1 0 57408 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_636
timestamp 1624635492
transform 1 0 59616 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1624635492
transform 1 0 61548 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_648
timestamp 1624635492
transform 1 0 60720 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1624635492
transform 1 0 61456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1624635492
transform 1 0 63756 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1624635492
transform 1 0 62652 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_555
timestamp 1624635492
transform 1 0 52164 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_562
timestamp 1624635492
transform 1 0 52808 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_550
timestamp 1624635492
transform 1 0 51704 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_579
timestamp 1624635492
transform 1 0 54372 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_567
timestamp 1624635492
transform 1 0 53268 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_583
timestamp 1624635492
transform 1 0 54740 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_571
timestamp 1624635492
transform 1 0 53636 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1624635492
transform 1 0 53544 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_600
timestamp 1624635492
transform 1 0 56304 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_591
timestamp 1624635492
transform 1 0 55476 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_595
timestamp 1624635492
transform 1 0 55844 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1624635492
transform 1 0 56212 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_624
timestamp 1624635492
transform 1 0 58512 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_612
timestamp 1624635492
transform 1 0 57408 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_619
timestamp 1624635492
transform 1 0 58052 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_607
timestamp 1624635492
transform 1 0 56948 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_636
timestamp 1624635492
transform 1 0 59616 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_640
timestamp 1624635492
transform 1 0 59984 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_628
timestamp 1624635492
transform 1 0 58880 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1624635492
transform 1 0 58788 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_657
timestamp 1624635492
transform 1 0 61548 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_652
timestamp 1624635492
transform 1 0 61088 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_648
timestamp 1624635492
transform 1 0 60720 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_664
timestamp 1624635492
transform 1 0 62192 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_652
timestamp 1624635492
transform 1 0 61088 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1624635492
transform 1 0 61456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _310_
timestamp 1624635492
transform -1 0 61088 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1624635492
transform 1 0 63756 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_669
timestamp 1624635492
transform 1 0 62652 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_676
timestamp 1624635492
transform 1 0 63296 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_562
timestamp 1624635492
transform 1 0 52808 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_550
timestamp 1624635492
transform 1 0 51704 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_583
timestamp 1624635492
transform 1 0 54740 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_571
timestamp 1624635492
transform 1 0 53636 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1624635492
transform 1 0 53544 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_596
timestamp 1624635492
transform 1 0 55936 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_591
timestamp 1624635492
transform 1 0 55476 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _288_
timestamp 1624635492
transform 1 0 55660 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_620
timestamp 1624635492
transform 1 0 58144 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_608
timestamp 1624635492
transform 1 0 57040 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_640
timestamp 1624635492
transform 1 0 59984 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_628
timestamp 1624635492
transform 1 0 58880 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_626
timestamp 1624635492
transform 1 0 58696 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1624635492
transform 1 0 58788 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_650
timestamp 1624635492
transform 1 0 60904 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__CLK
timestamp 1624635492
transform 1 0 60720 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _344_
timestamp 1624635492
transform 1 0 61272 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_61_681
timestamp 1624635492
transform 1 0 63756 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_673
timestamp 1624635492
transform 1 0 63020 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_562
timestamp 1624635492
transform 1 0 52808 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_550
timestamp 1624635492
transform 1 0 51704 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _225_
timestamp 1624635492
transform -1 0 51704 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_574
timestamp 1624635492
transform 1 0 53912 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_600
timestamp 1624635492
transform 1 0 56304 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_598
timestamp 1624635492
transform 1 0 56120 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_586
timestamp 1624635492
transform 1 0 55016 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1624635492
transform 1 0 56212 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_624
timestamp 1624635492
transform 1 0 58512 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_612
timestamp 1624635492
transform 1 0 57408 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_636
timestamp 1624635492
transform 1 0 59616 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1624635492
transform 1 0 61548 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_648
timestamp 1624635492
transform 1 0 60720 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1624635492
transform 1 0 61456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_681
timestamp 1624635492
transform 1 0 63756 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_669
timestamp 1624635492
transform 1 0 62652 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_562
timestamp 1624635492
transform 1 0 52808 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_550
timestamp 1624635492
transform 1 0 51704 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_583
timestamp 1624635492
transform 1 0 54740 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_571
timestamp 1624635492
transform 1 0 53636 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1624635492
transform 1 0 53544 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_595
timestamp 1624635492
transform 1 0 55844 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_619
timestamp 1624635492
transform 1 0 58052 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_607
timestamp 1624635492
transform 1 0 56948 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_640
timestamp 1624635492
transform 1 0 59984 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_628
timestamp 1624635492
transform 1 0 58880 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1624635492
transform 1 0 58788 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_664
timestamp 1624635492
transform 1 0 62192 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_652
timestamp 1624635492
transform 1 0 61088 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_676
timestamp 1624635492
transform 1 0 63296 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_555
timestamp 1624635492
transform 1 0 52164 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_579
timestamp 1624635492
transform 1 0 54372 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_567
timestamp 1624635492
transform 1 0 53268 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_600
timestamp 1624635492
transform 1 0 56304 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_591
timestamp 1624635492
transform 1 0 55476 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1624635492
transform 1 0 56212 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_624
timestamp 1624635492
transform 1 0 58512 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_612
timestamp 1624635492
transform 1 0 57408 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_636
timestamp 1624635492
transform 1 0 59616 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_657
timestamp 1624635492
transform 1 0 61548 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_648
timestamp 1624635492
transform 1 0 60720 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1624635492
transform 1 0 61456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_681
timestamp 1624635492
transform 1 0 63756 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_669
timestamp 1624635492
transform 1 0 62652 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_562
timestamp 1624635492
transform 1 0 52808 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_550
timestamp 1624635492
transform 1 0 51704 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_583
timestamp 1624635492
transform 1 0 54740 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_571
timestamp 1624635492
transform 1 0 53636 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1624635492
transform 1 0 53544 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_595
timestamp 1624635492
transform 1 0 55844 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_619
timestamp 1624635492
transform 1 0 58052 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_607
timestamp 1624635492
transform 1 0 56948 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_640
timestamp 1624635492
transform 1 0 59984 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_628
timestamp 1624635492
transform 1 0 58880 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1624635492
transform 1 0 58788 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_664
timestamp 1624635492
transform 1 0 62192 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_652
timestamp 1624635492
transform 1 0 61088 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_676
timestamp 1624635492
transform 1 0 63296 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_557
timestamp 1624635492
transform 1 0 52348 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_555
timestamp 1624635492
transform 1 0 52164 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_583
timestamp 1624635492
transform 1 0 54740 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_571
timestamp 1624635492
transform 1 0 53636 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_569
timestamp 1624635492
transform 1 0 53452 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_579
timestamp 1624635492
transform 1 0 54372 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_567
timestamp 1624635492
transform 1 0 53268 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1624635492
transform 1 0 53544 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_595
timestamp 1624635492
transform 1 0 55844 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_600
timestamp 1624635492
transform 1 0 56304 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_591
timestamp 1624635492
transform 1 0 55476 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1624635492
transform 1 0 56212 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_619
timestamp 1624635492
transform 1 0 58052 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_607
timestamp 1624635492
transform 1 0 56948 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_624
timestamp 1624635492
transform 1 0 58512 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_612
timestamp 1624635492
transform 1 0 57408 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_640
timestamp 1624635492
transform 1 0 59984 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_628
timestamp 1624635492
transform 1 0 58880 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_636
timestamp 1624635492
transform 1 0 59616 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1624635492
transform 1 0 58788 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_664
timestamp 1624635492
transform 1 0 62192 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_652
timestamp 1624635492
transform 1 0 61088 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_657
timestamp 1624635492
transform 1 0 61548 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_648
timestamp 1624635492
transform 1 0 60720 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1624635492
transform 1 0 61456 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_676
timestamp 1624635492
transform 1 0 63296 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_681
timestamp 1624635492
transform 1 0 63756 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_669
timestamp 1624635492
transform 1 0 62652 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_555
timestamp 1624635492
transform 1 0 52164 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_579
timestamp 1624635492
transform 1 0 54372 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_567
timestamp 1624635492
transform 1 0 53268 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_600
timestamp 1624635492
transform 1 0 56304 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_591
timestamp 1624635492
transform 1 0 55476 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1624635492
transform 1 0 56212 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_624
timestamp 1624635492
transform 1 0 58512 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_612
timestamp 1624635492
transform 1 0 57408 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_636
timestamp 1624635492
transform 1 0 59616 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_657
timestamp 1624635492
transform 1 0 61548 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_648
timestamp 1624635492
transform 1 0 60720 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1624635492
transform 1 0 61456 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_681
timestamp 1624635492
transform 1 0 63756 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_669
timestamp 1624635492
transform 1 0 62652 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_562
timestamp 1624635492
transform 1 0 52808 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_550
timestamp 1624635492
transform 1 0 51704 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_583
timestamp 1624635492
transform 1 0 54740 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_571
timestamp 1624635492
transform 1 0 53636 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1624635492
transform 1 0 53544 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_595
timestamp 1624635492
transform 1 0 55844 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_619
timestamp 1624635492
transform 1 0 58052 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_607
timestamp 1624635492
transform 1 0 56948 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_640
timestamp 1624635492
transform 1 0 59984 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_628
timestamp 1624635492
transform 1 0 58880 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1624635492
transform 1 0 58788 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_664
timestamp 1624635492
transform 1 0 62192 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_652
timestamp 1624635492
transform 1 0 61088 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_676
timestamp 1624635492
transform 1 0 63296 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_555
timestamp 1624635492
transform 1 0 52164 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_579
timestamp 1624635492
transform 1 0 54372 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_567
timestamp 1624635492
transform 1 0 53268 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_600
timestamp 1624635492
transform 1 0 56304 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_591
timestamp 1624635492
transform 1 0 55476 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1624635492
transform 1 0 56212 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_624
timestamp 1624635492
transform 1 0 58512 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_612
timestamp 1624635492
transform 1 0 57408 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_636
timestamp 1624635492
transform 1 0 59616 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_657
timestamp 1624635492
transform 1 0 61548 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_648
timestamp 1624635492
transform 1 0 60720 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1624635492
transform 1 0 61456 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_681
timestamp 1624635492
transform 1 0 63756 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_669
timestamp 1624635492
transform 1 0 62652 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_562
timestamp 1624635492
transform 1 0 52808 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_550
timestamp 1624635492
transform 1 0 51704 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_583
timestamp 1624635492
transform 1 0 54740 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_571
timestamp 1624635492
transform 1 0 53636 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1624635492
transform 1 0 53544 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_595
timestamp 1624635492
transform 1 0 55844 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_619
timestamp 1624635492
transform 1 0 58052 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_607
timestamp 1624635492
transform 1 0 56948 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_640
timestamp 1624635492
transform 1 0 59984 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_628
timestamp 1624635492
transform 1 0 58880 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1624635492
transform 1 0 58788 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_664
timestamp 1624635492
transform 1 0 62192 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_652
timestamp 1624635492
transform 1 0 61088 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_676
timestamp 1624635492
transform 1 0 63296 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_561
timestamp 1624635492
transform 1 0 52716 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_549
timestamp 1624635492
transform 1 0 51612 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_555
timestamp 1624635492
transform 1 0 52164 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_583
timestamp 1624635492
transform 1 0 54740 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_571
timestamp 1624635492
transform 1 0 53636 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_569
timestamp 1624635492
transform 1 0 53452 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_579
timestamp 1624635492
transform 1 0 54372 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_567
timestamp 1624635492
transform 1 0 53268 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1624635492
transform 1 0 53544 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_595
timestamp 1624635492
transform 1 0 55844 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_600
timestamp 1624635492
transform 1 0 56304 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_591
timestamp 1624635492
transform 1 0 55476 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1624635492
transform 1 0 56212 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_619
timestamp 1624635492
transform 1 0 58052 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_607
timestamp 1624635492
transform 1 0 56948 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_618
timestamp 1624635492
transform 1 0 57960 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_612
timestamp 1624635492
transform 1 0 57408 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _195_
timestamp 1624635492
transform -1 0 57960 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_640
timestamp 1624635492
transform 1 0 59984 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_628
timestamp 1624635492
transform 1 0 58880 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_642
timestamp 1624635492
transform 1 0 60168 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_630
timestamp 1624635492
transform 1 0 59064 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1624635492
transform 1 0 58788 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_664
timestamp 1624635492
transform 1 0 62192 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_652
timestamp 1624635492
transform 1 0 61088 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_657
timestamp 1624635492
transform 1 0 61548 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_654
timestamp 1624635492
transform 1 0 61272 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1624635492
transform 1 0 61456 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_676
timestamp 1624635492
transform 1 0 63296 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_681
timestamp 1624635492
transform 1 0 63756 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_669
timestamp 1624635492
transform 1 0 62652 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_555
timestamp 1624635492
transform 1 0 52164 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_579
timestamp 1624635492
transform 1 0 54372 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_567
timestamp 1624635492
transform 1 0 53268 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_600
timestamp 1624635492
transform 1 0 56304 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_591
timestamp 1624635492
transform 1 0 55476 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1624635492
transform 1 0 56212 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_624
timestamp 1624635492
transform 1 0 58512 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_612
timestamp 1624635492
transform 1 0 57408 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_636
timestamp 1624635492
transform 1 0 59616 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_657
timestamp 1624635492
transform 1 0 61548 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_648
timestamp 1624635492
transform 1 0 60720 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1624635492
transform 1 0 61456 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_681
timestamp 1624635492
transform 1 0 63756 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_669
timestamp 1624635492
transform 1 0 62652 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_557
timestamp 1624635492
transform 1 0 52348 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_583
timestamp 1624635492
transform 1 0 54740 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_571
timestamp 1624635492
transform 1 0 53636 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_569
timestamp 1624635492
transform 1 0 53452 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1624635492
transform 1 0 53544 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_595
timestamp 1624635492
transform 1 0 55844 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_619
timestamp 1624635492
transform 1 0 58052 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_607
timestamp 1624635492
transform 1 0 56948 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_640
timestamp 1624635492
transform 1 0 59984 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_628
timestamp 1624635492
transform 1 0 58880 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1624635492
transform 1 0 58788 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_664
timestamp 1624635492
transform 1 0 62192 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_652
timestamp 1624635492
transform 1 0 61088 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_676
timestamp 1624635492
transform 1 0 63296 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_555
timestamp 1624635492
transform 1 0 52164 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_579
timestamp 1624635492
transform 1 0 54372 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_567
timestamp 1624635492
transform 1 0 53268 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_600
timestamp 1624635492
transform 1 0 56304 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_591
timestamp 1624635492
transform 1 0 55476 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1624635492
transform 1 0 56212 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_624
timestamp 1624635492
transform 1 0 58512 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_612
timestamp 1624635492
transform 1 0 57408 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_636
timestamp 1624635492
transform 1 0 59616 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_657
timestamp 1624635492
transform 1 0 61548 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_648
timestamp 1624635492
transform 1 0 60720 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1624635492
transform 1 0 61456 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _071_
timestamp 1624635492
transform -1 0 62468 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_673
timestamp 1624635492
transform 1 0 63020 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_667
timestamp 1624635492
transform 1 0 62468 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1624635492
transform 1 0 62836 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_562
timestamp 1624635492
transform 1 0 52808 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_550
timestamp 1624635492
transform 1 0 51704 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_583
timestamp 1624635492
transform 1 0 54740 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_571
timestamp 1624635492
transform 1 0 53636 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1624635492
transform 1 0 53544 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_595
timestamp 1624635492
transform 1 0 55844 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_622
timestamp 1624635492
transform 1 0 58328 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_619
timestamp 1624635492
transform 1 0 58052 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_607
timestamp 1624635492
transform 1 0 56948 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A1
timestamp 1624635492
transform 1 0 58144 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_640
timestamp 1624635492
transform 1 0 59984 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_628
timestamp 1624635492
transform 1 0 58880 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_626
timestamp 1624635492
transform 1 0 58696 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1624635492
transform 1 0 58788 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_664
timestamp 1624635492
transform 1 0 62192 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_652
timestamp 1624635492
transform 1 0 61088 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_676
timestamp 1624635492
transform 1 0 63296 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_555
timestamp 1624635492
transform 1 0 52164 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_579
timestamp 1624635492
transform 1 0 54372 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_567
timestamp 1624635492
transform 1 0 53268 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_600
timestamp 1624635492
transform 1 0 56304 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_591
timestamp 1624635492
transform 1 0 55476 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1624635492
transform 1 0 56212 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_620
timestamp 1624635492
transform 1 0 58144 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_612
timestamp 1624635492
transform 1 0 57408 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A2
timestamp 1624635492
transform 1 0 57960 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 58512 0 -1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_78_637
timestamp 1624635492
transform 1 0 59708 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_631
timestamp 1624635492
transform 1 0 59156 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__B1
timestamp 1624635492
transform 1 0 59524 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_657
timestamp 1624635492
transform 1 0 61548 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_655
timestamp 1624635492
transform 1 0 61364 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_649
timestamp 1624635492
transform 1 0 60812 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1624635492
transform 1 0 61456 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_681
timestamp 1624635492
transform 1 0 63756 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_669
timestamp 1624635492
transform 1 0 62652 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_562
timestamp 1624635492
transform 1 0 52808 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_550
timestamp 1624635492
transform 1 0 51704 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_583
timestamp 1624635492
transform 1 0 54740 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_571
timestamp 1624635492
transform 1 0 53636 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1624635492
transform 1 0 53544 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_595
timestamp 1624635492
transform 1 0 55844 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_620
timestamp 1624635492
transform 1 0 58144 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_79_615
timestamp 1624635492
transform 1 0 57684 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_607
timestamp 1624635492
transform 1 0 56948 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__B2
timestamp 1624635492
transform 1 0 57960 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_640
timestamp 1624635492
transform 1 0 59984 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_628
timestamp 1624635492
transform 1 0 58880 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_626
timestamp 1624635492
transform 1 0 58696 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1624635492
transform 1 0 58788 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_664
timestamp 1624635492
transform 1 0 62192 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_652
timestamp 1624635492
transform 1 0 61088 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_676
timestamp 1624635492
transform 1 0 63296 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_693
timestamp 1624635492
transform 1 0 64860 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_685
timestamp 1624635492
transform 1 0 64124 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1624635492
transform 1 0 64032 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_705
timestamp 1624635492
transform 1 0 65964 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_697
timestamp 1624635492
transform 1 0 65228 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_714
timestamp 1624635492
transform 1 0 66792 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_721
timestamp 1624635492
transform 1 0 67436 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_709
timestamp 1624635492
transform 1 0 66332 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1624635492
transform 1 0 66700 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_732
timestamp 1624635492
transform 1 0 68448 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_726
timestamp 1624635492
transform 1 0 67896 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1624635492
transform -1 0 68816 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1624635492
transform -1 0 68816 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1624635492
transform 1 0 64124 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1624635492
transform 1 0 64032 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_697
timestamp 1624635492
transform 1 0 65228 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_721
timestamp 1624635492
transform 1 0 67436 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_709
timestamp 1624635492
transform 1 0 66332 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1624635492
transform 1 0 68172 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output403
timestamp 1624635492
transform 1 0 67804 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1624635492
transform -1 0 68816 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1624635492
transform 1 0 64124 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_683
timestamp 1624635492
transform 1 0 63940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1624635492
transform 1 0 64032 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _208_
timestamp 1624635492
transform -1 0 65136 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1624635492
transform 1 0 65228 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_708
timestamp 1624635492
transform 1 0 66240 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_696
timestamp 1624635492
transform 1 0 65136 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_721
timestamp 1624635492
transform 1 0 67436 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1624635492
transform 1 0 66332 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_714
timestamp 1624635492
transform 1 0 66792 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_712
timestamp 1624635492
transform 1 0 66608 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1624635492
transform 1 0 66700 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_732
timestamp 1624635492
transform 1 0 68448 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_726
timestamp 1624635492
transform 1 0 67896 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1624635492
transform -1 0 68816 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1624635492
transform -1 0 68816 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_693
timestamp 1624635492
transform 1 0 64860 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_705
timestamp 1624635492
transform 1 0 65964 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_714
timestamp 1624635492
transform 1 0 66792 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1624635492
transform 1 0 66700 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_732
timestamp 1624635492
transform 1 0 68448 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_726
timestamp 1624635492
transform 1 0 67896 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1624635492
transform -1 0 68816 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_692
timestamp 1624635492
transform 1 0 64768 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_685
timestamp 1624635492
transform 1 0 64124 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1624635492
transform 1 0 64032 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _112_
timestamp 1624635492
transform 1 0 64492 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_704
timestamp 1624635492
transform 1 0 65872 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_716
timestamp 1624635492
transform 1 0 66976 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_732
timestamp 1624635492
transform 1 0 68448 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_728
timestamp 1624635492
transform 1 0 68080 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1624635492
transform -1 0 68816 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1624635492
transform 1 0 64124 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_693
timestamp 1624635492
transform 1 0 64860 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1624635492
transform 1 0 64032 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_697
timestamp 1624635492
transform 1 0 65228 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_705
timestamp 1624635492
transform 1 0 65964 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_717
timestamp 1624635492
transform 1 0 67068 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_709
timestamp 1624635492
transform 1 0 66332 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_714
timestamp 1624635492
transform 1 0 66792 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 67528 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1624635492
transform 1 0 66700 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1624635492
transform 1 0 68172 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_722
timestamp 1624635492
transform 1 0 67528 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_729
timestamp 1624635492
transform 1 0 68172 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1624635492
transform -1 0 68172 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1624635492
transform -1 0 68816 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1624635492
transform -1 0 68816 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _299_
timestamp 1624635492
transform -1 0 68172 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_693
timestamp 1624635492
transform 1 0 64860 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_705
timestamp 1624635492
transform 1 0 65964 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_721
timestamp 1624635492
transform 1 0 67436 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_718
timestamp 1624635492
transform 1 0 67160 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_714
timestamp 1624635492
transform 1 0 66792 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output442_A
timestamp 1624635492
transform 1 0 67252 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1624635492
transform 1 0 66700 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_729
timestamp 1624635492
transform 1 0 68172 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output442
timestamp 1624635492
transform 1 0 67804 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1624635492
transform -1 0 68816 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_693
timestamp 1624635492
transform 1 0 64860 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_685
timestamp 1624635492
transform 1 0 64124 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1624635492
transform 1 0 64032 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_705
timestamp 1624635492
transform 1 0 65964 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_697
timestamp 1624635492
transform 1 0 65228 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_714
timestamp 1624635492
transform 1 0 66792 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_721
timestamp 1624635492
transform 1 0 67436 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_709
timestamp 1624635492
transform 1 0 66332 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1624635492
transform 1 0 66700 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_732
timestamp 1624635492
transform 1 0 68448 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_726
timestamp 1624635492
transform 1 0 67896 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1624635492
transform -1 0 68816 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1624635492
transform -1 0 68816 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_685
timestamp 1624635492
transform 1 0 64124 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1624635492
transform 1 0 64032 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_697
timestamp 1624635492
transform 1 0 65228 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_721
timestamp 1624635492
transform 1 0 67436 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_709
timestamp 1624635492
transform 1 0 66332 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1624635492
transform 1 0 68172 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output404
timestamp 1624635492
transform 1 0 67804 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1624635492
transform -1 0 68816 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_693
timestamp 1624635492
transform 1 0 64860 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_705
timestamp 1624635492
transform 1 0 65964 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_714
timestamp 1624635492
transform 1 0 66792 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1624635492
transform 1 0 66700 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_732
timestamp 1624635492
transform 1 0 68448 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_726
timestamp 1624635492
transform 1 0 67896 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1624635492
transform -1 0 68816 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_693
timestamp 1624635492
transform 1 0 64860 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_685
timestamp 1624635492
transform 1 0 64124 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1624635492
transform 1 0 64032 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_705
timestamp 1624635492
transform 1 0 65964 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_697
timestamp 1624635492
transform 1 0 65228 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_714
timestamp 1624635492
transform 1 0 66792 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_721
timestamp 1624635492
transform 1 0 67436 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_709
timestamp 1624635492
transform 1 0 66332 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1624635492
transform 1 0 66700 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_732
timestamp 1624635492
transform 1 0 68448 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_726
timestamp 1624635492
transform 1 0 67896 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1624635492
transform -1 0 68816 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1624635492
transform -1 0 68816 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_685
timestamp 1624635492
transform 1 0 64124 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1624635492
transform 1 0 64032 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_697
timestamp 1624635492
transform 1 0 65228 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_717
timestamp 1624635492
transform 1 0 67068 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_709
timestamp 1624635492
transform 1 0 66332 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 67528 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1624635492
transform 1 0 68172 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_722
timestamp 1624635492
transform 1 0 67528 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1624635492
transform -1 0 68172 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1624635492
transform -1 0 68816 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_685
timestamp 1624635492
transform 1 0 64124 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_693
timestamp 1624635492
transform 1 0 64860 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1624635492
transform 1 0 64032 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_705
timestamp 1624635492
transform 1 0 65964 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_697
timestamp 1624635492
transform 1 0 65228 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_705
timestamp 1624635492
transform 1 0 65964 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _189_
timestamp 1624635492
transform -1 0 66424 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_710
timestamp 1624635492
transform 1 0 66424 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_714
timestamp 1624635492
transform 1 0 66792 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1624635492
transform 1 0 66700 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_730
timestamp 1624635492
transform 1 0 68264 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_722
timestamp 1624635492
transform 1 0 67528 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_732
timestamp 1624635492
transform 1 0 68448 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_726
timestamp 1624635492
transform 1 0 67896 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1624635492
transform -1 0 68816 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1624635492
transform -1 0 68816 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_693
timestamp 1624635492
transform 1 0 64860 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_705
timestamp 1624635492
transform 1 0 65964 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_721
timestamp 1624635492
transform 1 0 67436 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_718
timestamp 1624635492
transform 1 0 67160 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_714
timestamp 1624635492
transform 1 0 66792 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output443_A
timestamp 1624635492
transform -1 0 67436 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1624635492
transform 1 0 66700 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_729
timestamp 1624635492
transform 1 0 68172 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output443
timestamp 1624635492
transform 1 0 67804 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1624635492
transform -1 0 68816 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_685
timestamp 1624635492
transform 1 0 64124 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1624635492
transform 1 0 64032 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_697
timestamp 1624635492
transform 1 0 65228 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_721
timestamp 1624635492
transform 1 0 67436 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_709
timestamp 1624635492
transform 1 0 66332 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1624635492
transform -1 0 68816 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_685
timestamp 1624635492
transform 1 0 64124 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_693
timestamp 1624635492
transform 1 0 64860 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1624635492
transform 1 0 64032 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_697
timestamp 1624635492
transform 1 0 65228 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_705
timestamp 1624635492
transform 1 0 65964 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_721
timestamp 1624635492
transform 1 0 67436 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_709
timestamp 1624635492
transform 1 0 66332 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_714
timestamp 1624635492
transform 1 0 66792 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1624635492
transform 1 0 66700 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_729
timestamp 1624635492
transform 1 0 68172 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_722
timestamp 1624635492
transform 1 0 67528 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output405
timestamp 1624635492
transform 1 0 67804 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1624635492
transform -1 0 68816 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1624635492
transform -1 0 68816 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_685
timestamp 1624635492
transform 1 0 64124 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_700
timestamp 1624635492
transform 1 0 65504 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _146_
timestamp 1624635492
transform 1 0 65228 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_714
timestamp 1624635492
transform 1 0 66792 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_712
timestamp 1624635492
transform 1 0 66608 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1624635492
transform 1 0 66700 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_732
timestamp 1624635492
transform 1 0 68448 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_726
timestamp 1624635492
transform 1 0 67896 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1624635492
transform -1 0 68816 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_693
timestamp 1624635492
transform 1 0 64860 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_685
timestamp 1624635492
transform 1 0 64124 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1624635492
transform 1 0 64032 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_705
timestamp 1624635492
transform 1 0 65964 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_697
timestamp 1624635492
transform 1 0 65228 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_714
timestamp 1624635492
transform 1 0 66792 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_721
timestamp 1624635492
transform 1 0 67436 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_709
timestamp 1624635492
transform 1 0 66332 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1624635492
transform 1 0 66700 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_732
timestamp 1624635492
transform 1 0 68448 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_726
timestamp 1624635492
transform 1 0 67896 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1624635492
transform -1 0 68816 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1624635492
transform -1 0 68816 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_685
timestamp 1624635492
transform 1 0 64124 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1624635492
transform 1 0 64032 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_697
timestamp 1624635492
transform 1 0 65228 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_717
timestamp 1624635492
transform 1 0 67068 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_709
timestamp 1624635492
transform 1 0 66332 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 67528 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1624635492
transform 1 0 68172 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_722
timestamp 1624635492
transform 1 0 67528 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1624635492
transform -1 0 68172 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1624635492
transform -1 0 68816 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_11
timestamp 1624635492
transform 1 0 2116 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1624635492
transform 1 0 1380 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output426
timestamp 1624635492
transform -1 0 2116 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1624635492
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_17
timestamp 1624635492
transform 1 0 2668 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output426_A
timestamp 1624635492
transform -1 0 2668 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1624635492
transform 1 0 3772 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_42
timestamp 1624635492
transform 1 0 4968 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_30
timestamp 1624635492
transform 1 0 3864 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_54
timestamp 1624635492
transform 1 0 6072 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_66
timestamp 1624635492
transform 1 0 7176 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_87
timestamp 1624635492
transform 1 0 9108 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_78
timestamp 1624635492
transform 1 0 8280 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1624635492
transform 1 0 9016 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_99
timestamp 1624635492
transform 1 0 10212 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_111
timestamp 1624635492
transform 1 0 11316 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_123
timestamp 1624635492
transform 1 0 12420 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_135
timestamp 1624635492
transform 1 0 13524 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_7
timestamp 1624635492
transform 1 0 1748 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1624635492
transform 1 0 1380 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 1748 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1624635492
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_19
timestamp 1624635492
transform 1 0 2852 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_43
timestamp 1624635492
transform 1 0 5060 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_31
timestamp 1624635492
transform 1 0 3956 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_58
timestamp 1624635492
transform 1 0 6440 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_55
timestamp 1624635492
transform 1 0 6164 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1624635492
transform 1 0 6348 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_71
timestamp 1624635492
transform 1 0 7636 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_66
timestamp 1624635492
transform 1 0 7176 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _270_
timestamp 1624635492
transform 1 0 7360 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_83
timestamp 1624635492
transform 1 0 8740 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_95
timestamp 1624635492
transform 1 0 9844 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_115
timestamp 1624635492
transform 1 0 11684 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_113
timestamp 1624635492
transform 1 0 11500 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_107
timestamp 1624635492
transform 1 0 10948 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1624635492
transform 1 0 11592 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_127
timestamp 1624635492
transform 1 0 12788 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1624635492
transform 1 0 1380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_11
timestamp 1624635492
transform 1 0 2116 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1624635492
transform 1 0 1380 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1624635492
transform 1 0 1748 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1624635492
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1624635492
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1624635492
transform 1 0 3588 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1624635492
transform 1 0 2484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_23
timestamp 1624635492
transform 1 0 3220 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1624635492
transform 1 0 3772 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1624635492
transform 1 0 4692 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_42
timestamp 1624635492
transform 1 0 4968 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_30
timestamp 1624635492
transform 1 0 3864 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_58
timestamp 1624635492
transform 1 0 6440 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_51
timestamp 1624635492
transform 1 0 5796 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_54
timestamp 1624635492
transform 1 0 6072 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1624635492
transform 1 0 6348 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_70
timestamp 1624635492
transform 1 0 7544 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_66
timestamp 1624635492
transform 1 0 7176 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_82
timestamp 1624635492
transform 1 0 8648 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_87
timestamp 1624635492
transform 1 0 9108 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_78
timestamp 1624635492
transform 1 0 8280 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1624635492
transform 1 0 9016 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_94
timestamp 1624635492
transform 1 0 9752 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_99
timestamp 1624635492
transform 1 0 10212 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_115
timestamp 1624635492
transform 1 0 11684 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_106
timestamp 1624635492
transform 1 0 10856 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_111
timestamp 1624635492
transform 1 0 11316 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1624635492
transform 1 0 11592 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_127
timestamp 1624635492
transform 1 0 12788 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_123
timestamp 1624635492
transform 1 0 12420 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_135
timestamp 1624635492
transform 1 0 13524 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1624635492
transform 1 0 1380 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1624635492
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_27
timestamp 1624635492
transform 1 0 3588 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1624635492
transform 1 0 2484 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1624635492
transform 1 0 3772 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_42
timestamp 1624635492
transform 1 0 4968 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_30
timestamp 1624635492
transform 1 0 3864 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_54
timestamp 1624635492
transform 1 0 6072 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_66
timestamp 1624635492
transform 1 0 7176 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_87
timestamp 1624635492
transform 1 0 9108 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_78
timestamp 1624635492
transform 1 0 8280 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1624635492
transform 1 0 9016 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_99
timestamp 1624635492
transform 1 0 10212 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_111
timestamp 1624635492
transform 1 0 11316 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_123
timestamp 1624635492
transform 1 0 12420 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_135
timestamp 1624635492
transform 1 0 13524 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1624635492
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1624635492
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1624635492
transform 1 0 3588 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1624635492
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1624635492
transform 1 0 4692 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_58
timestamp 1624635492
transform 1 0 6440 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_51
timestamp 1624635492
transform 1 0 5796 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1624635492
transform 1 0 6348 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_70
timestamp 1624635492
transform 1 0 7544 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_82
timestamp 1624635492
transform 1 0 8648 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_94
timestamp 1624635492
transform 1 0 9752 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_115
timestamp 1624635492
transform 1 0 11684 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_106
timestamp 1624635492
transform 1 0 10856 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1624635492
transform 1 0 11592 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_127
timestamp 1624635492
transform 1 0 12788 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1624635492
transform 1 0 1380 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1624635492
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_27
timestamp 1624635492
transform 1 0 3588 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1624635492
transform 1 0 2484 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1624635492
transform 1 0 3772 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_42
timestamp 1624635492
transform 1 0 4968 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_30
timestamp 1624635492
transform 1 0 3864 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_54
timestamp 1624635492
transform 1 0 6072 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_66
timestamp 1624635492
transform 1 0 7176 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_87
timestamp 1624635492
transform 1 0 9108 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_78
timestamp 1624635492
transform 1 0 8280 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1624635492
transform 1 0 9016 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_99
timestamp 1624635492
transform 1 0 10212 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_111
timestamp 1624635492
transform 1 0 11316 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_123
timestamp 1624635492
transform 1 0 12420 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_135
timestamp 1624635492
transform 1 0 13524 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_87_11
timestamp 1624635492
transform 1 0 2116 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_3
timestamp 1624635492
transform 1 0 1380 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output387
timestamp 1624635492
transform -1 0 2116 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1624635492
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_29
timestamp 1624635492
transform 1 0 3772 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_17
timestamp 1624635492
transform 1 0 2668 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output387_A
timestamp 1624635492
transform -1 0 2668 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_41
timestamp 1624635492
transform 1 0 4876 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_58
timestamp 1624635492
transform 1 0 6440 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_53
timestamp 1624635492
transform 1 0 5980 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1624635492
transform 1 0 6348 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_70
timestamp 1624635492
transform 1 0 7544 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_82
timestamp 1624635492
transform 1 0 8648 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_94
timestamp 1624635492
transform 1 0 9752 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_115
timestamp 1624635492
transform 1 0 11684 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_106
timestamp 1624635492
transform 1 0 10856 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1624635492
transform 1 0 11592 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_127
timestamp 1624635492
transform 1 0 12788 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_11
timestamp 1624635492
transform 1 0 2116 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_3
timestamp 1624635492
transform 1 0 1380 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1624635492
transform 1 0 1380 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output425
timestamp 1624635492
transform -1 0 2116 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1624635492
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1624635492
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_29
timestamp 1624635492
transform 1 0 3772 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_17
timestamp 1624635492
transform 1 0 2668 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_25
timestamp 1624635492
transform 1 0 3404 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_21
timestamp 1624635492
transform 1 0 3036 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_15
timestamp 1624635492
transform 1 0 2484 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output425_A
timestamp 1624635492
transform 1 0 2484 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1624635492
transform 1 0 3772 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _133_
timestamp 1624635492
transform -1 0 3404 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_41
timestamp 1624635492
transform 1 0 4876 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_42
timestamp 1624635492
transform 1 0 4968 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_30
timestamp 1624635492
transform 1 0 3864 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_58
timestamp 1624635492
transform 1 0 6440 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_53
timestamp 1624635492
transform 1 0 5980 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_54
timestamp 1624635492
transform 1 0 6072 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1624635492
transform 1 0 6348 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_70
timestamp 1624635492
transform 1 0 7544 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_66
timestamp 1624635492
transform 1 0 7176 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_82
timestamp 1624635492
transform 1 0 8648 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_87
timestamp 1624635492
transform 1 0 9108 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_78
timestamp 1624635492
transform 1 0 8280 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1624635492
transform 1 0 9016 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_94
timestamp 1624635492
transform 1 0 9752 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_99
timestamp 1624635492
transform 1 0 10212 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_115
timestamp 1624635492
transform 1 0 11684 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_106
timestamp 1624635492
transform 1 0 10856 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_111
timestamp 1624635492
transform 1 0 11316 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1624635492
transform 1 0 11592 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_127
timestamp 1624635492
transform 1 0 12788 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_123
timestamp 1624635492
transform 1 0 12420 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_135
timestamp 1624635492
transform 1 0 13524 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1624635492
transform 1 0 1380 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1624635492
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_90_27
timestamp 1624635492
transform 1 0 3588 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1624635492
transform 1 0 2484 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1624635492
transform 1 0 3772 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_42
timestamp 1624635492
transform 1 0 4968 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_30
timestamp 1624635492
transform 1 0 3864 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_54
timestamp 1624635492
transform 1 0 6072 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_66
timestamp 1624635492
transform 1 0 7176 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_87
timestamp 1624635492
transform 1 0 9108 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_78
timestamp 1624635492
transform 1 0 8280 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1624635492
transform 1 0 9016 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_99
timestamp 1624635492
transform 1 0 10212 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_111
timestamp 1624635492
transform 1 0 11316 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_123
timestamp 1624635492
transform 1 0 12420 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_135
timestamp 1624635492
transform 1 0 13524 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1624635492
transform 1 0 1380 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1624635492
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1624635492
transform 1 0 3588 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1624635492
transform 1 0 2484 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_39
timestamp 1624635492
transform 1 0 4692 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_58
timestamp 1624635492
transform 1 0 6440 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_51
timestamp 1624635492
transform 1 0 5796 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1624635492
transform 1 0 6348 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_70
timestamp 1624635492
transform 1 0 7544 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_82
timestamp 1624635492
transform 1 0 8648 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_94
timestamp 1624635492
transform 1 0 9752 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_115
timestamp 1624635492
transform 1 0 11684 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_106
timestamp 1624635492
transform 1 0 10856 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1624635492
transform 1 0 11592 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_127
timestamp 1624635492
transform 1 0 12788 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_12
timestamp 1624635492
transform 1 0 2208 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_6
timestamp 1624635492
transform 1 0 1656 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 2208 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1624635492
transform -1 0 1656 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1624635492
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_92_28
timestamp 1624635492
transform 1 0 3680 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_24
timestamp 1624635492
transform 1 0 3312 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1624635492
transform 1 0 3772 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_42
timestamp 1624635492
transform 1 0 4968 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_30
timestamp 1624635492
transform 1 0 3864 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_54
timestamp 1624635492
transform 1 0 6072 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_66
timestamp 1624635492
transform 1 0 7176 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_87
timestamp 1624635492
transform 1 0 9108 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_78
timestamp 1624635492
transform 1 0 8280 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1624635492
transform 1 0 9016 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_99
timestamp 1624635492
transform 1 0 10212 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_111
timestamp 1624635492
transform 1 0 11316 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_123
timestamp 1624635492
transform 1 0 12420 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_135
timestamp 1624635492
transform 1 0 13524 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1624635492
transform 1 0 1380 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1624635492
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1624635492
transform 1 0 3588 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1624635492
transform 1 0 2484 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1624635492
transform 1 0 4692 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_58
timestamp 1624635492
transform 1 0 6440 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_51
timestamp 1624635492
transform 1 0 5796 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1624635492
transform 1 0 6348 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_70
timestamp 1624635492
transform 1 0 7544 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_82
timestamp 1624635492
transform 1 0 8648 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_94
timestamp 1624635492
transform 1 0 9752 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_115
timestamp 1624635492
transform 1 0 11684 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_106
timestamp 1624635492
transform 1 0 10856 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1624635492
transform 1 0 11592 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_127
timestamp 1624635492
transform 1 0 12788 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1624635492
transform 1 0 1380 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1624635492
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_27
timestamp 1624635492
transform 1 0 3588 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1624635492
transform 1 0 2484 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1624635492
transform 1 0 3772 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_42
timestamp 1624635492
transform 1 0 4968 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_30
timestamp 1624635492
transform 1 0 3864 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_54
timestamp 1624635492
transform 1 0 6072 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_73
timestamp 1624635492
transform 1 0 7820 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_66
timestamp 1624635492
transform 1 0 7176 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _322_
timestamp 1624635492
transform 1 0 7544 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_87
timestamp 1624635492
transform 1 0 9108 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_85
timestamp 1624635492
transform 1 0 8924 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1624635492
transform 1 0 9016 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_99
timestamp 1624635492
transform 1 0 10212 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_111
timestamp 1624635492
transform 1 0 11316 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_123
timestamp 1624635492
transform 1 0 12420 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_135
timestamp 1624635492
transform 1 0 13524 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1624635492
transform 1 0 1380 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1624635492
transform 1 0 1380 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1624635492
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1624635492
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_27
timestamp 1624635492
transform 1 0 3588 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1624635492
transform 1 0 2484 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1624635492
transform 1 0 3588 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1624635492
transform 1 0 2484 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1624635492
transform 1 0 3772 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_42
timestamp 1624635492
transform 1 0 4968 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_30
timestamp 1624635492
transform 1 0 3864 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_39
timestamp 1624635492
transform 1 0 4692 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_54
timestamp 1624635492
transform 1 0 6072 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_58
timestamp 1624635492
transform 1 0 6440 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_56
timestamp 1624635492
transform 1 0 6256 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_50
timestamp 1624635492
transform 1 0 5704 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1624635492
transform 1 0 6348 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _148_
timestamp 1624635492
transform 1 0 5428 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_66
timestamp 1624635492
transform 1 0 7176 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_70
timestamp 1624635492
transform 1 0 7544 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_87
timestamp 1624635492
transform 1 0 9108 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_78
timestamp 1624635492
transform 1 0 8280 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_82
timestamp 1624635492
transform 1 0 8648 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1624635492
transform 1 0 9016 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_99
timestamp 1624635492
transform 1 0 10212 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_94
timestamp 1624635492
transform 1 0 9752 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_111
timestamp 1624635492
transform 1 0 11316 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_115
timestamp 1624635492
transform 1 0 11684 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_106
timestamp 1624635492
transform 1 0 10856 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1624635492
transform 1 0 11592 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_123
timestamp 1624635492
transform 1 0 12420 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_127
timestamp 1624635492
transform 1 0 12788 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_135
timestamp 1624635492
transform 1 0 13524 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_97_11
timestamp 1624635492
transform 1 0 2116 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_3
timestamp 1624635492
transform 1 0 1380 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output386
timestamp 1624635492
transform -1 0 2116 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1624635492
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_29
timestamp 1624635492
transform 1 0 3772 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_17
timestamp 1624635492
transform 1 0 2668 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output386_A
timestamp 1624635492
transform 1 0 2484 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_41
timestamp 1624635492
transform 1 0 4876 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_58
timestamp 1624635492
transform 1 0 6440 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_53
timestamp 1624635492
transform 1 0 5980 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1624635492
transform 1 0 6348 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_70
timestamp 1624635492
transform 1 0 7544 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_82
timestamp 1624635492
transform 1 0 8648 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_100
timestamp 1624635492
transform 1 0 10304 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_94
timestamp 1624635492
transform 1 0 9752 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1624635492
transform 1 0 10120 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_115
timestamp 1624635492
transform 1 0 11684 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_112
timestamp 1624635492
transform 1 0 11408 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1624635492
transform 1 0 11592 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_127
timestamp 1624635492
transform 1 0 12788 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1624635492
transform 1 0 1380 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1624635492
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_27
timestamp 1624635492
transform 1 0 3588 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1624635492
transform 1 0 2484 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1624635492
transform 1 0 3772 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_42
timestamp 1624635492
transform 1 0 4968 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_30
timestamp 1624635492
transform 1 0 3864 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_54
timestamp 1624635492
transform 1 0 6072 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_66
timestamp 1624635492
transform 1 0 7176 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_87
timestamp 1624635492
transform 1 0 9108 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_78
timestamp 1624635492
transform 1 0 8280 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1624635492
transform 1 0 9016 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_98
timestamp 1624635492
transform 1 0 10120 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_4  _091_
timestamp 1624635492
transform -1 0 10120 0 -1 56032
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_98_109
timestamp 1624635492
transform 1 0 11132 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _198_
timestamp 1624635492
transform 1 0 10856 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_131
timestamp 1624635492
transform 1 0 13156 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_127
timestamp 1624635492
transform 1 0 12788 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_121
timestamp 1624635492
transform 1 0 12236 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _179_
timestamp 1624635492
transform 1 0 12880 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_11
timestamp 1624635492
transform 1 0 2116 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_3
timestamp 1624635492
transform 1 0 1380 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output424
timestamp 1624635492
transform -1 0 2116 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1624635492
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_29
timestamp 1624635492
transform 1 0 3772 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_17
timestamp 1624635492
transform 1 0 2668 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output424_A
timestamp 1624635492
transform -1 0 2668 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_41
timestamp 1624635492
transform 1 0 4876 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_58
timestamp 1624635492
transform 1 0 6440 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_53
timestamp 1624635492
transform 1 0 5980 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1247
timestamp 1624635492
transform 1 0 6348 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_70
timestamp 1624635492
transform 1 0 7544 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_82
timestamp 1624635492
transform 1 0 8648 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_94
timestamp 1624635492
transform 1 0 9752 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_115
timestamp 1624635492
transform 1 0 11684 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_106
timestamp 1624635492
transform 1 0 10856 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1248
timestamp 1624635492
transform 1 0 11592 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_127
timestamp 1624635492
transform 1 0 12788 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1624635492
transform 1 0 1380 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1624635492
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_27
timestamp 1624635492
transform 1 0 3588 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1624635492
transform 1 0 2484 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1259
timestamp 1624635492
transform 1 0 3772 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_42
timestamp 1624635492
transform 1 0 4968 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_30
timestamp 1624635492
transform 1 0 3864 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_54
timestamp 1624635492
transform 1 0 6072 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_66
timestamp 1624635492
transform 1 0 7176 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_87
timestamp 1624635492
transform 1 0 9108 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_78
timestamp 1624635492
transform 1 0 8280 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1260
timestamp 1624635492
transform 1 0 9016 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_99
timestamp 1624635492
transform 1 0 10212 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _170_
timestamp 1624635492
transform 1 0 10580 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_118
timestamp 1624635492
transform 1 0 11960 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_106
timestamp 1624635492
transform 1 0 10856 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_130
timestamp 1624635492
transform 1 0 13064 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_12
timestamp 1624635492
transform 1 0 2208 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_6
timestamp 1624635492
transform 1 0 1656 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 2208 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1624635492
transform -1 0 1656 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1624635492
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_24
timestamp 1624635492
transform 1 0 3312 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_36
timestamp 1624635492
transform 1 0 4416 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_58
timestamp 1624635492
transform 1 0 6440 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_56
timestamp 1624635492
transform 1 0 6256 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_48
timestamp 1624635492
transform 1 0 5520 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1272
timestamp 1624635492
transform 1 0 6348 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_64
timestamp 1624635492
transform 1 0 6992 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A3
timestamp 1624635492
transform 1 0 6808 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_88
timestamp 1624635492
transform 1 0 9200 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_76
timestamp 1624635492
transform 1 0 8096 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_100
timestamp 1624635492
transform 1 0 10304 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_115
timestamp 1624635492
transform 1 0 11684 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_112
timestamp 1624635492
transform 1 0 11408 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1273
timestamp 1624635492
transform 1 0 11592 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_127
timestamp 1624635492
transform 1 0 12788 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1624635492
transform 1 0 1380 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1624635492
transform 1 0 1380 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1624635492
transform 1 0 1104 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1624635492
transform 1 0 1104 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_27
timestamp 1624635492
transform 1 0 3588 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_15
timestamp 1624635492
transform 1 0 2484 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_27
timestamp 1624635492
transform 1 0 3588 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1624635492
transform 1 0 2484 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1284
timestamp 1624635492
transform 1 0 3772 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_39
timestamp 1624635492
transform 1 0 4692 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_40
timestamp 1624635492
transform 1 0 4784 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_102_30
timestamp 1624635492
transform 1 0 3864 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B1
timestamp 1624635492
transform 1 0 4600 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_4  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 6440 0 -1 58208
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_103_58
timestamp 1624635492
transform 1 0 6440 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_51
timestamp 1624635492
transform 1 0 5796 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_102_58
timestamp 1624635492
transform 1 0 6440 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1297
timestamp 1624635492
transform 1 0 6348 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_70
timestamp 1624635492
transform 1 0 7544 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_74
timestamp 1624635492
transform 1 0 7912 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_70
timestamp 1624635492
transform 1 0 7544 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_64
timestamp 1624635492
transform 1 0 6992 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A2
timestamp 1624635492
transform 1 0 7360 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A1
timestamp 1624635492
transform 1 0 6808 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_82
timestamp 1624635492
transform 1 0 8648 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_87
timestamp 1624635492
transform 1 0 9108 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_78
timestamp 1624635492
transform 1 0 8280 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1285
timestamp 1624635492
transform 1 0 9016 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _234_
timestamp 1624635492
transform 1 0 8004 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_94
timestamp 1624635492
transform 1 0 9752 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_99
timestamp 1624635492
transform 1 0 10212 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_115
timestamp 1624635492
transform 1 0 11684 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_106
timestamp 1624635492
transform 1 0 10856 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_111
timestamp 1624635492
transform 1 0 11316 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1298
timestamp 1624635492
transform 1 0 11592 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_127
timestamp 1624635492
transform 1 0 12788 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_123
timestamp 1624635492
transform 1 0 12420 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_135
timestamp 1624635492
transform 1 0 13524 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1624635492
transform 1 0 1380 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1624635492
transform 1 0 1104 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_104_27
timestamp 1624635492
transform 1 0 3588 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1624635492
transform 1 0 2484 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1309
timestamp 1624635492
transform 1 0 3772 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_42
timestamp 1624635492
transform 1 0 4968 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_30
timestamp 1624635492
transform 1 0 3864 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_54
timestamp 1624635492
transform 1 0 6072 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_66
timestamp 1624635492
transform 1 0 7176 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_87
timestamp 1624635492
transform 1 0 9108 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_78
timestamp 1624635492
transform 1 0 8280 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1310
timestamp 1624635492
transform 1 0 9016 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_103
timestamp 1624635492
transform 1 0 10580 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_99
timestamp 1624635492
transform 1 0 10212 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _143_
timestamp 1624635492
transform 1 0 10304 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_115
timestamp 1624635492
transform 1 0 11684 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_133
timestamp 1624635492
transform 1 0 13340 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_127
timestamp 1624635492
transform 1 0 12788 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _313_
timestamp 1624635492
transform -1 0 13708 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1624635492
transform 1 0 1380 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1624635492
transform 1 0 1104 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1624635492
transform 1 0 3588 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1624635492
transform 1 0 2484 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1624635492
transform 1 0 4692 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_58
timestamp 1624635492
transform 1 0 6440 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_51
timestamp 1624635492
transform 1 0 5796 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1322
timestamp 1624635492
transform 1 0 6348 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_70
timestamp 1624635492
transform 1 0 7544 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_82
timestamp 1624635492
transform 1 0 8648 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_94
timestamp 1624635492
transform 1 0 9752 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_115
timestamp 1624635492
transform 1 0 11684 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_106
timestamp 1624635492
transform 1 0 10856 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1323
timestamp 1624635492
transform 1 0 11592 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_127
timestamp 1624635492
transform 1 0 12788 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_11
timestamp 1624635492
transform 1 0 2116 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_3
timestamp 1624635492
transform 1 0 1380 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output385
timestamp 1624635492
transform -1 0 2116 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1624635492
transform 1 0 1104 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_17
timestamp 1624635492
transform 1 0 2668 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output385_A
timestamp 1624635492
transform 1 0 2484 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1334
timestamp 1624635492
transform 1 0 3772 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_42
timestamp 1624635492
transform 1 0 4968 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_30
timestamp 1624635492
transform 1 0 3864 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_54
timestamp 1624635492
transform 1 0 6072 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_66
timestamp 1624635492
transform 1 0 7176 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_87
timestamp 1624635492
transform 1 0 9108 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_78
timestamp 1624635492
transform 1 0 8280 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1335
timestamp 1624635492
transform 1 0 9016 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_99
timestamp 1624635492
transform 1 0 10212 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_111
timestamp 1624635492
transform 1 0 11316 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_123
timestamp 1624635492
transform 1 0 12420 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_135
timestamp 1624635492
transform 1 0 13524 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1624635492
transform 1 0 15456 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1624635492
transform 1 0 14352 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1624635492
transform 1 0 14260 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1624635492
transform 1 0 16560 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_192
timestamp 1624635492
transform 1 0 18768 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1624635492
transform 1 0 17664 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_213
timestamp 1624635492
transform 1 0 20700 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_201
timestamp 1624635492
transform 1 0 19596 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1624635492
transform 1 0 19504 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_225
timestamp 1624635492
transform 1 0 21804 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_249
timestamp 1624635492
transform 1 0 24012 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_237
timestamp 1624635492
transform 1 0 22908 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_270
timestamp 1624635492
transform 1 0 25944 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_258
timestamp 1624635492
transform 1 0 24840 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1624635492
transform 1 0 24748 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_151
timestamp 1624635492
transform 1 0 14996 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_139
timestamp 1624635492
transform 1 0 13892 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_172
timestamp 1624635492
transform 1 0 16928 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_163
timestamp 1624635492
transform 1 0 16100 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1624635492
transform 1 0 16836 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_196
timestamp 1624635492
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_184
timestamp 1624635492
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_208
timestamp 1624635492
transform 1 0 20240 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_229
timestamp 1624635492
transform 1 0 22172 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_220
timestamp 1624635492
transform 1 0 21344 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_216
timestamp 1624635492
transform 1 0 20976 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1624635492
transform 1 0 22080 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _105_
timestamp 1624635492
transform 1 0 21068 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_253
timestamp 1624635492
transform 1 0 24380 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_241
timestamp 1624635492
transform 1 0 23276 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_265
timestamp 1624635492
transform 1 0 25484 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_151
timestamp 1624635492
transform 1 0 14996 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_139
timestamp 1624635492
transform 1 0 13892 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_156
timestamp 1624635492
transform 1 0 15456 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_144
timestamp 1624635492
transform 1 0 14352 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1624635492
transform 1 0 14260 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_172
timestamp 1624635492
transform 1 0 16928 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_163
timestamp 1624635492
transform 1 0 16100 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_168
timestamp 1624635492
transform 1 0 16560 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1624635492
transform 1 0 16836 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_196
timestamp 1624635492
transform 1 0 19136 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_184
timestamp 1624635492
transform 1 0 18032 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_192
timestamp 1624635492
transform 1 0 18768 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_180
timestamp 1624635492
transform 1 0 17664 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_208
timestamp 1624635492
transform 1 0 20240 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_213
timestamp 1624635492
transform 1 0 20700 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_201
timestamp 1624635492
transform 1 0 19596 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1624635492
transform 1 0 19504 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_229
timestamp 1624635492
transform 1 0 22172 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_220
timestamp 1624635492
transform 1 0 21344 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1624635492
transform 1 0 21804 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1624635492
transform 1 0 22080 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_253
timestamp 1624635492
transform 1 0 24380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_241
timestamp 1624635492
transform 1 0 23276 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_249
timestamp 1624635492
transform 1 0 24012 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1624635492
transform 1 0 22908 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_265
timestamp 1624635492
transform 1 0 25484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_272
timestamp 1624635492
transform 1 0 26128 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_265
timestamp 1624635492
transform 1 0 25484 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_258
timestamp 1624635492
transform 1 0 24840 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1624635492
transform 1 0 24748 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _233_
timestamp 1624635492
transform 1 0 25852 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _229_
timestamp 1624635492
transform 1 0 25208 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_156
timestamp 1624635492
transform 1 0 15456 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_144
timestamp 1624635492
transform 1 0 14352 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1624635492
transform 1 0 14260 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_168
timestamp 1624635492
transform 1 0 16560 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_192
timestamp 1624635492
transform 1 0 18768 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_180
timestamp 1624635492
transform 1 0 17664 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_213
timestamp 1624635492
transform 1 0 20700 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_201
timestamp 1624635492
transform 1 0 19596 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1624635492
transform 1 0 19504 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_225
timestamp 1624635492
transform 1 0 21804 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_249
timestamp 1624635492
transform 1 0 24012 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_237
timestamp 1624635492
transform 1 0 22908 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_270
timestamp 1624635492
transform 1 0 25944 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_258
timestamp 1624635492
transform 1 0 24840 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1624635492
transform 1 0 24748 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_151
timestamp 1624635492
transform 1 0 14996 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_139
timestamp 1624635492
transform 1 0 13892 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_172
timestamp 1624635492
transform 1 0 16928 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_163
timestamp 1624635492
transform 1 0 16100 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1624635492
transform 1 0 16836 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_196
timestamp 1624635492
transform 1 0 19136 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_184
timestamp 1624635492
transform 1 0 18032 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_208
timestamp 1624635492
transform 1 0 20240 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_229
timestamp 1624635492
transform 1 0 22172 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_220
timestamp 1624635492
transform 1 0 21344 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1624635492
transform 1 0 22080 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_253
timestamp 1624635492
transform 1 0 24380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_241
timestamp 1624635492
transform 1 0 23276 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_265
timestamp 1624635492
transform 1 0 25484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_156
timestamp 1624635492
transform 1 0 15456 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_144
timestamp 1624635492
transform 1 0 14352 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1624635492
transform 1 0 14260 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_168
timestamp 1624635492
transform 1 0 16560 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_192
timestamp 1624635492
transform 1 0 18768 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_180
timestamp 1624635492
transform 1 0 17664 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_213
timestamp 1624635492
transform 1 0 20700 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_201
timestamp 1624635492
transform 1 0 19596 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1624635492
transform 1 0 19504 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_225
timestamp 1624635492
transform 1 0 21804 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_249
timestamp 1624635492
transform 1 0 24012 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_237
timestamp 1624635492
transform 1 0 22908 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_270
timestamp 1624635492
transform 1 0 25944 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_258
timestamp 1624635492
transform 1 0 24840 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1624635492
transform 1 0 24748 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_151
timestamp 1624635492
transform 1 0 14996 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_139
timestamp 1624635492
transform 1 0 13892 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_172
timestamp 1624635492
transform 1 0 16928 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_163
timestamp 1624635492
transform 1 0 16100 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1624635492
transform 1 0 16836 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_196
timestamp 1624635492
transform 1 0 19136 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_184
timestamp 1624635492
transform 1 0 18032 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_215
timestamp 1624635492
transform 1 0 20884 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 20884 0 1 49504
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_87_229
timestamp 1624635492
transform 1 0 22172 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_227
timestamp 1624635492
transform 1 0 21988 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_221
timestamp 1624635492
transform 1 0 21436 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1624635492
transform 1 0 21252 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1624635492
transform 1 0 22080 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_253
timestamp 1624635492
transform 1 0 24380 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_241
timestamp 1624635492
transform 1 0 23276 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_265
timestamp 1624635492
transform 1 0 25484 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_151
timestamp 1624635492
transform 1 0 14996 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_139
timestamp 1624635492
transform 1 0 13892 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_156
timestamp 1624635492
transform 1 0 15456 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_144
timestamp 1624635492
transform 1 0 14352 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1624635492
transform 1 0 14260 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_172
timestamp 1624635492
transform 1 0 16928 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_163
timestamp 1624635492
transform 1 0 16100 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_168
timestamp 1624635492
transform 1 0 16560 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1624635492
transform 1 0 16836 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _052_
timestamp 1624635492
transform -1 0 18124 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_89_191
timestamp 1624635492
transform 1 0 18676 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_185
timestamp 1624635492
transform 1 0 18124 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_192
timestamp 1624635492
transform 1 0 18768 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_180
timestamp 1624635492
transform 1 0 17664 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__A
timestamp 1624635492
transform 1 0 18492 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_215
timestamp 1624635492
transform 1 0 20884 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_203
timestamp 1624635492
transform 1 0 19780 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_213
timestamp 1624635492
transform 1 0 20700 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_201
timestamp 1624635492
transform 1 0 19596 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1624635492
transform 1 0 19504 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_229
timestamp 1624635492
transform 1 0 22172 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_227
timestamp 1624635492
transform 1 0 21988 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_225
timestamp 1624635492
transform 1 0 21804 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1624635492
transform 1 0 22080 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_253
timestamp 1624635492
transform 1 0 24380 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_241
timestamp 1624635492
transform 1 0 23276 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_254
timestamp 1624635492
transform 1 0 24472 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_242
timestamp 1624635492
transform 1 0 23368 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_237
timestamp 1624635492
transform 1 0 22908 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _297_
timestamp 1624635492
transform 1 0 23092 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_265
timestamp 1624635492
transform 1 0 25484 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_270
timestamp 1624635492
transform 1 0 25944 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_258
timestamp 1624635492
transform 1 0 24840 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1624635492
transform 1 0 24748 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_155
timestamp 1624635492
transform 1 0 15364 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_148
timestamp 1624635492
transform 1 0 14720 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_144
timestamp 1624635492
transform 1 0 14352 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1624635492
transform 1 0 14260 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _070_
timestamp 1624635492
transform -1 0 15364 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_173
timestamp 1624635492
transform 1 0 17020 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_161
timestamp 1624635492
transform 1 0 15916 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1624635492
transform 1 0 15732 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_90_185
timestamp 1624635492
transform 1 0 18124 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_213
timestamp 1624635492
transform 1 0 20700 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_201
timestamp 1624635492
transform 1 0 19596 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_197
timestamp 1624635492
transform 1 0 19228 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1624635492
transform 1 0 19504 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_225
timestamp 1624635492
transform 1 0 21804 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_249
timestamp 1624635492
transform 1 0 24012 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_237
timestamp 1624635492
transform 1 0 22908 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_270
timestamp 1624635492
transform 1 0 25944 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_258
timestamp 1624635492
transform 1 0 24840 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1624635492
transform 1 0 24748 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_151
timestamp 1624635492
transform 1 0 14996 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_91_139
timestamp 1624635492
transform 1 0 13892 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_172
timestamp 1624635492
transform 1 0 16928 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_169
timestamp 1624635492
transform 1 0 16652 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_161
timestamp 1624635492
transform 1 0 15916 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_157
timestamp 1624635492
transform 1 0 15548 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1624635492
transform 1 0 16836 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _104_
timestamp 1624635492
transform 1 0 15640 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_196
timestamp 1624635492
transform 1 0 19136 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_184
timestamp 1624635492
transform 1 0 18032 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_208
timestamp 1624635492
transform 1 0 20240 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_229
timestamp 1624635492
transform 1 0 22172 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_220
timestamp 1624635492
transform 1 0 21344 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1624635492
transform 1 0 22080 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_253
timestamp 1624635492
transform 1 0 24380 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_241
timestamp 1624635492
transform 1 0 23276 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_265
timestamp 1624635492
transform 1 0 25484 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_156
timestamp 1624635492
transform 1 0 15456 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_144
timestamp 1624635492
transform 1 0 14352 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1624635492
transform 1 0 14260 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_168
timestamp 1624635492
transform 1 0 16560 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_192
timestamp 1624635492
transform 1 0 18768 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_180
timestamp 1624635492
transform 1 0 17664 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_213
timestamp 1624635492
transform 1 0 20700 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_201
timestamp 1624635492
transform 1 0 19596 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1624635492
transform 1 0 19504 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_225
timestamp 1624635492
transform 1 0 21804 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_249
timestamp 1624635492
transform 1 0 24012 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_237
timestamp 1624635492
transform 1 0 22908 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_270
timestamp 1624635492
transform 1 0 25944 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_258
timestamp 1624635492
transform 1 0 24840 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1624635492
transform 1 0 24748 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_151
timestamp 1624635492
transform 1 0 14996 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_139
timestamp 1624635492
transform 1 0 13892 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_172
timestamp 1624635492
transform 1 0 16928 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_163
timestamp 1624635492
transform 1 0 16100 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1624635492
transform 1 0 16836 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_196
timestamp 1624635492
transform 1 0 19136 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_184
timestamp 1624635492
transform 1 0 18032 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_208
timestamp 1624635492
transform 1 0 20240 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_229
timestamp 1624635492
transform 1 0 22172 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_220
timestamp 1624635492
transform 1 0 21344 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1624635492
transform 1 0 22080 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_253
timestamp 1624635492
transform 1 0 24380 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_241
timestamp 1624635492
transform 1 0 23276 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_265
timestamp 1624635492
transform 1 0 25484 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_156
timestamp 1624635492
transform 1 0 15456 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_144
timestamp 1624635492
transform 1 0 14352 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1624635492
transform 1 0 14260 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_168
timestamp 1624635492
transform 1 0 16560 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_192
timestamp 1624635492
transform 1 0 18768 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_180
timestamp 1624635492
transform 1 0 17664 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_213
timestamp 1624635492
transform 1 0 20700 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_201
timestamp 1624635492
transform 1 0 19596 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1624635492
transform 1 0 19504 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_225
timestamp 1624635492
transform 1 0 21804 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_249
timestamp 1624635492
transform 1 0 24012 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_237
timestamp 1624635492
transform 1 0 22908 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_270
timestamp 1624635492
transform 1 0 25944 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_258
timestamp 1624635492
transform 1 0 24840 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1624635492
transform 1 0 24748 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_156
timestamp 1624635492
transform 1 0 15456 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_144
timestamp 1624635492
transform 1 0 14352 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_151
timestamp 1624635492
transform 1 0 14996 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_139
timestamp 1624635492
transform 1 0 13892 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1624635492
transform 1 0 14260 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_168
timestamp 1624635492
transform 1 0 16560 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_172
timestamp 1624635492
transform 1 0 16928 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_163
timestamp 1624635492
transform 1 0 16100 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1624635492
transform 1 0 16836 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_192
timestamp 1624635492
transform 1 0 18768 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_180
timestamp 1624635492
transform 1 0 17664 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_196
timestamp 1624635492
transform 1 0 19136 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_184
timestamp 1624635492
transform 1 0 18032 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_213
timestamp 1624635492
transform 1 0 20700 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_201
timestamp 1624635492
transform 1 0 19596 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_208
timestamp 1624635492
transform 1 0 20240 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1624635492
transform 1 0 19504 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_225
timestamp 1624635492
transform 1 0 21804 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_229
timestamp 1624635492
transform 1 0 22172 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_220
timestamp 1624635492
transform 1 0 21344 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1624635492
transform 1 0 22080 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_249
timestamp 1624635492
transform 1 0 24012 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_237
timestamp 1624635492
transform 1 0 22908 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_253
timestamp 1624635492
transform 1 0 24380 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_241
timestamp 1624635492
transform 1 0 23276 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_270
timestamp 1624635492
transform 1 0 25944 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_258
timestamp 1624635492
transform 1 0 24840 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_265
timestamp 1624635492
transform 1 0 25484 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1624635492
transform 1 0 24748 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_151
timestamp 1624635492
transform 1 0 14996 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_139
timestamp 1624635492
transform 1 0 13892 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_172
timestamp 1624635492
transform 1 0 16928 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_163
timestamp 1624635492
transform 1 0 16100 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1624635492
transform 1 0 16836 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_196
timestamp 1624635492
transform 1 0 19136 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_184
timestamp 1624635492
transform 1 0 18032 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_208
timestamp 1624635492
transform 1 0 20240 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_229
timestamp 1624635492
transform 1 0 22172 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_220
timestamp 1624635492
transform 1 0 21344 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1624635492
transform 1 0 22080 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_253
timestamp 1624635492
transform 1 0 24380 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_241
timestamp 1624635492
transform 1 0 23276 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_265
timestamp 1624635492
transform 1 0 25484 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_156
timestamp 1624635492
transform 1 0 15456 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_144
timestamp 1624635492
transform 1 0 14352 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1624635492
transform 1 0 14260 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_168
timestamp 1624635492
transform 1 0 16560 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_192
timestamp 1624635492
transform 1 0 18768 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_180
timestamp 1624635492
transform 1 0 17664 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_213
timestamp 1624635492
transform 1 0 20700 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_201
timestamp 1624635492
transform 1 0 19596 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1624635492
transform 1 0 19504 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_225
timestamp 1624635492
transform 1 0 21804 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_249
timestamp 1624635492
transform 1 0 24012 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_237
timestamp 1624635492
transform 1 0 22908 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_270
timestamp 1624635492
transform 1 0 25944 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_258
timestamp 1624635492
transform 1 0 24840 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1624635492
transform 1 0 24748 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_151
timestamp 1624635492
transform 1 0 14996 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_139
timestamp 1624635492
transform 1 0 13892 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_172
timestamp 1624635492
transform 1 0 16928 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_163
timestamp 1624635492
transform 1 0 16100 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1249
timestamp 1624635492
transform 1 0 16836 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_187
timestamp 1624635492
transform 1 0 18308 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _230_
timestamp 1624635492
transform 1 0 18032 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_211
timestamp 1624635492
transform 1 0 20516 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_199
timestamp 1624635492
transform 1 0 19412 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_229
timestamp 1624635492
transform 1 0 22172 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_227
timestamp 1624635492
transform 1 0 21988 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_223
timestamp 1624635492
transform 1 0 21620 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1250
timestamp 1624635492
transform 1 0 22080 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_253
timestamp 1624635492
transform 1 0 24380 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_241
timestamp 1624635492
transform 1 0 23276 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_265
timestamp 1624635492
transform 1 0 25484 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_156
timestamp 1624635492
transform 1 0 15456 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_144
timestamp 1624635492
transform 1 0 14352 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_142
timestamp 1624635492
transform 1 0 14168 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1261
timestamp 1624635492
transform 1 0 14260 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_168
timestamp 1624635492
transform 1 0 16560 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_192
timestamp 1624635492
transform 1 0 18768 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_180
timestamp 1624635492
transform 1 0 17664 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_213
timestamp 1624635492
transform 1 0 20700 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_201
timestamp 1624635492
transform 1 0 19596 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1262
timestamp 1624635492
transform 1 0 19504 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_225
timestamp 1624635492
transform 1 0 21804 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_249
timestamp 1624635492
transform 1 0 24012 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_237
timestamp 1624635492
transform 1 0 22908 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_270
timestamp 1624635492
transform 1 0 25944 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_258
timestamp 1624635492
transform 1 0 24840 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1263
timestamp 1624635492
transform 1 0 24748 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_151
timestamp 1624635492
transform 1 0 14996 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_139
timestamp 1624635492
transform 1 0 13892 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_172
timestamp 1624635492
transform 1 0 16928 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_163
timestamp 1624635492
transform 1 0 16100 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1274
timestamp 1624635492
transform 1 0 16836 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _124_
timestamp 1624635492
transform -1 0 17572 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_191
timestamp 1624635492
transform 1 0 18676 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_179
timestamp 1624635492
transform 1 0 17572 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_215
timestamp 1624635492
transform 1 0 20884 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_203
timestamp 1624635492
transform 1 0 19780 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_229
timestamp 1624635492
transform 1 0 22172 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_227
timestamp 1624635492
transform 1 0 21988 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1275
timestamp 1624635492
transform 1 0 22080 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_253
timestamp 1624635492
transform 1 0 24380 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_241
timestamp 1624635492
transform 1 0 23276 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_268
timestamp 1624635492
transform 1 0 25760 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _128_
timestamp 1624635492
transform -1 0 25760 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_151
timestamp 1624635492
transform 1 0 14996 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_139
timestamp 1624635492
transform 1 0 13892 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_156
timestamp 1624635492
transform 1 0 15456 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_144
timestamp 1624635492
transform 1 0 14352 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1286
timestamp 1624635492
transform 1 0 14260 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_172
timestamp 1624635492
transform 1 0 16928 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_163
timestamp 1624635492
transform 1 0 16100 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_168
timestamp 1624635492
transform 1 0 16560 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1299
timestamp 1624635492
transform 1 0 16836 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_196
timestamp 1624635492
transform 1 0 19136 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_184
timestamp 1624635492
transform 1 0 18032 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_192
timestamp 1624635492
transform 1 0 18768 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_180
timestamp 1624635492
transform 1 0 17664 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_208
timestamp 1624635492
transform 1 0 20240 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_213
timestamp 1624635492
transform 1 0 20700 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_201
timestamp 1624635492
transform 1 0 19596 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1287
timestamp 1624635492
transform 1 0 19504 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_229
timestamp 1624635492
transform 1 0 22172 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_103_220
timestamp 1624635492
transform 1 0 21344 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_225
timestamp 1624635492
transform 1 0 21804 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1300
timestamp 1624635492
transform 1 0 22080 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _109_
timestamp 1624635492
transform 1 0 22540 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_255
timestamp 1624635492
transform 1 0 24564 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_243
timestamp 1624635492
transform 1 0 23460 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_236
timestamp 1624635492
transform 1 0 22816 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_102_249
timestamp 1624635492
transform 1 0 24012 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_237
timestamp 1624635492
transform 1 0 22908 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _126_
timestamp 1624635492
transform -1 0 23460 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_267
timestamp 1624635492
transform 1 0 25668 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_270
timestamp 1624635492
transform 1 0 25944 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_258
timestamp 1624635492
transform 1 0 24840 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1288
timestamp 1624635492
transform 1 0 24748 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_156
timestamp 1624635492
transform 1 0 15456 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_144
timestamp 1624635492
transform 1 0 14352 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_137
timestamp 1624635492
transform 1 0 13708 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1311
timestamp 1624635492
transform 1 0 14260 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_168
timestamp 1624635492
transform 1 0 16560 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_192
timestamp 1624635492
transform 1 0 18768 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_180
timestamp 1624635492
transform 1 0 17664 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_213
timestamp 1624635492
transform 1 0 20700 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_201
timestamp 1624635492
transform 1 0 19596 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1312
timestamp 1624635492
transform 1 0 19504 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_225
timestamp 1624635492
transform 1 0 21804 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_249
timestamp 1624635492
transform 1 0 24012 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_237
timestamp 1624635492
transform 1 0 22908 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_270
timestamp 1624635492
transform 1 0 25944 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_258
timestamp 1624635492
transform 1 0 24840 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1313
timestamp 1624635492
transform 1 0 24748 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_147
timestamp 1624635492
transform 1 0 14628 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_139
timestamp 1624635492
transform 1 0 13892 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _338_
timestamp 1624635492
transform -1 0 16468 0 1 59296
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_105_174
timestamp 1624635492
transform 1 0 17112 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_167
timestamp 1624635492
transform 1 0 16468 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__D
timestamp 1624635492
transform 1 0 16928 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1324
timestamp 1624635492
transform 1 0 16836 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_192
timestamp 1624635492
transform 1 0 18768 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_180
timestamp 1624635492
transform 1 0 17664 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__CLK
timestamp 1624635492
transform 1 0 17480 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_204
timestamp 1624635492
transform 1 0 19872 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_229
timestamp 1624635492
transform 1 0 22172 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_216
timestamp 1624635492
transform 1 0 20976 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1325
timestamp 1624635492
transform 1 0 22080 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_253
timestamp 1624635492
transform 1 0 24380 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_241
timestamp 1624635492
transform 1 0 23276 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_265
timestamp 1624635492
transform 1 0 25484 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_156
timestamp 1624635492
transform 1 0 15456 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_144
timestamp 1624635492
transform 1 0 14352 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1336
timestamp 1624635492
transform 1 0 14260 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_173
timestamp 1624635492
transform 1 0 17020 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_161
timestamp 1624635492
transform 1 0 15916 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _103_
timestamp 1624635492
transform 1 0 15640 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_185
timestamp 1624635492
transform 1 0 18124 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_213
timestamp 1624635492
transform 1 0 20700 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_201
timestamp 1624635492
transform 1 0 19596 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_197
timestamp 1624635492
transform 1 0 19228 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1337
timestamp 1624635492
transform 1 0 19504 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_225
timestamp 1624635492
transform 1 0 21804 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_249
timestamp 1624635492
transform 1 0 24012 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_237
timestamp 1624635492
transform 1 0 22908 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_270
timestamp 1624635492
transform 1 0 25944 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_258
timestamp 1624635492
transform 1 0 24840 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1338
timestamp 1624635492
transform 1 0 24748 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_282
timestamp 1624635492
transform 1 0 27048 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_294
timestamp 1624635492
transform 1 0 28152 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_306
timestamp 1624635492
transform 1 0 29256 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_315
timestamp 1624635492
transform 1 0 30084 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1624635492
transform 1 0 29992 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_327
timestamp 1624635492
transform 1 0 31188 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_339
timestamp 1624635492
transform 1 0 32292 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_363
timestamp 1624635492
transform 1 0 34500 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_351
timestamp 1624635492
transform 1 0 33396 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_372
timestamp 1624635492
transform 1 0 35328 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1624635492
transform 1 0 35236 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_384
timestamp 1624635492
transform 1 0 36432 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_396
timestamp 1624635492
transform 1 0 37536 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_408
timestamp 1624635492
transform 1 0 38640 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_277
timestamp 1624635492
transform 1 0 26588 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1624635492
transform 1 0 27324 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_298
timestamp 1624635492
transform 1 0 28520 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_286
timestamp 1624635492
transform 1 0 27416 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_310
timestamp 1624635492
transform 1 0 29624 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_322
timestamp 1624635492
transform 1 0 30728 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_334
timestamp 1624635492
transform 1 0 31832 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_343
timestamp 1624635492
transform 1 0 32660 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1624635492
transform 1 0 32568 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_355
timestamp 1624635492
transform 1 0 33764 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_367
timestamp 1624635492
transform 1 0 34868 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_379
timestamp 1624635492
transform 1 0 35972 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_400
timestamp 1624635492
transform 1 0 37904 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_391
timestamp 1624635492
transform 1 0 37076 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1624635492
transform 1 0 37812 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_277
timestamp 1624635492
transform 1 0 26588 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_284
timestamp 1624635492
transform 1 0 27232 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1624635492
transform 1 0 27324 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_298
timestamp 1624635492
transform 1 0 28520 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_286
timestamp 1624635492
transform 1 0 27416 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_296
timestamp 1624635492
transform 1 0 28336 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_310
timestamp 1624635492
transform 1 0 29624 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_308
timestamp 1624635492
transform 1 0 29440 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_322
timestamp 1624635492
transform 1 0 30728 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_315
timestamp 1624635492
transform 1 0 30084 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1624635492
transform 1 0 29992 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_334
timestamp 1624635492
transform 1 0 31832 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_335
timestamp 1624635492
transform 1 0 31924 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_327
timestamp 1624635492
transform 1 0 31188 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1624635492
transform 1 0 31740 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_343
timestamp 1624635492
transform 1 0 32660 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_346
timestamp 1624635492
transform 1 0 32936 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1624635492
transform 1 0 32568 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _061_
timestamp 1624635492
transform -1 0 32936 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_83_355
timestamp 1624635492
transform 1 0 33764 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_358
timestamp 1624635492
transform 1 0 34040 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_367
timestamp 1624635492
transform 1 0 34868 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_372
timestamp 1624635492
transform 1 0 35328 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_370
timestamp 1624635492
transform 1 0 35144 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1624635492
transform 1 0 35236 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_379
timestamp 1624635492
transform 1 0 35972 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_384
timestamp 1624635492
transform 1 0 36432 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_400
timestamp 1624635492
transform 1 0 37904 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_391
timestamp 1624635492
transform 1 0 37076 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_396
timestamp 1624635492
transform 1 0 37536 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1624635492
transform 1 0 37812 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_408
timestamp 1624635492
transform 1 0 38640 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_282
timestamp 1624635492
transform 1 0 27048 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_294
timestamp 1624635492
transform 1 0 28152 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_306
timestamp 1624635492
transform 1 0 29256 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_315
timestamp 1624635492
transform 1 0 30084 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1624635492
transform 1 0 29992 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_327
timestamp 1624635492
transform 1 0 31188 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_339
timestamp 1624635492
transform 1 0 32292 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_363
timestamp 1624635492
transform 1 0 34500 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_351
timestamp 1624635492
transform 1 0 33396 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_372
timestamp 1624635492
transform 1 0 35328 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1624635492
transform 1 0 35236 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_384
timestamp 1624635492
transform 1 0 36432 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_396
timestamp 1624635492
transform 1 0 37536 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_408
timestamp 1624635492
transform 1 0 38640 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_277
timestamp 1624635492
transform 1 0 26588 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1624635492
transform 1 0 27324 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_298
timestamp 1624635492
transform 1 0 28520 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_286
timestamp 1624635492
transform 1 0 27416 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_310
timestamp 1624635492
transform 1 0 29624 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_322
timestamp 1624635492
transform 1 0 30728 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_334
timestamp 1624635492
transform 1 0 31832 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_343
timestamp 1624635492
transform 1 0 32660 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1624635492
transform 1 0 32568 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_355
timestamp 1624635492
transform 1 0 33764 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_367
timestamp 1624635492
transform 1 0 34868 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_379
timestamp 1624635492
transform 1 0 35972 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_400
timestamp 1624635492
transform 1 0 37904 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_391
timestamp 1624635492
transform 1 0 37076 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1624635492
transform 1 0 37812 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_282
timestamp 1624635492
transform 1 0 27048 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_294
timestamp 1624635492
transform 1 0 28152 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_306
timestamp 1624635492
transform 1 0 29256 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_315
timestamp 1624635492
transform 1 0 30084 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1624635492
transform 1 0 29992 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_327
timestamp 1624635492
transform 1 0 31188 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_339
timestamp 1624635492
transform 1 0 32292 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_359
timestamp 1624635492
transform 1 0 34132 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_351
timestamp 1624635492
transform 1 0 33396 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B1
timestamp 1624635492
transform 1 0 33948 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_372
timestamp 1624635492
transform 1 0 35328 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1624635492
transform 1 0 35236 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_384
timestamp 1624635492
transform 1 0 36432 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_396
timestamp 1624635492
transform 1 0 37536 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_408
timestamp 1624635492
transform 1 0 38640 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_277
timestamp 1624635492
transform 1 0 26588 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1624635492
transform 1 0 27324 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_298
timestamp 1624635492
transform 1 0 28520 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_286
timestamp 1624635492
transform 1 0 27416 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_310
timestamp 1624635492
transform 1 0 29624 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_322
timestamp 1624635492
transform 1 0 30728 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_334
timestamp 1624635492
transform 1 0 31832 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_343
timestamp 1624635492
transform 1 0 32660 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1624635492
transform 1 0 32568 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_357
timestamp 1624635492
transform 1 0 33948 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A1
timestamp 1624635492
transform 1 0 33764 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _098_
timestamp 1624635492
transform 1 0 34316 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_87_375
timestamp 1624635492
transform 1 0 35604 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_369
timestamp 1624635492
transform 1 0 35052 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B2
timestamp 1624635492
transform 1 0 35420 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_381
timestamp 1624635492
transform 1 0 36156 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A2
timestamp 1624635492
transform -1 0 36156 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_400
timestamp 1624635492
transform 1 0 37904 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_393
timestamp 1624635492
transform 1 0 37260 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1624635492
transform 1 0 37812 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_277
timestamp 1624635492
transform 1 0 26588 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_282
timestamp 1624635492
transform 1 0 27048 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1624635492
transform 1 0 27324 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_298
timestamp 1624635492
transform 1 0 28520 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_286
timestamp 1624635492
transform 1 0 27416 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_294
timestamp 1624635492
transform 1 0 28152 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_310
timestamp 1624635492
transform 1 0 29624 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_306
timestamp 1624635492
transform 1 0 29256 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_322
timestamp 1624635492
transform 1 0 30728 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_315
timestamp 1624635492
transform 1 0 30084 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1624635492
transform 1 0 29992 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_334
timestamp 1624635492
transform 1 0 31832 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_327
timestamp 1624635492
transform 1 0 31188 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_343
timestamp 1624635492
transform 1 0 32660 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_339
timestamp 1624635492
transform 1 0 32292 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1624635492
transform 1 0 32568 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_361
timestamp 1624635492
transform 1 0 34316 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_355
timestamp 1624635492
transform 1 0 33764 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_88_359
timestamp 1624635492
transform 1 0 34132 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_88_351
timestamp 1624635492
transform 1 0 33396 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _324_
timestamp 1624635492
transform -1 0 34684 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _123_
timestamp 1624635492
transform -1 0 34684 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_365
timestamp 1624635492
transform 1 0 34684 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_372
timestamp 1624635492
transform 1 0 35328 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_365
timestamp 1624635492
transform 1 0 34684 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1624635492
transform 1 0 35236 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_377
timestamp 1624635492
transform 1 0 35788 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_384
timestamp 1624635492
transform 1 0 36432 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_400
timestamp 1624635492
transform 1 0 37904 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_397
timestamp 1624635492
transform 1 0 37628 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_389
timestamp 1624635492
transform 1 0 36892 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_396
timestamp 1624635492
transform 1 0 37536 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1624635492
transform 1 0 37812 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_408
timestamp 1624635492
transform 1 0 38640 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_282
timestamp 1624635492
transform 1 0 27048 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_294
timestamp 1624635492
transform 1 0 28152 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_306
timestamp 1624635492
transform 1 0 29256 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_315
timestamp 1624635492
transform 1 0 30084 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1624635492
transform 1 0 29992 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_331
timestamp 1624635492
transform 1 0 31556 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_327
timestamp 1624635492
transform 1 0 31188 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _142_
timestamp 1624635492
transform 1 0 31280 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_343
timestamp 1624635492
transform 1 0 32660 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_355
timestamp 1624635492
transform 1 0 33764 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_372
timestamp 1624635492
transform 1 0 35328 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_367
timestamp 1624635492
transform 1 0 34868 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1624635492
transform 1 0 35236 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_384
timestamp 1624635492
transform 1 0 36432 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_396
timestamp 1624635492
transform 1 0 37536 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_408
timestamp 1624635492
transform 1 0 38640 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_277
timestamp 1624635492
transform 1 0 26588 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1624635492
transform 1 0 27324 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_298
timestamp 1624635492
transform 1 0 28520 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_286
timestamp 1624635492
transform 1 0 27416 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_310
timestamp 1624635492
transform 1 0 29624 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_322
timestamp 1624635492
transform 1 0 30728 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_334
timestamp 1624635492
transform 1 0 31832 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_343
timestamp 1624635492
transform 1 0 32660 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1624635492
transform 1 0 32568 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_355
timestamp 1624635492
transform 1 0 33764 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_367
timestamp 1624635492
transform 1 0 34868 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_379
timestamp 1624635492
transform 1 0 35972 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_400
timestamp 1624635492
transform 1 0 37904 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_391
timestamp 1624635492
transform 1 0 37076 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1624635492
transform 1 0 37812 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_283
timestamp 1624635492
transform 1 0 27140 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_278
timestamp 1624635492
transform 1 0 26680 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _296_
timestamp 1624635492
transform 1 0 26864 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_295
timestamp 1624635492
transform 1 0 28244 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_307
timestamp 1624635492
transform 1 0 29348 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_92_315
timestamp 1624635492
transform 1 0 30084 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_313
timestamp 1624635492
transform 1 0 29900 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1624635492
transform 1 0 29992 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_327
timestamp 1624635492
transform 1 0 31188 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_339
timestamp 1624635492
transform 1 0 32292 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_363
timestamp 1624635492
transform 1 0 34500 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_351
timestamp 1624635492
transform 1 0 33396 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_372
timestamp 1624635492
transform 1 0 35328 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1624635492
transform 1 0 35236 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_384
timestamp 1624635492
transform 1 0 36432 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_396
timestamp 1624635492
transform 1 0 37536 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_408
timestamp 1624635492
transform 1 0 38640 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_277
timestamp 1624635492
transform 1 0 26588 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1624635492
transform 1 0 27324 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_298
timestamp 1624635492
transform 1 0 28520 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_286
timestamp 1624635492
transform 1 0 27416 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_310
timestamp 1624635492
transform 1 0 29624 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_322
timestamp 1624635492
transform 1 0 30728 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_334
timestamp 1624635492
transform 1 0 31832 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B1
timestamp 1624635492
transform 1 0 32016 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_345
timestamp 1624635492
transform 1 0 32844 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_338
timestamp 1624635492
transform 1 0 32200 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A3
timestamp 1624635492
transform 1 0 32660 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1624635492
transform 1 0 32568 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_357
timestamp 1624635492
transform 1 0 33948 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_369
timestamp 1624635492
transform 1 0 35052 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_381
timestamp 1624635492
transform 1 0 36156 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_400
timestamp 1624635492
transform 1 0 37904 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_393
timestamp 1624635492
transform 1 0 37260 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1624635492
transform 1 0 37812 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_282
timestamp 1624635492
transform 1 0 27048 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_94_294
timestamp 1624635492
transform 1 0 28152 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_290
timestamp 1624635492
transform 1 0 27784 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1624635492
transform 1 0 27968 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  _072_
timestamp 1624635492
transform 1 0 28520 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_310
timestamp 1624635492
transform 1 0 29624 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_315
timestamp 1624635492
transform 1 0 30084 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1624635492
transform 1 0 29992 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_334
timestamp 1624635492
transform 1 0 31832 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_331
timestamp 1624635492
transform 1 0 31556 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_327
timestamp 1624635492
transform 1 0 31188 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A2
timestamp 1624635492
transform 1 0 31648 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_340
timestamp 1624635492
transform 1 0 32384 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A1
timestamp 1624635492
transform 1 0 32200 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 33396 0 -1 53856
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_94_363
timestamp 1624635492
transform 1 0 34500 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_351
timestamp 1624635492
transform 1 0 33396 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_372
timestamp 1624635492
transform 1 0 35328 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1624635492
transform 1 0 35236 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_384
timestamp 1624635492
transform 1 0 36432 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_396
timestamp 1624635492
transform 1 0 37536 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_408
timestamp 1624635492
transform 1 0 38640 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_282
timestamp 1624635492
transform 1 0 27048 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_277
timestamp 1624635492
transform 1 0 26588 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1624635492
transform 1 0 27324 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_294
timestamp 1624635492
transform 1 0 28152 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_298
timestamp 1624635492
transform 1 0 28520 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_286
timestamp 1624635492
transform 1 0 27416 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_306
timestamp 1624635492
transform 1 0 29256 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_310
timestamp 1624635492
transform 1 0 29624 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_315
timestamp 1624635492
transform 1 0 30084 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_322
timestamp 1624635492
transform 1 0 30728 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1624635492
transform 1 0 29992 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_327
timestamp 1624635492
transform 1 0 31188 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_334
timestamp 1624635492
transform 1 0 31832 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_339
timestamp 1624635492
transform 1 0 32292 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_343
timestamp 1624635492
transform 1 0 32660 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1624635492
transform 1 0 32568 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_363
timestamp 1624635492
transform 1 0 34500 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_351
timestamp 1624635492
transform 1 0 33396 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_355
timestamp 1624635492
transform 1 0 33764 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_372
timestamp 1624635492
transform 1 0 35328 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_367
timestamp 1624635492
transform 1 0 34868 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1624635492
transform 1 0 35236 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_384
timestamp 1624635492
transform 1 0 36432 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_379
timestamp 1624635492
transform 1 0 35972 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_396
timestamp 1624635492
transform 1 0 37536 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_400
timestamp 1624635492
transform 1 0 37904 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_391
timestamp 1624635492
transform 1 0 37076 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1624635492
transform 1 0 37812 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_404
timestamp 1624635492
transform 1 0 38272 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A2
timestamp 1624635492
transform 1 0 38088 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_277
timestamp 1624635492
transform 1 0 26588 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1624635492
transform 1 0 27324 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_298
timestamp 1624635492
transform 1 0 28520 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_286
timestamp 1624635492
transform 1 0 27416 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_310
timestamp 1624635492
transform 1 0 29624 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_322
timestamp 1624635492
transform 1 0 30728 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_334
timestamp 1624635492
transform 1 0 31832 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_343
timestamp 1624635492
transform 1 0 32660 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1624635492
transform 1 0 32568 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_355
timestamp 1624635492
transform 1 0 33764 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_367
timestamp 1624635492
transform 1 0 34868 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_379
timestamp 1624635492
transform 1 0 35972 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_400
timestamp 1624635492
transform 1 0 37904 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_395
timestamp 1624635492
transform 1 0 37444 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_391
timestamp 1624635492
transform 1 0 37076 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A3
timestamp 1624635492
transform 1 0 37260 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1624635492
transform 1 0 37812 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_2  _090_
timestamp 1624635492
transform 1 0 38272 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_98_282
timestamp 1624635492
transform 1 0 27048 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_294
timestamp 1624635492
transform 1 0 28152 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_306
timestamp 1624635492
transform 1 0 29256 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_315
timestamp 1624635492
transform 1 0 30084 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1624635492
transform 1 0 29992 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_327
timestamp 1624635492
transform 1 0 31188 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_339
timestamp 1624635492
transform 1 0 32292 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_363
timestamp 1624635492
transform 1 0 34500 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_351
timestamp 1624635492
transform 1 0 33396 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_372
timestamp 1624635492
transform 1 0 35328 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1624635492
transform 1 0 35236 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_384
timestamp 1624635492
transform 1 0 36432 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_396
timestamp 1624635492
transform 1 0 37536 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A1
timestamp 1624635492
transform -1 0 38088 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_98_402
timestamp 1624635492
transform 1 0 38088 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_277
timestamp 1624635492
transform 1 0 26588 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1251
timestamp 1624635492
transform 1 0 27324 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_298
timestamp 1624635492
transform 1 0 28520 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_286
timestamp 1624635492
transform 1 0 27416 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_310
timestamp 1624635492
transform 1 0 29624 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_320
timestamp 1624635492
transform 1 0 30544 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_316
timestamp 1624635492
transform 1 0 30176 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _323_
timestamp 1624635492
transform -1 0 30544 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_332
timestamp 1624635492
transform 1 0 31648 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_343
timestamp 1624635492
transform 1 0 32660 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_340
timestamp 1624635492
transform 1 0 32384 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1252
timestamp 1624635492
transform 1 0 32568 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_355
timestamp 1624635492
transform 1 0 33764 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_367
timestamp 1624635492
transform 1 0 34868 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_379
timestamp 1624635492
transform 1 0 35972 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_400
timestamp 1624635492
transform 1 0 37904 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_391
timestamp 1624635492
transform 1 0 37076 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1253
timestamp 1624635492
transform 1 0 37812 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_282
timestamp 1624635492
transform 1 0 27048 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_294
timestamp 1624635492
transform 1 0 28152 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_306
timestamp 1624635492
transform 1 0 29256 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_315
timestamp 1624635492
transform 1 0 30084 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1264
timestamp 1624635492
transform 1 0 29992 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_327
timestamp 1624635492
transform 1 0 31188 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_339
timestamp 1624635492
transform 1 0 32292 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_363
timestamp 1624635492
transform 1 0 34500 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_351
timestamp 1624635492
transform 1 0 33396 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_372
timestamp 1624635492
transform 1 0 35328 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1265
timestamp 1624635492
transform 1 0 35236 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_384
timestamp 1624635492
transform 1 0 36432 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_396
timestamp 1624635492
transform 1 0 37536 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_408
timestamp 1624635492
transform 1 0 38640 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_284
timestamp 1624635492
transform 1 0 27232 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_280
timestamp 1624635492
transform 1 0 26864 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1276
timestamp 1624635492
transform 1 0 27324 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_298
timestamp 1624635492
transform 1 0 28520 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_286
timestamp 1624635492
transform 1 0 27416 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_310
timestamp 1624635492
transform 1 0 29624 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_322
timestamp 1624635492
transform 1 0 30728 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_334
timestamp 1624635492
transform 1 0 31832 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_343
timestamp 1624635492
transform 1 0 32660 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1277
timestamp 1624635492
transform 1 0 32568 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_355
timestamp 1624635492
transform 1 0 33764 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_367
timestamp 1624635492
transform 1 0 34868 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _315_
timestamp 1624635492
transform -1 0 35880 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_378
timestamp 1624635492
transform 1 0 35880 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_400
timestamp 1624635492
transform 1 0 37904 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_398
timestamp 1624635492
transform 1 0 37720 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_390
timestamp 1624635492
transform 1 0 36984 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1278
timestamp 1624635492
transform 1 0 37812 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_103_279
timestamp 1624635492
transform 1 0 26772 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_102_282
timestamp 1624635492
transform 1 0 27048 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1301
timestamp 1624635492
transform 1 0 27324 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_293
timestamp 1624635492
transform 1 0 28060 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_286
timestamp 1624635492
transform 1 0 27416 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_296
timestamp 1624635492
transform 1 0 28336 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_102_290
timestamp 1624635492
transform 1 0 27784 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _238_
timestamp 1624635492
transform 1 0 27784 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _122_
timestamp 1624635492
transform -1 0 28336 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_305
timestamp 1624635492
transform 1 0 29164 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_308
timestamp 1624635492
transform 1 0 29440 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_103_317
timestamp 1624635492
transform 1 0 30268 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_315
timestamp 1624635492
transform 1 0 30084 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1289
timestamp 1624635492
transform 1 0 29992 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_329
timestamp 1624635492
transform 1 0 31372 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_327
timestamp 1624635492
transform 1 0 31188 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_343
timestamp 1624635492
transform 1 0 32660 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_341
timestamp 1624635492
transform 1 0 32476 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_339
timestamp 1624635492
transform 1 0 32292 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1302
timestamp 1624635492
transform 1 0 32568 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_103_355
timestamp 1624635492
transform 1 0 33764 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_102_363
timestamp 1624635492
transform 1 0 34500 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_351
timestamp 1624635492
transform 1 0 33396 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _235_
timestamp 1624635492
transform 1 0 34316 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_364
timestamp 1624635492
transform 1 0 34592 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_372
timestamp 1624635492
transform 1 0 35328 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1290
timestamp 1624635492
transform 1 0 35236 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_388
timestamp 1624635492
transform 1 0 36800 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_376
timestamp 1624635492
transform 1 0 35696 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_382
timestamp 1624635492
transform 1 0 36248 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_378
timestamp 1624635492
transform 1 0 35880 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _242_
timestamp 1624635492
transform 1 0 35972 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_400
timestamp 1624635492
transform 1 0 37904 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_396
timestamp 1624635492
transform 1 0 37536 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_394
timestamp 1624635492
transform 1 0 37352 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1303
timestamp 1624635492
transform 1 0 37812 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_406
timestamp 1624635492
transform 1 0 38456 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_282
timestamp 1624635492
transform 1 0 27048 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_294
timestamp 1624635492
transform 1 0 28152 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_306
timestamp 1624635492
transform 1 0 29256 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_315
timestamp 1624635492
transform 1 0 30084 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1314
timestamp 1624635492
transform 1 0 29992 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_327
timestamp 1624635492
transform 1 0 31188 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_339
timestamp 1624635492
transform 1 0 32292 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_363
timestamp 1624635492
transform 1 0 34500 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_351
timestamp 1624635492
transform 1 0 33396 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_372
timestamp 1624635492
transform 1 0 35328 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1315
timestamp 1624635492
transform 1 0 35236 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_384
timestamp 1624635492
transform 1 0 36432 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_396
timestamp 1624635492
transform 1 0 37536 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_408
timestamp 1624635492
transform 1 0 38640 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_277
timestamp 1624635492
transform 1 0 26588 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1326
timestamp 1624635492
transform 1 0 27324 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_298
timestamp 1624635492
transform 1 0 28520 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_286
timestamp 1624635492
transform 1 0 27416 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_310
timestamp 1624635492
transform 1 0 29624 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_322
timestamp 1624635492
transform 1 0 30728 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_334
timestamp 1624635492
transform 1 0 31832 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_343
timestamp 1624635492
transform 1 0 32660 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1327
timestamp 1624635492
transform 1 0 32568 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_355
timestamp 1624635492
transform 1 0 33764 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_367
timestamp 1624635492
transform 1 0 34868 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_379
timestamp 1624635492
transform 1 0 35972 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_400
timestamp 1624635492
transform 1 0 37904 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_391
timestamp 1624635492
transform 1 0 37076 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1328
timestamp 1624635492
transform 1 0 37812 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_282
timestamp 1624635492
transform 1 0 27048 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_294
timestamp 1624635492
transform 1 0 28152 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_306
timestamp 1624635492
transform 1 0 29256 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_315
timestamp 1624635492
transform 1 0 30084 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1339
timestamp 1624635492
transform 1 0 29992 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_327
timestamp 1624635492
transform 1 0 31188 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_339
timestamp 1624635492
transform 1 0 32292 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_363
timestamp 1624635492
transform 1 0 34500 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_351
timestamp 1624635492
transform 1 0 33396 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_372
timestamp 1624635492
transform 1 0 35328 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1340
timestamp 1624635492
transform 1 0 35236 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_384
timestamp 1624635492
transform 1 0 36432 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_396
timestamp 1624635492
transform 1 0 37536 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_408
timestamp 1624635492
transform 1 0 38640 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_417
timestamp 1624635492
transform 1 0 39468 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_414
timestamp 1624635492
transform 1 0 39192 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A1
timestamp 1624635492
transform 1 0 39284 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_429
timestamp 1624635492
transform 1 0 40572 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_425
timestamp 1624635492
transform 1 0 40204 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1624635492
transform 1 0 40480 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_441
timestamp 1624635492
transform 1 0 41676 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_453
timestamp 1624635492
transform 1 0 42780 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_465
timestamp 1624635492
transform 1 0 43884 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_486
timestamp 1624635492
transform 1 0 45816 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_477
timestamp 1624635492
transform 1 0 44988 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1624635492
transform 1 0 45724 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_498
timestamp 1624635492
transform 1 0 46920 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_510
timestamp 1624635492
transform 1 0 48024 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_522
timestamp 1624635492
transform 1 0 49128 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_534
timestamp 1624635492
transform 1 0 50232 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_543
timestamp 1624635492
transform 1 0 51060 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1624635492
transform 1 0 50968 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_412
timestamp 1624635492
transform 1 0 39008 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_424
timestamp 1624635492
transform 1 0 40112 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_448
timestamp 1624635492
transform 1 0 42320 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_436
timestamp 1624635492
transform 1 0 41216 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_457
timestamp 1624635492
transform 1 0 43148 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1624635492
transform 1 0 43056 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_469
timestamp 1624635492
transform 1 0 44252 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_481
timestamp 1624635492
transform 1 0 45356 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_493
timestamp 1624635492
transform 1 0 46460 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1624635492
transform 1 0 47564 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_514
timestamp 1624635492
transform 1 0 48392 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1624635492
transform 1 0 48300 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_538
timestamp 1624635492
transform 1 0 50600 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_526
timestamp 1624635492
transform 1 0 49496 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_412
timestamp 1624635492
transform 1 0 39008 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_420
timestamp 1624635492
transform 1 0 39744 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_416
timestamp 1624635492
transform 1 0 39376 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _228_
timestamp 1624635492
transform 1 0 39468 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_424
timestamp 1624635492
transform 1 0 40112 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1624635492
transform 1 0 40572 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1624635492
transform 1 0 40480 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_448
timestamp 1624635492
transform 1 0 42320 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_436
timestamp 1624635492
transform 1 0 41216 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_441
timestamp 1624635492
transform 1 0 41676 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_457
timestamp 1624635492
transform 1 0 43148 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_453
timestamp 1624635492
transform 1 0 42780 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1624635492
transform 1 0 43056 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_469
timestamp 1624635492
transform 1 0 44252 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_465
timestamp 1624635492
transform 1 0 43884 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_481
timestamp 1624635492
transform 1 0 45356 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_486
timestamp 1624635492
transform 1 0 45816 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_477
timestamp 1624635492
transform 1 0 44988 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1624635492
transform 1 0 45724 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_493
timestamp 1624635492
transform 1 0 46460 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_498
timestamp 1624635492
transform 1 0 46920 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_505
timestamp 1624635492
transform 1 0 47564 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_510
timestamp 1624635492
transform 1 0 48024 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_514
timestamp 1624635492
transform 1 0 48392 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_522
timestamp 1624635492
transform 1 0 49128 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1624635492
transform 1 0 48300 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_538
timestamp 1624635492
transform 1 0 50600 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_526
timestamp 1624635492
transform 1 0 49496 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_530
timestamp 1624635492
transform 1 0 49864 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_526
timestamp 1624635492
transform 1 0 49496 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _192_
timestamp 1624635492
transform -1 0 49864 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_543
timestamp 1624635492
transform 1 0 51060 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1624635492
transform 1 0 50968 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_420
timestamp 1624635492
transform 1 0 39744 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_429
timestamp 1624635492
transform 1 0 40572 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1624635492
transform 1 0 40480 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_441
timestamp 1624635492
transform 1 0 41676 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_453
timestamp 1624635492
transform 1 0 42780 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_465
timestamp 1624635492
transform 1 0 43884 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_486
timestamp 1624635492
transform 1 0 45816 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_484
timestamp 1624635492
transform 1 0 45632 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_480
timestamp 1624635492
transform 1 0 45264 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1624635492
transform 1 0 45724 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _177_
timestamp 1624635492
transform -1 0 45264 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_498
timestamp 1624635492
transform 1 0 46920 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_510
timestamp 1624635492
transform 1 0 48024 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_522
timestamp 1624635492
transform 1 0 49128 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_534
timestamp 1624635492
transform 1 0 50232 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_543
timestamp 1624635492
transform 1 0 51060 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1624635492
transform 1 0 50968 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_412
timestamp 1624635492
transform 1 0 39008 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_424
timestamp 1624635492
transform 1 0 40112 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_448
timestamp 1624635492
transform 1 0 42320 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_436
timestamp 1624635492
transform 1 0 41216 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_457
timestamp 1624635492
transform 1 0 43148 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1624635492
transform 1 0 43056 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_469
timestamp 1624635492
transform 1 0 44252 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_481
timestamp 1624635492
transform 1 0 45356 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_493
timestamp 1624635492
transform 1 0 46460 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_505
timestamp 1624635492
transform 1 0 47564 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_514
timestamp 1624635492
transform 1 0 48392 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1624635492
transform 1 0 48300 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_538
timestamp 1624635492
transform 1 0 50600 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_526
timestamp 1624635492
transform 1 0 49496 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_420
timestamp 1624635492
transform 1 0 39744 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_429
timestamp 1624635492
transform 1 0 40572 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1624635492
transform 1 0 40480 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_441
timestamp 1624635492
transform 1 0 41676 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_453
timestamp 1624635492
transform 1 0 42780 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_465
timestamp 1624635492
transform 1 0 43884 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_486
timestamp 1624635492
transform 1 0 45816 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_477
timestamp 1624635492
transform 1 0 44988 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1624635492
transform 1 0 45724 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_498
timestamp 1624635492
transform 1 0 46920 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_510
timestamp 1624635492
transform 1 0 48024 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_522
timestamp 1624635492
transform 1 0 49128 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_534
timestamp 1624635492
transform 1 0 50232 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_543
timestamp 1624635492
transform 1 0 51060 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1624635492
transform 1 0 50968 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_412
timestamp 1624635492
transform 1 0 39008 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_424
timestamp 1624635492
transform 1 0 40112 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_448
timestamp 1624635492
transform 1 0 42320 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_436
timestamp 1624635492
transform 1 0 41216 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_457
timestamp 1624635492
transform 1 0 43148 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1624635492
transform 1 0 43056 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_469
timestamp 1624635492
transform 1 0 44252 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_481
timestamp 1624635492
transform 1 0 45356 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_493
timestamp 1624635492
transform 1 0 46460 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_505
timestamp 1624635492
transform 1 0 47564 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_514
timestamp 1624635492
transform 1 0 48392 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1624635492
transform 1 0 48300 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_538
timestamp 1624635492
transform 1 0 50600 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_526
timestamp 1624635492
transform 1 0 49496 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_412
timestamp 1624635492
transform 1 0 39008 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_420
timestamp 1624635492
transform 1 0 39744 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_424
timestamp 1624635492
transform 1 0 40112 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_429
timestamp 1624635492
transform 1 0 40572 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1624635492
transform 1 0 40480 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_448
timestamp 1624635492
transform 1 0 42320 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_436
timestamp 1624635492
transform 1 0 41216 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_441
timestamp 1624635492
transform 1 0 41676 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_457
timestamp 1624635492
transform 1 0 43148 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_453
timestamp 1624635492
transform 1 0 42780 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1624635492
transform 1 0 43056 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_469
timestamp 1624635492
transform 1 0 44252 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_465
timestamp 1624635492
transform 1 0 43884 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_481
timestamp 1624635492
transform 1 0 45356 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_486
timestamp 1624635492
transform 1 0 45816 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_477
timestamp 1624635492
transform 1 0 44988 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1624635492
transform 1 0 45724 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_493
timestamp 1624635492
transform 1 0 46460 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_498
timestamp 1624635492
transform 1 0 46920 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_505
timestamp 1624635492
transform 1 0 47564 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_510
timestamp 1624635492
transform 1 0 48024 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_514
timestamp 1624635492
transform 1 0 48392 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_522
timestamp 1624635492
transform 1 0 49128 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1624635492
transform 1 0 48300 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_538
timestamp 1624635492
transform 1 0 50600 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_526
timestamp 1624635492
transform 1 0 49496 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_534
timestamp 1624635492
transform 1 0 50232 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_543
timestamp 1624635492
transform 1 0 51060 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1624635492
transform 1 0 50968 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_420
timestamp 1624635492
transform 1 0 39744 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_429
timestamp 1624635492
transform 1 0 40572 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1624635492
transform 1 0 40480 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_441
timestamp 1624635492
transform 1 0 41676 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_453
timestamp 1624635492
transform 1 0 42780 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_465
timestamp 1624635492
transform 1 0 43884 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_486
timestamp 1624635492
transform 1 0 45816 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_477
timestamp 1624635492
transform 1 0 44988 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1624635492
transform 1 0 45724 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_493
timestamp 1624635492
transform 1 0 46460 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _211_
timestamp 1624635492
transform -1 0 46460 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_505
timestamp 1624635492
transform 1 0 47564 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_517
timestamp 1624635492
transform 1 0 48668 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_529
timestamp 1624635492
transform 1 0 49772 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_543
timestamp 1624635492
transform 1 0 51060 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_541
timestamp 1624635492
transform 1 0 50876 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1624635492
transform 1 0 50968 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_412
timestamp 1624635492
transform 1 0 39008 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_424
timestamp 1624635492
transform 1 0 40112 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_448
timestamp 1624635492
transform 1 0 42320 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_436
timestamp 1624635492
transform 1 0 41216 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_457
timestamp 1624635492
transform 1 0 43148 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1624635492
transform 1 0 43056 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_469
timestamp 1624635492
transform 1 0 44252 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_481
timestamp 1624635492
transform 1 0 45356 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_493
timestamp 1624635492
transform 1 0 46460 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_505
timestamp 1624635492
transform 1 0 47564 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_514
timestamp 1624635492
transform 1 0 48392 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1624635492
transform 1 0 48300 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_538
timestamp 1624635492
transform 1 0 50600 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_526
timestamp 1624635492
transform 1 0 49496 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_420
timestamp 1624635492
transform 1 0 39744 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_429
timestamp 1624635492
transform 1 0 40572 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1624635492
transform 1 0 40480 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_441
timestamp 1624635492
transform 1 0 41676 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_453
timestamp 1624635492
transform 1 0 42780 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_465
timestamp 1624635492
transform 1 0 43884 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_486
timestamp 1624635492
transform 1 0 45816 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_477
timestamp 1624635492
transform 1 0 44988 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1624635492
transform 1 0 45724 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_498
timestamp 1624635492
transform 1 0 46920 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_510
timestamp 1624635492
transform 1 0 48024 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_522
timestamp 1624635492
transform 1 0 49128 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_534
timestamp 1624635492
transform 1 0 50232 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_543
timestamp 1624635492
transform 1 0 51060 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1624635492
transform 1 0 50968 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_412
timestamp 1624635492
transform 1 0 39008 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_431
timestamp 1624635492
transform 1 0 40756 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_424
timestamp 1624635492
transform 1 0 40112 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _232_
timestamp 1624635492
transform 1 0 41124 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _153_
timestamp 1624635492
transform 1 0 40480 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_438
timestamp 1624635492
transform 1 0 41400 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_457
timestamp 1624635492
transform 1 0 43148 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_450
timestamp 1624635492
transform 1 0 42504 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1624635492
transform 1 0 43056 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_469
timestamp 1624635492
transform 1 0 44252 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_481
timestamp 1624635492
transform 1 0 45356 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_493
timestamp 1624635492
transform 1 0 46460 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_505
timestamp 1624635492
transform 1 0 47564 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_514
timestamp 1624635492
transform 1 0 48392 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1624635492
transform 1 0 48300 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_538
timestamp 1624635492
transform 1 0 50600 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_526
timestamp 1624635492
transform 1 0 49496 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_544
timestamp 1624635492
transform 1 0 51152 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _249_
timestamp 1624635492
transform 1 0 50876 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_94_420
timestamp 1624635492
transform 1 0 39744 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_429
timestamp 1624635492
transform 1 0 40572 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1624635492
transform 1 0 40480 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_441
timestamp 1624635492
transform 1 0 41676 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_453
timestamp 1624635492
transform 1 0 42780 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_465
timestamp 1624635492
transform 1 0 43884 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_486
timestamp 1624635492
transform 1 0 45816 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_477
timestamp 1624635492
transform 1 0 44988 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1624635492
transform 1 0 45724 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_498
timestamp 1624635492
transform 1 0 46920 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_510
timestamp 1624635492
transform 1 0 48024 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_522
timestamp 1624635492
transform 1 0 49128 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_534
timestamp 1624635492
transform 1 0 50232 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_543
timestamp 1624635492
transform 1 0 51060 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1624635492
transform 1 0 50968 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_416
timestamp 1624635492
transform 1 0 39376 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_412
timestamp 1624635492
transform 1 0 39008 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_429
timestamp 1624635492
transform 1 0 40572 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_424
timestamp 1624635492
transform 1 0 40112 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1624635492
transform 1 0 40480 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_441
timestamp 1624635492
transform 1 0 41676 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_448
timestamp 1624635492
transform 1 0 42320 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_436
timestamp 1624635492
transform 1 0 41216 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_453
timestamp 1624635492
transform 1 0 42780 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_457
timestamp 1624635492
transform 1 0 43148 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1624635492
transform 1 0 43056 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_473
timestamp 1624635492
transform 1 0 44620 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_96_465
timestamp 1624635492
transform 1 0 43884 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_469
timestamp 1624635492
transform 1 0 44252 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_486
timestamp 1624635492
transform 1 0 45816 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_484
timestamp 1624635492
transform 1 0 45632 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_478
timestamp 1624635492
transform 1 0 45080 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_481
timestamp 1624635492
transform 1 0 45356 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1624635492
transform 1 0 45724 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _166_
timestamp 1624635492
transform -1 0 45080 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_498
timestamp 1624635492
transform 1 0 46920 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_493
timestamp 1624635492
transform 1 0 46460 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_510
timestamp 1624635492
transform 1 0 48024 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_505
timestamp 1624635492
transform 1 0 47564 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_522
timestamp 1624635492
transform 1 0 49128 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_521
timestamp 1624635492
transform 1 0 49036 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_514
timestamp 1624635492
transform 1 0 48392 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1624635492
transform 1 0 48300 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _182_
timestamp 1624635492
transform -1 0 49036 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_96_534
timestamp 1624635492
transform 1 0 50232 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_533
timestamp 1624635492
transform 1 0 50140 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_543
timestamp 1624635492
transform 1 0 51060 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_545
timestamp 1624635492
transform 1 0 51244 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1624635492
transform 1 0 50968 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_419
timestamp 1624635492
transform 1 0 39652 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_413
timestamp 1624635492
transform 1 0 39100 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B1
timestamp 1624635492
transform 1 0 39468 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_431
timestamp 1624635492
transform 1 0 40756 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_447
timestamp 1624635492
transform 1 0 42228 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_443
timestamp 1624635492
transform 1 0 41860 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _220_
timestamp 1624635492
transform -1 0 42228 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_457
timestamp 1624635492
transform 1 0 43148 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_455
timestamp 1624635492
transform 1 0 42964 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1624635492
transform 1 0 43056 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_469
timestamp 1624635492
transform 1 0 44252 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_481
timestamp 1624635492
transform 1 0 45356 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_493
timestamp 1624635492
transform 1 0 46460 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_505
timestamp 1624635492
transform 1 0 47564 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_514
timestamp 1624635492
transform 1 0 48392 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1624635492
transform 1 0 48300 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_538
timestamp 1624635492
transform 1 0 50600 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_526
timestamp 1624635492
transform 1 0 49496 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_414
timestamp 1624635492
transform 1 0 39192 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_429
timestamp 1624635492
transform 1 0 40572 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_426
timestamp 1624635492
transform 1 0 40296 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1624635492
transform 1 0 40480 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_441
timestamp 1624635492
transform 1 0 41676 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_453
timestamp 1624635492
transform 1 0 42780 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_465
timestamp 1624635492
transform 1 0 43884 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_486
timestamp 1624635492
transform 1 0 45816 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_477
timestamp 1624635492
transform 1 0 44988 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1624635492
transform 1 0 45724 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_498
timestamp 1624635492
transform 1 0 46920 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_510
timestamp 1624635492
transform 1 0 48024 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_522
timestamp 1624635492
transform 1 0 49128 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_534
timestamp 1624635492
transform 1 0 50232 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_543
timestamp 1624635492
transform 1 0 51060 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1624635492
transform 1 0 50968 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_412
timestamp 1624635492
transform 1 0 39008 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_424
timestamp 1624635492
transform 1 0 40112 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_448
timestamp 1624635492
transform 1 0 42320 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_436
timestamp 1624635492
transform 1 0 41216 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_457
timestamp 1624635492
transform 1 0 43148 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1254
timestamp 1624635492
transform 1 0 43056 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_469
timestamp 1624635492
transform 1 0 44252 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_481
timestamp 1624635492
transform 1 0 45356 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_493
timestamp 1624635492
transform 1 0 46460 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_505
timestamp 1624635492
transform 1 0 47564 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_514
timestamp 1624635492
transform 1 0 48392 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1255
timestamp 1624635492
transform 1 0 48300 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_538
timestamp 1624635492
transform 1 0 50600 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_526
timestamp 1624635492
transform 1 0 49496 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_420
timestamp 1624635492
transform 1 0 39744 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_429
timestamp 1624635492
transform 1 0 40572 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1266
timestamp 1624635492
transform 1 0 40480 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_441
timestamp 1624635492
transform 1 0 41676 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_453
timestamp 1624635492
transform 1 0 42780 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_465
timestamp 1624635492
transform 1 0 43884 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_486
timestamp 1624635492
transform 1 0 45816 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_477
timestamp 1624635492
transform 1 0 44988 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1267
timestamp 1624635492
transform 1 0 45724 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_498
timestamp 1624635492
transform 1 0 46920 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_510
timestamp 1624635492
transform 1 0 48024 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_522
timestamp 1624635492
transform 1 0 49128 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_534
timestamp 1624635492
transform 1 0 50232 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_543
timestamp 1624635492
transform 1 0 51060 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1268
timestamp 1624635492
transform 1 0 50968 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_412
timestamp 1624635492
transform 1 0 39008 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_424
timestamp 1624635492
transform 1 0 40112 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_448
timestamp 1624635492
transform 1 0 42320 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_436
timestamp 1624635492
transform 1 0 41216 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_457
timestamp 1624635492
transform 1 0 43148 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1279
timestamp 1624635492
transform 1 0 43056 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_469
timestamp 1624635492
transform 1 0 44252 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_481
timestamp 1624635492
transform 1 0 45356 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_493
timestamp 1624635492
transform 1 0 46460 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_505
timestamp 1624635492
transform 1 0 47564 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_514
timestamp 1624635492
transform 1 0 48392 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1280
timestamp 1624635492
transform 1 0 48300 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_538
timestamp 1624635492
transform 1 0 50600 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_526
timestamp 1624635492
transform 1 0 49496 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_412
timestamp 1624635492
transform 1 0 39008 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_418
timestamp 1624635492
transform 1 0 39560 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_424
timestamp 1624635492
transform 1 0 40112 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_429
timestamp 1624635492
transform 1 0 40572 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_426
timestamp 1624635492
transform 1 0 40296 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1291
timestamp 1624635492
transform 1 0 40480 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_448
timestamp 1624635492
transform 1 0 42320 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_436
timestamp 1624635492
transform 1 0 41216 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_441
timestamp 1624635492
transform 1 0 41676 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_460
timestamp 1624635492
transform 1 0 43424 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_457
timestamp 1624635492
transform 1 0 43148 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_452
timestamp 1624635492
transform 1 0 42688 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_459
timestamp 1624635492
transform 1 0 43332 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_453
timestamp 1624635492
transform 1 0 42780 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B1
timestamp 1624635492
transform -1 0 42688 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A2
timestamp 1624635492
transform 1 0 43424 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A1
timestamp 1624635492
transform 1 0 43240 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1304
timestamp 1624635492
transform 1 0 43056 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_471
timestamp 1624635492
transform 1 0 44436 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_462
timestamp 1624635492
transform 1 0 43608 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _086_
timestamp 1624635492
transform 1 0 43792 0 1 58208
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_103_483
timestamp 1624635492
transform 1 0 45540 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_486
timestamp 1624635492
transform 1 0 45816 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_481
timestamp 1624635492
transform 1 0 45356 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_474
timestamp 1624635492
transform 1 0 44712 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1292
timestamp 1624635492
transform 1 0 45724 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _139_
timestamp 1624635492
transform 1 0 45080 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_495
timestamp 1624635492
transform 1 0 46644 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_498
timestamp 1624635492
transform 1 0 46920 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_507
timestamp 1624635492
transform 1 0 47748 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_102_510
timestamp 1624635492
transform 1 0 48024 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_521
timestamp 1624635492
transform 1 0 49036 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_514
timestamp 1624635492
transform 1 0 48392 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_522
timestamp 1624635492
transform 1 0 49128 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1305
timestamp 1624635492
transform 1 0 48300 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _300_
timestamp 1624635492
transform -1 0 49036 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_533
timestamp 1624635492
transform 1 0 50140 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_534
timestamp 1624635492
transform 1 0 50232 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_545
timestamp 1624635492
transform 1 0 51244 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_543
timestamp 1624635492
transform 1 0 51060 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1293
timestamp 1624635492
transform 1 0 50968 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_420
timestamp 1624635492
transform 1 0 39744 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_429
timestamp 1624635492
transform 1 0 40572 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1316
timestamp 1624635492
transform 1 0 40480 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_441
timestamp 1624635492
transform 1 0 41676 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_460
timestamp 1624635492
transform 1 0 43424 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_457
timestamp 1624635492
transform 1 0 43148 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_453
timestamp 1624635492
transform 1 0 42780 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A3
timestamp 1624635492
transform 1 0 43240 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_104_472
timestamp 1624635492
transform 1 0 44528 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_486
timestamp 1624635492
transform 1 0 45816 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_484
timestamp 1624635492
transform 1 0 45632 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1317
timestamp 1624635492
transform 1 0 45724 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_498
timestamp 1624635492
transform 1 0 46920 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_510
timestamp 1624635492
transform 1 0 48024 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_522
timestamp 1624635492
transform 1 0 49128 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_534
timestamp 1624635492
transform 1 0 50232 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_543
timestamp 1624635492
transform 1 0 51060 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1318
timestamp 1624635492
transform 1 0 50968 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_412
timestamp 1624635492
transform 1 0 39008 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_424
timestamp 1624635492
transform 1 0 40112 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_448
timestamp 1624635492
transform 1 0 42320 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_436
timestamp 1624635492
transform 1 0 41216 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_457
timestamp 1624635492
transform 1 0 43148 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1329
timestamp 1624635492
transform 1 0 43056 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_469
timestamp 1624635492
transform 1 0 44252 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_481
timestamp 1624635492
transform 1 0 45356 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_493
timestamp 1624635492
transform 1 0 46460 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_505
timestamp 1624635492
transform 1 0 47564 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_514
timestamp 1624635492
transform 1 0 48392 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1330
timestamp 1624635492
transform 1 0 48300 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_538
timestamp 1624635492
transform 1 0 50600 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_526
timestamp 1624635492
transform 1 0 49496 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_546
timestamp 1624635492
transform 1 0 51336 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_420
timestamp 1624635492
transform 1 0 39744 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_429
timestamp 1624635492
transform 1 0 40572 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1341
timestamp 1624635492
transform 1 0 40480 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_441
timestamp 1624635492
transform 1 0 41676 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_453
timestamp 1624635492
transform 1 0 42780 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_473
timestamp 1624635492
transform 1 0 44620 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_469
timestamp 1624635492
transform 1 0 44252 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_465
timestamp 1624635492
transform 1 0 43884 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _130_
timestamp 1624635492
transform -1 0 44620 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_486
timestamp 1624635492
transform 1 0 45816 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1342
timestamp 1624635492
transform 1 0 45724 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_498
timestamp 1624635492
transform 1 0 46920 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_506
timestamp 1624635492
transform 1 0 47656 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_502
timestamp 1624635492
transform 1 0 47288 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _168_
timestamp 1624635492
transform -1 0 47656 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_518
timestamp 1624635492
transform 1 0 48760 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_530
timestamp 1624635492
transform 1 0 49864 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_543
timestamp 1624635492
transform 1 0 51060 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1343
timestamp 1624635492
transform 1 0 50968 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_555
timestamp 1624635492
transform 1 0 52164 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_567
timestamp 1624635492
transform 1 0 53268 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_579
timestamp 1624635492
transform 1 0 54372 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_591
timestamp 1624635492
transform 1 0 55476 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_600
timestamp 1624635492
transform 1 0 56304 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1624635492
transform 1 0 56212 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_612
timestamp 1624635492
transform 1 0 57408 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_636
timestamp 1624635492
transform 1 0 59616 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_624
timestamp 1624635492
transform 1 0 58512 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_648
timestamp 1624635492
transform 1 0 60720 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_657
timestamp 1624635492
transform 1 0 61548 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1624635492
transform 1 0 61456 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_669
timestamp 1624635492
transform 1 0 62652 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_681
timestamp 1624635492
transform 1 0 63756 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_550
timestamp 1624635492
transform 1 0 51704 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_571
timestamp 1624635492
transform 1 0 53636 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_562
timestamp 1624635492
transform 1 0 52808 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1624635492
transform 1 0 53544 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_583
timestamp 1624635492
transform 1 0 54740 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_595
timestamp 1624635492
transform 1 0 55844 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_607
timestamp 1624635492
transform 1 0 56948 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_619
timestamp 1624635492
transform 1 0 58052 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_628
timestamp 1624635492
transform 1 0 58880 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1624635492
transform 1 0 58788 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_640
timestamp 1624635492
transform 1 0 59984 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_652
timestamp 1624635492
transform 1 0 61088 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_664
timestamp 1624635492
transform 1 0 62192 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_676
timestamp 1624635492
transform 1 0 63296 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_550
timestamp 1624635492
transform 1 0 51704 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_555
timestamp 1624635492
transform 1 0 52164 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_571
timestamp 1624635492
transform 1 0 53636 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_562
timestamp 1624635492
transform 1 0 52808 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_567
timestamp 1624635492
transform 1 0 53268 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1624635492
transform 1 0 53544 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_583
timestamp 1624635492
transform 1 0 54740 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_579
timestamp 1624635492
transform 1 0 54372 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_595
timestamp 1624635492
transform 1 0 55844 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_591
timestamp 1624635492
transform 1 0 55476 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_607
timestamp 1624635492
transform 1 0 56948 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_600
timestamp 1624635492
transform 1 0 56304 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1624635492
transform 1 0 56212 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_619
timestamp 1624635492
transform 1 0 58052 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_612
timestamp 1624635492
transform 1 0 57408 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_628
timestamp 1624635492
transform 1 0 58880 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_636
timestamp 1624635492
transform 1 0 59616 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_624
timestamp 1624635492
transform 1 0 58512 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1624635492
transform 1 0 58788 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_640
timestamp 1624635492
transform 1 0 59984 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_648
timestamp 1624635492
transform 1 0 60720 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_652
timestamp 1624635492
transform 1 0 61088 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_657
timestamp 1624635492
transform 1 0 61548 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1624635492
transform 1 0 61456 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_664
timestamp 1624635492
transform 1 0 62192 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_669
timestamp 1624635492
transform 1 0 62652 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_676
timestamp 1624635492
transform 1 0 63296 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_681
timestamp 1624635492
transform 1 0 63756 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_555
timestamp 1624635492
transform 1 0 52164 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_567
timestamp 1624635492
transform 1 0 53268 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_579
timestamp 1624635492
transform 1 0 54372 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_591
timestamp 1624635492
transform 1 0 55476 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_600
timestamp 1624635492
transform 1 0 56304 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1624635492
transform 1 0 56212 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_612
timestamp 1624635492
transform 1 0 57408 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_636
timestamp 1624635492
transform 1 0 59616 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_624
timestamp 1624635492
transform 1 0 58512 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_648
timestamp 1624635492
transform 1 0 60720 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_657
timestamp 1624635492
transform 1 0 61548 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1624635492
transform 1 0 61456 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_669
timestamp 1624635492
transform 1 0 62652 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_681
timestamp 1624635492
transform 1 0 63756 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_550
timestamp 1624635492
transform 1 0 51704 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_571
timestamp 1624635492
transform 1 0 53636 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_562
timestamp 1624635492
transform 1 0 52808 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1624635492
transform 1 0 53544 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_583
timestamp 1624635492
transform 1 0 54740 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_595
timestamp 1624635492
transform 1 0 55844 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_607
timestamp 1624635492
transform 1 0 56948 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_619
timestamp 1624635492
transform 1 0 58052 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_628
timestamp 1624635492
transform 1 0 58880 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1624635492
transform 1 0 58788 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_640
timestamp 1624635492
transform 1 0 59984 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_652
timestamp 1624635492
transform 1 0 61088 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_664
timestamp 1624635492
transform 1 0 62192 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_676
timestamp 1624635492
transform 1 0 63296 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_555
timestamp 1624635492
transform 1 0 52164 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_567
timestamp 1624635492
transform 1 0 53268 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_579
timestamp 1624635492
transform 1 0 54372 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_591
timestamp 1624635492
transform 1 0 55476 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_600
timestamp 1624635492
transform 1 0 56304 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1624635492
transform 1 0 56212 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_612
timestamp 1624635492
transform 1 0 57408 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_636
timestamp 1624635492
transform 1 0 59616 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_624
timestamp 1624635492
transform 1 0 58512 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_648
timestamp 1624635492
transform 1 0 60720 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_657
timestamp 1624635492
transform 1 0 61548 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1624635492
transform 1 0 61456 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_669
timestamp 1624635492
transform 1 0 62652 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_681
timestamp 1624635492
transform 1 0 63756 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_550
timestamp 1624635492
transform 1 0 51704 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_571
timestamp 1624635492
transform 1 0 53636 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_562
timestamp 1624635492
transform 1 0 52808 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1624635492
transform 1 0 53544 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_583
timestamp 1624635492
transform 1 0 54740 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_595
timestamp 1624635492
transform 1 0 55844 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_607
timestamp 1624635492
transform 1 0 56948 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_619
timestamp 1624635492
transform 1 0 58052 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_628
timestamp 1624635492
transform 1 0 58880 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1624635492
transform 1 0 58788 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_640
timestamp 1624635492
transform 1 0 59984 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_652
timestamp 1624635492
transform 1 0 61088 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_664
timestamp 1624635492
transform 1 0 62192 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_676
timestamp 1624635492
transform 1 0 63296 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_550
timestamp 1624635492
transform 1 0 51704 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_555
timestamp 1624635492
transform 1 0 52164 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_571
timestamp 1624635492
transform 1 0 53636 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_562
timestamp 1624635492
transform 1 0 52808 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_567
timestamp 1624635492
transform 1 0 53268 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1624635492
transform 1 0 53544 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_578
timestamp 1624635492
transform 1 0 54280 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_579
timestamp 1624635492
transform 1 0 54372 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _106_
timestamp 1624635492
transform 1 0 54004 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_590
timestamp 1624635492
transform 1 0 55384 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_591
timestamp 1624635492
transform 1 0 55476 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_602
timestamp 1624635492
transform 1 0 56488 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_600
timestamp 1624635492
transform 1 0 56304 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1624635492
transform 1 0 56212 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_614
timestamp 1624635492
transform 1 0 57592 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_612
timestamp 1624635492
transform 1 0 57408 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_628
timestamp 1624635492
transform 1 0 58880 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_626
timestamp 1624635492
transform 1 0 58696 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_636
timestamp 1624635492
transform 1 0 59616 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_624
timestamp 1624635492
transform 1 0 58512 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1624635492
transform 1 0 58788 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_640
timestamp 1624635492
transform 1 0 59984 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_648
timestamp 1624635492
transform 1 0 60720 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_652
timestamp 1624635492
transform 1 0 61088 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_657
timestamp 1624635492
transform 1 0 61548 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1624635492
transform 1 0 61456 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_664
timestamp 1624635492
transform 1 0 62192 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_669
timestamp 1624635492
transform 1 0 62652 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_676
timestamp 1624635492
transform 1 0 63296 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_681
timestamp 1624635492
transform 1 0 63756 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_555
timestamp 1624635492
transform 1 0 52164 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_567
timestamp 1624635492
transform 1 0 53268 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_579
timestamp 1624635492
transform 1 0 54372 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_591
timestamp 1624635492
transform 1 0 55476 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_600
timestamp 1624635492
transform 1 0 56304 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1624635492
transform 1 0 56212 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_612
timestamp 1624635492
transform 1 0 57408 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_636
timestamp 1624635492
transform 1 0 59616 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_624
timestamp 1624635492
transform 1 0 58512 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_648
timestamp 1624635492
transform 1 0 60720 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_657
timestamp 1624635492
transform 1 0 61548 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1624635492
transform 1 0 61456 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_669
timestamp 1624635492
transform 1 0 62652 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_681
timestamp 1624635492
transform 1 0 63756 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_550
timestamp 1624635492
transform 1 0 51704 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_571
timestamp 1624635492
transform 1 0 53636 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_562
timestamp 1624635492
transform 1 0 52808 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1624635492
transform 1 0 53544 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_583
timestamp 1624635492
transform 1 0 54740 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_595
timestamp 1624635492
transform 1 0 55844 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_607
timestamp 1624635492
transform 1 0 56948 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_619
timestamp 1624635492
transform 1 0 58052 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_628
timestamp 1624635492
transform 1 0 58880 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1624635492
transform 1 0 58788 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_640
timestamp 1624635492
transform 1 0 59984 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_652
timestamp 1624635492
transform 1 0 61088 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_664
timestamp 1624635492
transform 1 0 62192 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_676
timestamp 1624635492
transform 1 0 63296 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_555
timestamp 1624635492
transform 1 0 52164 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_567
timestamp 1624635492
transform 1 0 53268 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_92_577
timestamp 1624635492
transform 1 0 54188 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A2
timestamp 1624635492
transform 1 0 54004 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_590
timestamp 1624635492
transform 1 0 55384 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_585
timestamp 1624635492
transform 1 0 54924 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B1
timestamp 1624635492
transform 1 0 55200 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_600
timestamp 1624635492
transform 1 0 56304 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_598
timestamp 1624635492
transform 1 0 56120 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1624635492
transform 1 0 56212 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_612
timestamp 1624635492
transform 1 0 57408 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_636
timestamp 1624635492
transform 1 0 59616 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_624
timestamp 1624635492
transform 1 0 58512 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_648
timestamp 1624635492
transform 1 0 60720 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_657
timestamp 1624635492
transform 1 0 61548 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1624635492
transform 1 0 61456 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_669
timestamp 1624635492
transform 1 0 62652 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_92_677
timestamp 1624635492
transform 1 0 63388 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1624635492
transform 1 0 63204 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_556
timestamp 1624635492
transform 1 0 52256 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_571
timestamp 1624635492
transform 1 0 53636 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_566
timestamp 1624635492
transform 1 0 53176 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__C1
timestamp 1624635492
transform -1 0 53176 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1624635492
transform 1 0 53544 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_575
timestamp 1624635492
transform 1 0 54004 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A1
timestamp 1624635492
transform -1 0 54004 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_2  _075_
timestamp 1624635492
transform -1 0 55200 0 1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_93_596
timestamp 1624635492
transform 1 0 55936 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_588
timestamp 1624635492
transform 1 0 55200 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _331_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 55568 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_608
timestamp 1624635492
transform 1 0 57040 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_620
timestamp 1624635492
transform 1 0 58144 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_628
timestamp 1624635492
transform 1 0 58880 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_626
timestamp 1624635492
transform 1 0 58696 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1624635492
transform 1 0 58788 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_640
timestamp 1624635492
transform 1 0 59984 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_652
timestamp 1624635492
transform 1 0 61088 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_664
timestamp 1624635492
transform 1 0 62192 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__inv_4  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 63204 0 1 52768
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_93_675
timestamp 1624635492
transform 1 0 63204 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_555
timestamp 1624635492
transform 1 0 52164 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_567
timestamp 1624635492
transform 1 0 53268 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_575
timestamp 1624635492
transform 1 0 54004 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A3
timestamp 1624635492
transform -1 0 54004 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_592
timestamp 1624635492
transform 1 0 55568 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_94_587
timestamp 1624635492
transform 1 0 55108 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1624635492
transform 1 0 55384 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_600
timestamp 1624635492
transform 1 0 56304 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_598
timestamp 1624635492
transform 1 0 56120 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1624635492
transform 1 0 56212 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_612
timestamp 1624635492
transform 1 0 57408 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_636
timestamp 1624635492
transform 1 0 59616 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_624
timestamp 1624635492
transform 1 0 58512 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_648
timestamp 1624635492
transform 1 0 60720 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_657
timestamp 1624635492
transform 1 0 61548 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1624635492
transform 1 0 61456 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_669
timestamp 1624635492
transform 1 0 62652 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_681
timestamp 1624635492
transform 1 0 63756 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_555
timestamp 1624635492
transform 1 0 52164 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_557
timestamp 1624635492
transform 1 0 52348 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_567
timestamp 1624635492
transform 1 0 53268 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_571
timestamp 1624635492
transform 1 0 53636 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_569
timestamp 1624635492
transform 1 0 53452 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1624635492
transform 1 0 53544 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_579
timestamp 1624635492
transform 1 0 54372 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_583
timestamp 1624635492
transform 1 0 54740 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_591
timestamp 1624635492
transform 1 0 55476 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_595
timestamp 1624635492
transform 1 0 55844 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_600
timestamp 1624635492
transform 1 0 56304 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_607
timestamp 1624635492
transform 1 0 56948 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1624635492
transform 1 0 56212 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_612
timestamp 1624635492
transform 1 0 57408 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_619
timestamp 1624635492
transform 1 0 58052 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_636
timestamp 1624635492
transform 1 0 59616 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_624
timestamp 1624635492
transform 1 0 58512 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_628
timestamp 1624635492
transform 1 0 58880 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1624635492
transform 1 0 58788 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_648
timestamp 1624635492
transform 1 0 60720 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_640
timestamp 1624635492
transform 1 0 59984 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_657
timestamp 1624635492
transform 1 0 61548 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_652
timestamp 1624635492
transform 1 0 61088 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1624635492
transform 1 0 61456 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _283_
timestamp 1624635492
transform 1 0 61916 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_664
timestamp 1624635492
transform 1 0 62192 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_664
timestamp 1624635492
transform 1 0 62192 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_676
timestamp 1624635492
transform 1 0 63296 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_676
timestamp 1624635492
transform 1 0 63296 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_550
timestamp 1624635492
transform 1 0 51704 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_571
timestamp 1624635492
transform 1 0 53636 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_562
timestamp 1624635492
transform 1 0 52808 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1624635492
transform 1 0 53544 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_583
timestamp 1624635492
transform 1 0 54740 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_595
timestamp 1624635492
transform 1 0 55844 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_607
timestamp 1624635492
transform 1 0 56948 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_619
timestamp 1624635492
transform 1 0 58052 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_628
timestamp 1624635492
transform 1 0 58880 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1624635492
transform 1 0 58788 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_648
timestamp 1624635492
transform 1 0 60720 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_640
timestamp 1624635492
transform 1 0 59984 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_653
timestamp 1624635492
transform 1 0 61180 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _145_
timestamp 1624635492
transform 1 0 60904 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_665
timestamp 1624635492
transform 1 0 62284 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_677
timestamp 1624635492
transform 1 0 63388 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_555
timestamp 1624635492
transform 1 0 52164 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_567
timestamp 1624635492
transform 1 0 53268 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_579
timestamp 1624635492
transform 1 0 54372 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_591
timestamp 1624635492
transform 1 0 55476 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_600
timestamp 1624635492
transform 1 0 56304 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1244
timestamp 1624635492
transform 1 0 56212 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_612
timestamp 1624635492
transform 1 0 57408 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_636
timestamp 1624635492
transform 1 0 59616 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_624
timestamp 1624635492
transform 1 0 58512 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_648
timestamp 1624635492
transform 1 0 60720 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_657
timestamp 1624635492
transform 1 0 61548 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1245
timestamp 1624635492
transform 1 0 61456 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_669
timestamp 1624635492
transform 1 0 62652 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_681
timestamp 1624635492
transform 1 0 63756 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_550
timestamp 1624635492
transform 1 0 51704 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_571
timestamp 1624635492
transform 1 0 53636 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_562
timestamp 1624635492
transform 1 0 52808 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1256
timestamp 1624635492
transform 1 0 53544 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_583
timestamp 1624635492
transform 1 0 54740 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_595
timestamp 1624635492
transform 1 0 55844 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_607
timestamp 1624635492
transform 1 0 56948 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_619
timestamp 1624635492
transform 1 0 58052 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_628
timestamp 1624635492
transform 1 0 58880 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1257
timestamp 1624635492
transform 1 0 58788 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_640
timestamp 1624635492
transform 1 0 59984 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_652
timestamp 1624635492
transform 1 0 61088 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_664
timestamp 1624635492
transform 1 0 62192 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_676
timestamp 1624635492
transform 1 0 63296 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_555
timestamp 1624635492
transform 1 0 52164 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_567
timestamp 1624635492
transform 1 0 53268 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_579
timestamp 1624635492
transform 1 0 54372 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_591
timestamp 1624635492
transform 1 0 55476 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_600
timestamp 1624635492
transform 1 0 56304 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1269
timestamp 1624635492
transform 1 0 56212 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_612
timestamp 1624635492
transform 1 0 57408 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_636
timestamp 1624635492
transform 1 0 59616 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_624
timestamp 1624635492
transform 1 0 58512 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_648
timestamp 1624635492
transform 1 0 60720 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_657
timestamp 1624635492
transform 1 0 61548 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1270
timestamp 1624635492
transform 1 0 61456 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_669
timestamp 1624635492
transform 1 0 62652 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_681
timestamp 1624635492
transform 1 0 63756 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_550
timestamp 1624635492
transform 1 0 51704 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_571
timestamp 1624635492
transform 1 0 53636 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_562
timestamp 1624635492
transform 1 0 52808 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1281
timestamp 1624635492
transform 1 0 53544 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_583
timestamp 1624635492
transform 1 0 54740 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_595
timestamp 1624635492
transform 1 0 55844 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_607
timestamp 1624635492
transform 1 0 56948 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_619
timestamp 1624635492
transform 1 0 58052 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_628
timestamp 1624635492
transform 1 0 58880 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1282
timestamp 1624635492
transform 1 0 58788 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_640
timestamp 1624635492
transform 1 0 59984 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_652
timestamp 1624635492
transform 1 0 61088 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_664
timestamp 1624635492
transform 1 0 62192 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_676
timestamp 1624635492
transform 1 0 63296 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_557
timestamp 1624635492
transform 1 0 52348 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_555
timestamp 1624635492
transform 1 0 52164 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_571
timestamp 1624635492
transform 1 0 53636 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_569
timestamp 1624635492
transform 1 0 53452 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_567
timestamp 1624635492
transform 1 0 53268 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1306
timestamp 1624635492
transform 1 0 53544 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_583
timestamp 1624635492
transform 1 0 54740 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_579
timestamp 1624635492
transform 1 0 54372 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_595
timestamp 1624635492
transform 1 0 55844 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_590
timestamp 1624635492
transform 1 0 55384 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _185_
timestamp 1624635492
transform -1 0 55384 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_607
timestamp 1624635492
transform 1 0 56948 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_600
timestamp 1624635492
transform 1 0 56304 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_598
timestamp 1624635492
transform 1 0 56120 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1294
timestamp 1624635492
transform 1 0 56212 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_619
timestamp 1624635492
transform 1 0 58052 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_612
timestamp 1624635492
transform 1 0 57408 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_628
timestamp 1624635492
transform 1 0 58880 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_636
timestamp 1624635492
transform 1 0 59616 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_624
timestamp 1624635492
transform 1 0 58512 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1307
timestamp 1624635492
transform 1 0 58788 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_640
timestamp 1624635492
transform 1 0 59984 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_648
timestamp 1624635492
transform 1 0 60720 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_652
timestamp 1624635492
transform 1 0 61088 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_657
timestamp 1624635492
transform 1 0 61548 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1295
timestamp 1624635492
transform 1 0 61456 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_664
timestamp 1624635492
transform 1 0 62192 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_669
timestamp 1624635492
transform 1 0 62652 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_676
timestamp 1624635492
transform 1 0 63296 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_102_681
timestamp 1624635492
transform 1 0 63756 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_104_555
timestamp 1624635492
transform 1 0 52164 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_567
timestamp 1624635492
transform 1 0 53268 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_579
timestamp 1624635492
transform 1 0 54372 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_591
timestamp 1624635492
transform 1 0 55476 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_600
timestamp 1624635492
transform 1 0 56304 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1319
timestamp 1624635492
transform 1 0 56212 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_612
timestamp 1624635492
transform 1 0 57408 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_636
timestamp 1624635492
transform 1 0 59616 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_624
timestamp 1624635492
transform 1 0 58512 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_648
timestamp 1624635492
transform 1 0 60720 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_657
timestamp 1624635492
transform 1 0 61548 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1320
timestamp 1624635492
transform 1 0 61456 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_669
timestamp 1624635492
transform 1 0 62652 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_681
timestamp 1624635492
transform 1 0 63756 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_105_559
timestamp 1624635492
transform 1 0 52532 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_105_551
timestamp 1624635492
transform 1 0 51796 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__B1
timestamp 1624635492
transform 1 0 51612 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_571
timestamp 1624635492
transform 1 0 53636 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_569
timestamp 1624635492
transform 1 0 53452 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_105_563
timestamp 1624635492
transform 1 0 52900 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A1
timestamp 1624635492
transform 1 0 52716 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1331
timestamp 1624635492
transform 1 0 53544 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_583
timestamp 1624635492
transform 1 0 54740 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_595
timestamp 1624635492
transform 1 0 55844 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_607
timestamp 1624635492
transform 1 0 56948 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_619
timestamp 1624635492
transform 1 0 58052 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_628
timestamp 1624635492
transform 1 0 58880 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1332
timestamp 1624635492
transform 1 0 58788 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_640
timestamp 1624635492
transform 1 0 59984 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_652
timestamp 1624635492
transform 1 0 61088 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_664
timestamp 1624635492
transform 1 0 62192 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_676
timestamp 1624635492
transform 1 0 63296 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_106_549
timestamp 1624635492
transform 1 0 51612 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A2
timestamp 1624635492
transform 1 0 51428 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _060_
timestamp 1624635492
transform -1 0 52716 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_569
timestamp 1624635492
transform 1 0 53452 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_565
timestamp 1624635492
transform 1 0 53084 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_561
timestamp 1624635492
transform 1 0 52716 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _223_
timestamp 1624635492
transform -1 0 53452 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_581
timestamp 1624635492
transform 1 0 54556 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_593
timestamp 1624635492
transform 1 0 55660 0 -1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_608
timestamp 1624635492
transform 1 0 57040 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_600
timestamp 1624635492
transform 1 0 56304 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1344
timestamp 1624635492
transform 1 0 56212 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _119_
timestamp 1624635492
transform -1 0 57408 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_612
timestamp 1624635492
transform 1 0 57408 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_636
timestamp 1624635492
transform 1 0 59616 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_624
timestamp 1624635492
transform 1 0 58512 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_648
timestamp 1624635492
transform 1 0 60720 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_657
timestamp 1624635492
transform 1 0 61548 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1345
timestamp 1624635492
transform 1 0 61456 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_669
timestamp 1624635492
transform 1 0 62652 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_681
timestamp 1624635492
transform 1 0 63756 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_685
timestamp 1624635492
transform 1 0 64124 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_693
timestamp 1624635492
transform 1 0 64860 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1624635492
transform 1 0 64032 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_697
timestamp 1624635492
transform 1 0 65228 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_705
timestamp 1624635492
transform 1 0 65964 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_721
timestamp 1624635492
transform 1 0 67436 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_709
timestamp 1624635492
transform 1 0 66332 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_714
timestamp 1624635492
transform 1 0 66792 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1624635492
transform 1 0 66700 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_732
timestamp 1624635492
transform 1 0 68448 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_726
timestamp 1624635492
transform 1 0 67896 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1624635492
transform -1 0 68816 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1624635492
transform -1 0 68816 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_693
timestamp 1624635492
transform 1 0 64860 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_705
timestamp 1624635492
transform 1 0 65964 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_721
timestamp 1624635492
transform 1 0 67436 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_718
timestamp 1624635492
transform 1 0 67160 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_714
timestamp 1624635492
transform 1 0 66792 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output407_A
timestamp 1624635492
transform 1 0 67252 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1624635492
transform 1 0 66700 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_729
timestamp 1624635492
transform 1 0 68172 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output407
timestamp 1624635492
transform 1 0 67804 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1624635492
transform -1 0 68816 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_685
timestamp 1624635492
transform 1 0 64124 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1624635492
transform 1 0 64032 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_697
timestamp 1624635492
transform 1 0 65228 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_721
timestamp 1624635492
transform 1 0 67436 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_709
timestamp 1624635492
transform 1 0 66332 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1624635492
transform -1 0 68816 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_685
timestamp 1624635492
transform 1 0 64124 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_693
timestamp 1624635492
transform 1 0 64860 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1624635492
transform 1 0 64032 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_697
timestamp 1624635492
transform 1 0 65228 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_705
timestamp 1624635492
transform 1 0 65964 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_721
timestamp 1624635492
transform 1 0 67436 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_709
timestamp 1624635492
transform 1 0 66332 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_714
timestamp 1624635492
transform 1 0 66792 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1624635492
transform 1 0 66700 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_729
timestamp 1624635492
transform 1 0 68172 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_84_722
timestamp 1624635492
transform 1 0 67528 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output369
timestamp 1624635492
transform 1 0 67804 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1624635492
transform -1 0 68816 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1624635492
transform -1 0 68816 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_693
timestamp 1624635492
transform 1 0 64860 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_705
timestamp 1624635492
transform 1 0 65964 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_714
timestamp 1624635492
transform 1 0 66792 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1624635492
transform 1 0 66700 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_732
timestamp 1624635492
transform 1 0 68448 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_726
timestamp 1624635492
transform 1 0 67896 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1624635492
transform -1 0 68816 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_693
timestamp 1624635492
transform 1 0 64860 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_685
timestamp 1624635492
transform 1 0 64124 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1624635492
transform 1 0 64032 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_705
timestamp 1624635492
transform 1 0 65964 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_697
timestamp 1624635492
transform 1 0 65228 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_714
timestamp 1624635492
transform 1 0 66792 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_721
timestamp 1624635492
transform 1 0 67436 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_709
timestamp 1624635492
transform 1 0 66332 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1624635492
transform 1 0 66700 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_732
timestamp 1624635492
transform 1 0 68448 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_726
timestamp 1624635492
transform 1 0 67896 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1624635492
transform -1 0 68816 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1624635492
transform -1 0 68816 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_685
timestamp 1624635492
transform 1 0 64124 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1624635492
transform 1 0 64032 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_697
timestamp 1624635492
transform 1 0 65228 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_717
timestamp 1624635492
transform 1 0 67068 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_709
timestamp 1624635492
transform 1 0 66332 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 67528 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1624635492
transform 1 0 68172 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_722
timestamp 1624635492
transform 1 0 67528 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform -1 0 68172 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1624635492
transform -1 0 68816 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_693
timestamp 1624635492
transform 1 0 64860 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_705
timestamp 1624635492
transform 1 0 65964 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_90_714
timestamp 1624635492
transform 1 0 66792 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1624635492
transform 1 0 66700 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _165_
timestamp 1624635492
transform -1 0 67620 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_90_731
timestamp 1624635492
transform 1 0 68356 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_90_723
timestamp 1624635492
transform 1 0 67620 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1624635492
transform -1 0 68816 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_689
timestamp 1624635492
transform 1 0 64492 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_685
timestamp 1624635492
transform 1 0 64124 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1624635492
transform 1 0 64032 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_701
timestamp 1624635492
transform 1 0 65596 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_697
timestamp 1624635492
transform 1 0 65228 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_714
timestamp 1624635492
transform 1 0 66792 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_721
timestamp 1624635492
transform 1 0 67436 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_717
timestamp 1624635492
transform 1 0 67068 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_709
timestamp 1624635492
transform 1 0 66332 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output408_A
timestamp 1624635492
transform 1 0 67252 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1624635492
transform 1 0 66700 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_732
timestamp 1624635492
transform 1 0 68448 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_726
timestamp 1624635492
transform 1 0 67896 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1624635492
transform 1 0 68172 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output408
timestamp 1624635492
transform 1 0 67804 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1624635492
transform -1 0 68816 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1624635492
transform -1 0 68816 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_685
timestamp 1624635492
transform 1 0 64124 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_683
timestamp 1624635492
transform 1 0 63940 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1624635492
transform 1 0 64032 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_700
timestamp 1624635492
transform 1 0 65504 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _201_
timestamp 1624635492
transform -1 0 65504 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_712
timestamp 1624635492
transform 1 0 66608 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_732
timestamp 1624635492
transform 1 0 68448 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_724
timestamp 1624635492
transform 1 0 67712 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1624635492
transform -1 0 68816 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_685
timestamp 1624635492
transform 1 0 64124 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_693
timestamp 1624635492
transform 1 0 64860 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1624635492
transform 1 0 64032 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_697
timestamp 1624635492
transform 1 0 65228 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_705
timestamp 1624635492
transform 1 0 65964 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_721
timestamp 1624635492
transform 1 0 67436 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_709
timestamp 1624635492
transform 1 0 66332 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_721
timestamp 1624635492
transform 1 0 67436 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_718
timestamp 1624635492
transform 1 0 67160 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_714
timestamp 1624635492
transform 1 0 66792 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output370_A
timestamp 1624635492
transform 1 0 67252 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1624635492
transform 1 0 66700 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_729
timestamp 1624635492
transform 1 0 68172 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output370
timestamp 1624635492
transform 1 0 67804 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1624635492
transform -1 0 68816 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1624635492
transform -1 0 68816 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_688
timestamp 1624635492
transform 1 0 64400 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_700
timestamp 1624635492
transform 1 0 65504 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_714
timestamp 1624635492
transform 1 0 66792 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_712
timestamp 1624635492
transform 1 0 66608 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1624635492
transform 1 0 66700 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_732
timestamp 1624635492
transform 1 0 68448 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_726
timestamp 1624635492
transform 1 0 67896 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1624635492
transform -1 0 68816 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_685
timestamp 1624635492
transform 1 0 64124 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_683
timestamp 1624635492
transform 1 0 63940 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1624635492
transform 1 0 64032 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_697
timestamp 1624635492
transform 1 0 65228 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_721
timestamp 1624635492
transform 1 0 67436 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_717
timestamp 1624635492
transform 1 0 67068 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_709
timestamp 1624635492
transform 1 0 66332 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _252_
timestamp 1624635492
transform -1 0 67436 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1624635492
transform -1 0 68816 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_685
timestamp 1624635492
transform 1 0 64124 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_693
timestamp 1624635492
transform 1 0 64860 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1258
timestamp 1624635492
transform 1 0 64032 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_697
timestamp 1624635492
transform 1 0 65228 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_705
timestamp 1624635492
transform 1 0 65964 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_717
timestamp 1624635492
transform 1 0 67068 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_709
timestamp 1624635492
transform 1 0 66332 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_714
timestamp 1624635492
transform 1 0 66792 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 67528 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1246
timestamp 1624635492
transform 1 0 66700 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1624635492
transform 1 0 68172 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_722
timestamp 1624635492
transform 1 0 67528 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_732
timestamp 1624635492
transform 1 0 68448 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_726
timestamp 1624635492
transform 1 0 67896 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform -1 0 68172 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1624635492
transform -1 0 68816 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1624635492
transform -1 0 68816 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_693
timestamp 1624635492
transform 1 0 64860 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_705
timestamp 1624635492
transform 1 0 65964 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_714
timestamp 1624635492
transform 1 0 66792 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1271
timestamp 1624635492
transform 1 0 66700 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_732
timestamp 1624635492
transform 1 0 68448 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_726
timestamp 1624635492
transform 1 0 67896 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1624635492
transform -1 0 68816 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_102_690
timestamp 1624635492
transform 1 0 64584 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_687
timestamp 1624635492
transform 1 0 64308 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_685
timestamp 1624635492
transform 1 0 64124 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__A
timestamp 1624635492
transform 1 0 64400 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1283
timestamp 1624635492
transform 1 0 64032 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _053_
timestamp 1624635492
transform 1 0 64952 0 -1 58208
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_102_703
timestamp 1624635492
transform 1 0 65780 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_697
timestamp 1624635492
transform 1 0 65228 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_714
timestamp 1624635492
transform 1 0 66792 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_711
timestamp 1624635492
transform 1 0 66516 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_721
timestamp 1624635492
transform 1 0 67436 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_717
timestamp 1624635492
transform 1 0 67068 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_709
timestamp 1624635492
transform 1 0 66332 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output409_A
timestamp 1624635492
transform 1 0 67252 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1296
timestamp 1624635492
transform 1 0 66700 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_102_732
timestamp 1624635492
transform 1 0 68448 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_726
timestamp 1624635492
transform 1 0 67896 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1624635492
transform 1 0 68172 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output409
timestamp 1624635492
transform 1 0 67804 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1624635492
transform -1 0 68816 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1624635492
transform -1 0 68816 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_685
timestamp 1624635492
transform 1 0 64124 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1308
timestamp 1624635492
transform 1 0 64032 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_697
timestamp 1624635492
transform 1 0 65228 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_721
timestamp 1624635492
transform 1 0 67436 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_103_717
timestamp 1624635492
transform 1 0 67068 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_103_709
timestamp 1624635492
transform 1 0 66332 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output371_A
timestamp 1624635492
transform -1 0 67436 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_729
timestamp 1624635492
transform 1 0 68172 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output371
timestamp 1624635492
transform 1 0 67804 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1624635492
transform -1 0 68816 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_690
timestamp 1624635492
transform 1 0 64584 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _241_
timestamp 1624635492
transform -1 0 64584 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_104_702
timestamp 1624635492
transform 1 0 65688 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_714
timestamp 1624635492
transform 1 0 66792 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_104_710
timestamp 1624635492
transform 1 0 66424 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1321
timestamp 1624635492
transform 1 0 66700 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_732
timestamp 1624635492
transform 1 0 68448 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_726
timestamp 1624635492
transform 1 0 67896 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1624635492
transform -1 0 68816 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_693
timestamp 1624635492
transform 1 0 64860 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_685
timestamp 1624635492
transform 1 0 64124 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1333
timestamp 1624635492
transform 1 0 64032 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_705
timestamp 1624635492
transform 1 0 65964 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_697
timestamp 1624635492
transform 1 0 65228 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_714
timestamp 1624635492
transform 1 0 66792 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_718
timestamp 1624635492
transform 1 0 67160 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_709
timestamp 1624635492
transform 1 0 66332 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1346
timestamp 1624635492
transform 1 0 66700 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _111_
timestamp 1624635492
transform 1 0 66884 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_106_732
timestamp 1624635492
transform 1 0 68448 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_106_726
timestamp 1624635492
transform 1 0 67896 0 -1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_105_730
timestamp 1624635492
transform 1 0 68264 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1624635492
transform -1 0 68816 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1624635492
transform -1 0 68816 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_15
timestamp 1624635492
transform 1 0 2484 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_3
timestamp 1624635492
transform 1 0 1380 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1624635492
transform 1 0 1104 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_39
timestamp 1624635492
transform 1 0 4692 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_27
timestamp 1624635492
transform 1 0 3588 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_58
timestamp 1624635492
transform 1 0 6440 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_51
timestamp 1624635492
transform 1 0 5796 0 1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1347
timestamp 1624635492
transform 1 0 6348 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_70
timestamp 1624635492
transform 1 0 7544 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_94
timestamp 1624635492
transform 1 0 9752 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_82
timestamp 1624635492
transform 1 0 8648 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_115
timestamp 1624635492
transform 1 0 11684 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_106
timestamp 1624635492
transform 1 0 10856 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1348
timestamp 1624635492
transform 1 0 11592 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_127
timestamp 1624635492
transform 1 0 12788 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1624635492
transform 1 0 2484 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1624635492
transform 1 0 1380 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1624635492
transform 1 0 1104 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_30
timestamp 1624635492
transform 1 0 3864 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_108_27
timestamp 1624635492
transform 1 0 3588 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1359
timestamp 1624635492
transform 1 0 3772 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_54
timestamp 1624635492
transform 1 0 6072 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_42
timestamp 1624635492
transform 1 0 4968 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_78
timestamp 1624635492
transform 1 0 8280 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_66
timestamp 1624635492
transform 1 0 7176 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_99
timestamp 1624635492
transform 1 0 10212 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_87
timestamp 1624635492
transform 1 0 9108 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1360
timestamp 1624635492
transform 1 0 9016 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_111
timestamp 1624635492
transform 1 0 11316 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_135
timestamp 1624635492
transform 1 0 13524 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_123
timestamp 1624635492
transform 1 0 12420 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_17
timestamp 1624635492
transform 1 0 2668 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_11
timestamp 1624635492
transform 1 0 2116 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_3
timestamp 1624635492
transform 1 0 1380 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output423_A
timestamp 1624635492
transform -1 0 2668 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output423
timestamp 1624635492
transform -1 0 2116 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1624635492
transform 1 0 1104 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_29
timestamp 1624635492
transform 1 0 3772 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_58
timestamp 1624635492
transform 1 0 6440 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_53
timestamp 1624635492
transform 1 0 5980 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_41
timestamp 1624635492
transform 1 0 4876 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1372
timestamp 1624635492
transform 1 0 6348 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_70
timestamp 1624635492
transform 1 0 7544 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_94
timestamp 1624635492
transform 1 0 9752 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_82
timestamp 1624635492
transform 1 0 8648 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_115
timestamp 1624635492
transform 1 0 11684 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_106
timestamp 1624635492
transform 1 0 10856 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1373
timestamp 1624635492
transform 1 0 11592 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_127
timestamp 1624635492
transform 1 0 12788 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1624635492
transform 1 0 2484 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1624635492
transform 1 0 1380 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1624635492
transform 1 0 1104 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_30
timestamp 1624635492
transform 1 0 3864 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_110_27
timestamp 1624635492
transform 1 0 3588 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1384
timestamp 1624635492
transform 1 0 3772 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_54
timestamp 1624635492
transform 1 0 6072 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_42
timestamp 1624635492
transform 1 0 4968 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_78
timestamp 1624635492
transform 1 0 8280 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_66
timestamp 1624635492
transform 1 0 7176 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_99
timestamp 1624635492
transform 1 0 10212 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_87
timestamp 1624635492
transform 1 0 9108 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1385
timestamp 1624635492
transform 1 0 9016 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_111
timestamp 1624635492
transform 1 0 11316 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_136
timestamp 1624635492
transform 1 0 13616 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_110_131
timestamp 1624635492
transform 1 0 13156 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_110_123
timestamp 1624635492
transform 1 0 12420 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _256_
timestamp 1624635492
transform 1 0 13340 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_15
timestamp 1624635492
transform 1 0 2484 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_3
timestamp 1624635492
transform 1 0 1380 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_12
timestamp 1624635492
transform 1 0 2208 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_6
timestamp 1624635492
transform 1 0 1656 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 2208 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1624635492
transform -1 0 1656 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1624635492
transform 1 0 1104 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1624635492
transform 1 0 1104 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_30
timestamp 1624635492
transform 1 0 3864 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_112_27
timestamp 1624635492
transform 1 0 3588 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_36
timestamp 1624635492
transform 1 0 4416 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_24
timestamp 1624635492
transform 1 0 3312 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1409
timestamp 1624635492
transform 1 0 3772 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_54
timestamp 1624635492
transform 1 0 6072 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_42
timestamp 1624635492
transform 1 0 4968 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_58
timestamp 1624635492
transform 1 0 6440 0 1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_56
timestamp 1624635492
transform 1 0 6256 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_48
timestamp 1624635492
transform 1 0 5520 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1397
timestamp 1624635492
transform 1 0 6348 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_78
timestamp 1624635492
transform 1 0 8280 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_66
timestamp 1624635492
transform 1 0 7176 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_79
timestamp 1624635492
transform 1 0 8372 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_67
timestamp 1624635492
transform 1 0 7268 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _132_
timestamp 1624635492
transform -1 0 7268 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_112_99
timestamp 1624635492
transform 1 0 10212 0 -1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_112_87
timestamp 1624635492
transform 1 0 9108 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_95
timestamp 1624635492
transform 1 0 9844 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_91
timestamp 1624635492
transform 1 0 9476 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1410
timestamp 1624635492
transform 1 0 9016 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _284_
timestamp 1624635492
transform 1 0 9568 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_115
timestamp 1624635492
transform 1 0 11684 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_113
timestamp 1624635492
transform 1 0 11500 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_111_107
timestamp 1624635492
transform 1 0 10948 0 1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1398
timestamp 1624635492
transform 1 0 11592 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_8  _050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 10764 0 -1 63648
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_112_133
timestamp 1624635492
transform 1 0 13340 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_112_127
timestamp 1624635492
transform 1 0 12788 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_121
timestamp 1624635492
transform 1 0 12236 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_127
timestamp 1624635492
transform 1 0 12788 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__B
timestamp 1624635492
transform 1 0 13156 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__A
timestamp 1624635492
transform 1 0 12604 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1624635492
transform 1 0 2484 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1624635492
transform 1 0 1380 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1624635492
transform 1 0 1104 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_39
timestamp 1624635492
transform 1 0 4692 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1624635492
transform 1 0 3588 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_58
timestamp 1624635492
transform 1 0 6440 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_51
timestamp 1624635492
transform 1 0 5796 0 1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1422
timestamp 1624635492
transform 1 0 6348 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_70
timestamp 1624635492
transform 1 0 7544 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_94
timestamp 1624635492
transform 1 0 9752 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_82
timestamp 1624635492
transform 1 0 8648 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_115
timestamp 1624635492
transform 1 0 11684 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_113_106
timestamp 1624635492
transform 1 0 10856 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1423
timestamp 1624635492
transform 1 0 11592 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_113_123
timestamp 1624635492
transform 1 0 12420 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _350_
timestamp 1624635492
transform -1 0 14352 0 1 63648
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_114_13
timestamp 1624635492
transform 1 0 2300 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_9
timestamp 1624635492
transform 1 0 1932 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_3
timestamp 1624635492
transform 1 0 1380 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1624635492
transform 1 0 1104 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _218_
timestamp 1624635492
transform 1 0 2024 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_30
timestamp 1624635492
transform 1 0 3864 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_25
timestamp 1624635492
transform 1 0 3404 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1434
timestamp 1624635492
transform 1 0 3772 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_54
timestamp 1624635492
transform 1 0 6072 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_42
timestamp 1624635492
transform 1 0 4968 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_78
timestamp 1624635492
transform 1 0 8280 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_66
timestamp 1624635492
transform 1 0 7176 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_99
timestamp 1624635492
transform 1 0 10212 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_87
timestamp 1624635492
transform 1 0 9108 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1435
timestamp 1624635492
transform 1 0 9016 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_111
timestamp 1624635492
transform 1 0 11316 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_135
timestamp 1624635492
transform 1 0 13524 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_123
timestamp 1624635492
transform 1 0 12420 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_15
timestamp 1624635492
transform 1 0 2484 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_3
timestamp 1624635492
transform 1 0 1380 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1624635492
transform 1 0 1104 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_39
timestamp 1624635492
transform 1 0 4692 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_27
timestamp 1624635492
transform 1 0 3588 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_58
timestamp 1624635492
transform 1 0 6440 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_51
timestamp 1624635492
transform 1 0 5796 0 1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1447
timestamp 1624635492
transform 1 0 6348 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_70
timestamp 1624635492
transform 1 0 7544 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_94
timestamp 1624635492
transform 1 0 9752 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_82
timestamp 1624635492
transform 1 0 8648 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_115
timestamp 1624635492
transform 1 0 11684 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_106
timestamp 1624635492
transform 1 0 10856 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1448
timestamp 1624635492
transform 1 0 11592 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_127
timestamp 1624635492
transform 1 0 12788 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_17
timestamp 1624635492
transform 1 0 2668 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_11
timestamp 1624635492
transform 1 0 2116 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_3
timestamp 1624635492
transform 1 0 1380 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output384_A
timestamp 1624635492
transform 1 0 2484 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output384
timestamp 1624635492
transform -1 0 2116 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1624635492
transform 1 0 1104 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_30
timestamp 1624635492
transform 1 0 3864 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1459
timestamp 1624635492
transform 1 0 3772 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_54
timestamp 1624635492
transform 1 0 6072 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_42
timestamp 1624635492
transform 1 0 4968 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_78
timestamp 1624635492
transform 1 0 8280 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_66
timestamp 1624635492
transform 1 0 7176 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_99
timestamp 1624635492
transform 1 0 10212 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_87
timestamp 1624635492
transform 1 0 9108 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1460
timestamp 1624635492
transform 1 0 9016 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_111
timestamp 1624635492
transform 1 0 11316 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_135
timestamp 1624635492
transform 1 0 13524 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_123
timestamp 1624635492
transform 1 0 12420 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_13
timestamp 1624635492
transform 1 0 2300 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_10
timestamp 1624635492
transform 1 0 2024 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_6
timestamp 1624635492
transform 1 0 1656 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output422_A
timestamp 1624635492
transform 1 0 2116 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1624635492
transform 1 0 1104 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _107_
timestamp 1624635492
transform 1 0 1380 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_117_37
timestamp 1624635492
transform 1 0 4508 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_25
timestamp 1624635492
transform 1 0 3404 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_58
timestamp 1624635492
transform 1 0 6440 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_49
timestamp 1624635492
transform 1 0 5612 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1472
timestamp 1624635492
transform 1 0 6348 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_70
timestamp 1624635492
transform 1 0 7544 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_94
timestamp 1624635492
transform 1 0 9752 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_82
timestamp 1624635492
transform 1 0 8648 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_115
timestamp 1624635492
transform 1 0 11684 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_106
timestamp 1624635492
transform 1 0 10856 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1473
timestamp 1624635492
transform 1 0 11592 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_127
timestamp 1624635492
transform 1 0 12788 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1624635492
transform 1 0 1104 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1624635492
transform 1 0 1104 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output383
timestamp 1624635492
transform -1 0 2116 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output422
timestamp 1624635492
transform -1 0 2116 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_3
timestamp 1624635492
transform 1 0 1380 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_3
timestamp 1624635492
transform 1 0 1380 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform -1 0 2760 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_11
timestamp 1624635492
transform 1 0 2116 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_119_11
timestamp 1624635492
transform 1 0 2116 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output421
timestamp 1624635492
transform -1 0 3220 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_18
timestamp 1624635492
transform 1 0 2760 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1484
timestamp 1624635492
transform 1 0 3772 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1497
timestamp 1624635492
transform 1 0 3772 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 3312 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_118_24
timestamp 1624635492
transform 1 0 3312 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_28
timestamp 1624635492
transform 1 0 3680 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_23
timestamp 1624635492
transform 1 0 3220 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output383_A
timestamp 1624635492
transform -1 0 4048 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output421_A
timestamp 1624635492
transform 1 0 3864 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_119_32
timestamp 1624635492
transform 1 0 4048 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_32
timestamp 1624635492
transform 1 0 4048 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_59
timestamp 1624635492
transform 1 0 6532 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_57
timestamp 1624635492
transform 1 0 6348 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_49
timestamp 1624635492
transform 1 0 5612 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_119_43
timestamp 1624635492
transform 1 0 5060 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_56
timestamp 1624635492
transform 1 0 6256 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_44
timestamp 1624635492
transform 1 0 5152 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 5612 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1624635492
transform -1 0 5060 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1498
timestamp 1624635492
transform 1 0 6440 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_71
timestamp 1624635492
transform 1 0 7636 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_68
timestamp 1624635492
transform 1 0 7360 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output382
timestamp 1624635492
transform 1 0 8372 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_90
timestamp 1624635492
transform 1 0 9384 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_83
timestamp 1624635492
transform 1 0 8740 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_99
timestamp 1624635492
transform 1 0 10212 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_87
timestamp 1624635492
transform 1 0 9108 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_80
timestamp 1624635492
transform 1 0 8464 0 -1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output382_A
timestamp 1624635492
transform -1 0 9384 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1499
timestamp 1624635492
transform 1 0 9108 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1485
timestamp 1624635492
transform 1 0 9016 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_117
timestamp 1624635492
transform 1 0 11868 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_115
timestamp 1624635492
transform 1 0 11684 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_107
timestamp 1624635492
transform 1 0 10948 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_102
timestamp 1624635492
transform 1 0 10488 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_109
timestamp 1624635492
transform 1 0 11132 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output420_A
timestamp 1624635492
transform 1 0 10948 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output420
timestamp 1624635492
transform -1 0 10948 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1500
timestamp 1624635492
transform 1 0 11776 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_133
timestamp 1624635492
transform 1 0 13340 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_127
timestamp 1624635492
transform 1 0 12788 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_123
timestamp 1624635492
transform 1 0 12420 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_133
timestamp 1624635492
transform 1 0 13340 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_121
timestamp 1624635492
transform 1 0 12236 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 13340 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform -1 0 12788 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_139
timestamp 1624635492
transform 1 0 13892 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_151
timestamp 1624635492
transform 1 0 14996 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_172
timestamp 1624635492
transform 1 0 16928 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_163
timestamp 1624635492
transform 1 0 16100 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1349
timestamp 1624635492
transform 1 0 16836 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_184
timestamp 1624635492
transform 1 0 18032 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_196
timestamp 1624635492
transform 1 0 19136 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_208
timestamp 1624635492
transform 1 0 20240 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_220
timestamp 1624635492
transform 1 0 21344 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_229
timestamp 1624635492
transform 1 0 22172 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1350
timestamp 1624635492
transform 1 0 22080 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_241
timestamp 1624635492
transform 1 0 23276 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_253
timestamp 1624635492
transform 1 0 24380 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_265
timestamp 1624635492
transform 1 0 25484 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_144
timestamp 1624635492
transform 1 0 14352 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1361
timestamp 1624635492
transform 1 0 14260 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_156
timestamp 1624635492
transform 1 0 15456 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_168
timestamp 1624635492
transform 1 0 16560 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_180
timestamp 1624635492
transform 1 0 17664 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_192
timestamp 1624635492
transform 1 0 18768 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1362
timestamp 1624635492
transform 1 0 19504 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_213
timestamp 1624635492
transform 1 0 20700 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_201
timestamp 1624635492
transform 1 0 19596 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_225
timestamp 1624635492
transform 1 0 21804 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_237
timestamp 1624635492
transform 1 0 22908 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_249
timestamp 1624635492
transform 1 0 24012 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_258
timestamp 1624635492
transform 1 0 24840 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1363
timestamp 1624635492
transform 1 0 24748 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_270
timestamp 1624635492
transform 1 0 25944 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_144
timestamp 1624635492
transform 1 0 14352 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_142
timestamp 1624635492
transform 1 0 14168 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_139
timestamp 1624635492
transform 1 0 13892 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1386
timestamp 1624635492
transform 1 0 14260 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_156
timestamp 1624635492
transform 1 0 15456 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_151
timestamp 1624635492
transform 1 0 14996 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_168
timestamp 1624635492
transform 1 0 16560 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_172
timestamp 1624635492
transform 1 0 16928 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_109_163
timestamp 1624635492
transform 1 0 16100 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1374
timestamp 1624635492
transform 1 0 16836 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_180
timestamp 1624635492
transform 1 0 17664 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_179
timestamp 1624635492
transform 1 0 17572 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _151_
timestamp 1624635492
transform 1 0 17296 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_110_192
timestamp 1624635492
transform 1 0 18768 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_191
timestamp 1624635492
transform 1 0 18676 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1387
timestamp 1624635492
transform 1 0 19504 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_211
timestamp 1624635492
transform 1 0 20516 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_207
timestamp 1624635492
transform 1 0 20148 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_110_201
timestamp 1624635492
transform 1 0 19596 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_109_203
timestamp 1624635492
transform 1 0 19780 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1624635492
transform 1 0 20240 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_217
timestamp 1624635492
transform 1 0 21068 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_215
timestamp 1624635492
transform 1 0 20884 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1624635492
transform 1 0 20884 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_110_229
timestamp 1624635492
transform 1 0 22172 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_229
timestamp 1624635492
transform 1 0 22172 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_227
timestamp 1624635492
transform 1 0 21988 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1375
timestamp 1624635492
transform 1 0 22080 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_241
timestamp 1624635492
transform 1 0 23276 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_241
timestamp 1624635492
transform 1 0 23276 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_258
timestamp 1624635492
transform 1 0 24840 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_253
timestamp 1624635492
transform 1 0 24380 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_253
timestamp 1624635492
transform 1 0 24380 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1388
timestamp 1624635492
transform 1 0 24748 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_270
timestamp 1624635492
transform 1 0 25944 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_265
timestamp 1624635492
transform 1 0 25484 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_139
timestamp 1624635492
transform 1 0 13892 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_151
timestamp 1624635492
transform 1 0 14996 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_172
timestamp 1624635492
transform 1 0 16928 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_163
timestamp 1624635492
transform 1 0 16100 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1399
timestamp 1624635492
transform 1 0 16836 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_184
timestamp 1624635492
transform 1 0 18032 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_196
timestamp 1624635492
transform 1 0 19136 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_208
timestamp 1624635492
transform 1 0 20240 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_220
timestamp 1624635492
transform 1 0 21344 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_229
timestamp 1624635492
transform 1 0 22172 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1400
timestamp 1624635492
transform 1 0 22080 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_241
timestamp 1624635492
transform 1 0 23276 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_253
timestamp 1624635492
transform 1 0 24380 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_265
timestamp 1624635492
transform 1 0 25484 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_144
timestamp 1624635492
transform 1 0 14352 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_112_141
timestamp 1624635492
transform 1 0 14076 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1411
timestamp 1624635492
transform 1 0 14260 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_156
timestamp 1624635492
transform 1 0 15456 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_168
timestamp 1624635492
transform 1 0 16560 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_180
timestamp 1624635492
transform 1 0 17664 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_192
timestamp 1624635492
transform 1 0 18768 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1412
timestamp 1624635492
transform 1 0 19504 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_213
timestamp 1624635492
transform 1 0 20700 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_201
timestamp 1624635492
transform 1 0 19596 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_225
timestamp 1624635492
transform 1 0 21804 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_237
timestamp 1624635492
transform 1 0 22908 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_249
timestamp 1624635492
transform 1 0 24012 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_258
timestamp 1624635492
transform 1 0 24840 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1413
timestamp 1624635492
transform 1 0 24748 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_270
timestamp 1624635492
transform 1 0 25944 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_144
timestamp 1624635492
transform 1 0 14352 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_144
timestamp 1624635492
transform 1 0 14352 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__D
timestamp 1624635492
transform 1 0 14720 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1436
timestamp 1624635492
transform 1 0 14260 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_156
timestamp 1624635492
transform 1 0 15456 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_156
timestamp 1624635492
transform 1 0 15456 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_150
timestamp 1624635492
transform 1 0 14904 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__CLK
timestamp 1624635492
transform 1 0 15272 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_168
timestamp 1624635492
transform 1 0 16560 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_172
timestamp 1624635492
transform 1 0 16928 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_113_168
timestamp 1624635492
transform 1 0 16560 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1424
timestamp 1624635492
transform 1 0 16836 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_180
timestamp 1624635492
transform 1 0 17664 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_184
timestamp 1624635492
transform 1 0 18032 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_192
timestamp 1624635492
transform 1 0 18768 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_196
timestamp 1624635492
transform 1 0 19136 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1437
timestamp 1624635492
transform 1 0 19504 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_213
timestamp 1624635492
transform 1 0 20700 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_201
timestamp 1624635492
transform 1 0 19596 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_208
timestamp 1624635492
transform 1 0 20240 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_225
timestamp 1624635492
transform 1 0 21804 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_220
timestamp 1624635492
transform 1 0 21344 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_237
timestamp 1624635492
transform 1 0 22908 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_229
timestamp 1624635492
transform 1 0 22172 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1425
timestamp 1624635492
transform 1 0 22080 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_249
timestamp 1624635492
transform 1 0 24012 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_241
timestamp 1624635492
transform 1 0 23276 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_258
timestamp 1624635492
transform 1 0 24840 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_253
timestamp 1624635492
transform 1 0 24380 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1438
timestamp 1624635492
transform 1 0 24748 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_270
timestamp 1624635492
transform 1 0 25944 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_265
timestamp 1624635492
transform 1 0 25484 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_139
timestamp 1624635492
transform 1 0 13892 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_151
timestamp 1624635492
transform 1 0 14996 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_172
timestamp 1624635492
transform 1 0 16928 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_115_163
timestamp 1624635492
transform 1 0 16100 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1449
timestamp 1624635492
transform 1 0 16836 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_179
timestamp 1624635492
transform 1 0 17572 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _328_
timestamp 1624635492
transform -1 0 17572 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_191
timestamp 1624635492
transform 1 0 18676 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_203
timestamp 1624635492
transform 1 0 19780 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_215
timestamp 1624635492
transform 1 0 20884 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_229
timestamp 1624635492
transform 1 0 22172 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_115_227
timestamp 1624635492
transform 1 0 21988 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1450
timestamp 1624635492
transform 1 0 22080 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_241
timestamp 1624635492
transform 1 0 23276 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_253
timestamp 1624635492
transform 1 0 24380 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_265
timestamp 1624635492
transform 1 0 25484 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_144
timestamp 1624635492
transform 1 0 14352 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1461
timestamp 1624635492
transform 1 0 14260 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_156
timestamp 1624635492
transform 1 0 15456 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_168
timestamp 1624635492
transform 1 0 16560 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_180
timestamp 1624635492
transform 1 0 17664 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_192
timestamp 1624635492
transform 1 0 18768 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1462
timestamp 1624635492
transform 1 0 19504 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_213
timestamp 1624635492
transform 1 0 20700 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_201
timestamp 1624635492
transform 1 0 19596 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_225
timestamp 1624635492
transform 1 0 21804 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_239
timestamp 1624635492
transform 1 0 23092 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_233
timestamp 1624635492
transform 1 0 22540 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _150_
timestamp 1624635492
transform 1 0 22816 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_116_251
timestamp 1624635492
transform 1 0 24196 0 -1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_116_258
timestamp 1624635492
transform 1 0 24840 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1463
timestamp 1624635492
transform 1 0 24748 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_270
timestamp 1624635492
transform 1 0 25944 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_144
timestamp 1624635492
transform 1 0 14352 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_118_141
timestamp 1624635492
transform 1 0 14076 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_117_147
timestamp 1624635492
transform 1 0 14628 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_117_139
timestamp 1624635492
transform 1 0 13892 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1486
timestamp 1624635492
transform 1 0 14260 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _329_
timestamp 1624635492
transform -1 0 15088 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_156
timestamp 1624635492
transform 1 0 15456 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_152
timestamp 1624635492
transform 1 0 15088 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_168
timestamp 1624635492
transform 1 0 16560 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_172
timestamp 1624635492
transform 1 0 16928 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_170
timestamp 1624635492
transform 1 0 16744 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_117_164
timestamp 1624635492
transform 1 0 16192 0 1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1474
timestamp 1624635492
transform 1 0 16836 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_180
timestamp 1624635492
transform 1 0 17664 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_184
timestamp 1624635492
transform 1 0 18032 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_192
timestamp 1624635492
transform 1 0 18768 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_196
timestamp 1624635492
transform 1 0 19136 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1487
timestamp 1624635492
transform 1 0 19504 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_213
timestamp 1624635492
transform 1 0 20700 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_201
timestamp 1624635492
transform 1 0 19596 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_208
timestamp 1624635492
transform 1 0 20240 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_225
timestamp 1624635492
transform 1 0 21804 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_220
timestamp 1624635492
transform 1 0 21344 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_237
timestamp 1624635492
transform 1 0 22908 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_229
timestamp 1624635492
transform 1 0 22172 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1475
timestamp 1624635492
transform 1 0 22080 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_249
timestamp 1624635492
transform 1 0 24012 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_241
timestamp 1624635492
transform 1 0 23276 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_258
timestamp 1624635492
transform 1 0 24840 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_253
timestamp 1624635492
transform 1 0 24380 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1488
timestamp 1624635492
transform 1 0 24748 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_270
timestamp 1624635492
transform 1 0 25944 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_265
timestamp 1624635492
transform 1 0 25484 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_146
timestamp 1624635492
transform 1 0 14536 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1501
timestamp 1624635492
transform 1 0 14444 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_158
timestamp 1624635492
transform 1 0 15640 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_119_170
timestamp 1624635492
transform 1 0 16744 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output381_A
timestamp 1624635492
transform -1 0 17388 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output381
timestamp 1624635492
transform -1 0 16744 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1502
timestamp 1624635492
transform 1 0 17112 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_119_185
timestamp 1624635492
transform 1 0 18124 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_119_177
timestamp 1624635492
transform 1 0 17388 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_119_198
timestamp 1624635492
transform 1 0 19320 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_192
timestamp 1624635492
transform 1 0 18768 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output419_A
timestamp 1624635492
transform -1 0 19320 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output419
timestamp 1624635492
transform -1 0 18768 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_212
timestamp 1624635492
transform 1 0 20608 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_208
timestamp 1624635492
transform 1 0 20240 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_204
timestamp 1624635492
transform 1 0 19872 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_202
timestamp 1624635492
transform 1 0 19688 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1624635492
transform -1 0 20608 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1503
timestamp 1624635492
transform 1 0 19780 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_218
timestamp 1624635492
transform 1 0 21160 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 21160 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_119_233
timestamp 1624635492
transform 1 0 22540 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_230
timestamp 1624635492
transform 1 0 22264 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1504
timestamp 1624635492
transform 1 0 22448 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_245
timestamp 1624635492
transform 1 0 23644 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output380
timestamp 1624635492
transform -1 0 24564 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_262
timestamp 1624635492
transform 1 0 25208 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_119_255
timestamp 1624635492
transform 1 0 24564 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1505
timestamp 1624635492
transform 1 0 25116 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_268
timestamp 1624635492
transform 1 0 25760 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output418_A
timestamp 1624635492
transform -1 0 25760 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output418
timestamp 1624635492
transform -1 0 26496 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_286
timestamp 1624635492
transform 1 0 27416 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_277
timestamp 1624635492
transform 1 0 26588 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1351
timestamp 1624635492
transform 1 0 27324 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_310
timestamp 1624635492
transform 1 0 29624 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_298
timestamp 1624635492
transform 1 0 28520 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_322
timestamp 1624635492
transform 1 0 30728 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_343
timestamp 1624635492
transform 1 0 32660 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_334
timestamp 1624635492
transform 1 0 31832 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1352
timestamp 1624635492
transform 1 0 32568 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_367
timestamp 1624635492
transform 1 0 34868 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_355
timestamp 1624635492
transform 1 0 33764 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_391
timestamp 1624635492
transform 1 0 37076 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_379
timestamp 1624635492
transform 1 0 35972 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_400
timestamp 1624635492
transform 1 0 37904 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1353
timestamp 1624635492
transform 1 0 37812 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_282
timestamp 1624635492
transform 1 0 27048 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_306
timestamp 1624635492
transform 1 0 29256 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_294
timestamp 1624635492
transform 1 0 28152 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_327
timestamp 1624635492
transform 1 0 31188 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_315
timestamp 1624635492
transform 1 0 30084 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1364
timestamp 1624635492
transform 1 0 29992 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_351
timestamp 1624635492
transform 1 0 33396 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_339
timestamp 1624635492
transform 1 0 32292 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_372
timestamp 1624635492
transform 1 0 35328 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_363
timestamp 1624635492
transform 1 0 34500 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1365
timestamp 1624635492
transform 1 0 35236 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_384
timestamp 1624635492
transform 1 0 36432 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_408
timestamp 1624635492
transform 1 0 38640 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_396
timestamp 1624635492
transform 1 0 37536 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_286
timestamp 1624635492
transform 1 0 27416 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_277
timestamp 1624635492
transform 1 0 26588 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1376
timestamp 1624635492
transform 1 0 27324 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_310
timestamp 1624635492
transform 1 0 29624 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_298
timestamp 1624635492
transform 1 0 28520 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_322
timestamp 1624635492
transform 1 0 30728 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_343
timestamp 1624635492
transform 1 0 32660 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_334
timestamp 1624635492
transform 1 0 31832 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1377
timestamp 1624635492
transform 1 0 32568 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_367
timestamp 1624635492
transform 1 0 34868 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_355
timestamp 1624635492
transform 1 0 33764 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_390
timestamp 1624635492
transform 1 0 36984 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_109_379
timestamp 1624635492
transform 1 0 35972 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _115_
timestamp 1624635492
transform 1 0 36708 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_400
timestamp 1624635492
transform 1 0 37904 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_398
timestamp 1624635492
transform 1 0 37720 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1378
timestamp 1624635492
transform 1 0 37812 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_282
timestamp 1624635492
transform 1 0 27048 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_306
timestamp 1624635492
transform 1 0 29256 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_294
timestamp 1624635492
transform 1 0 28152 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_327
timestamp 1624635492
transform 1 0 31188 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_315
timestamp 1624635492
transform 1 0 30084 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1389
timestamp 1624635492
transform 1 0 29992 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_351
timestamp 1624635492
transform 1 0 33396 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_339
timestamp 1624635492
transform 1 0 32292 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_372
timestamp 1624635492
transform 1 0 35328 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_363
timestamp 1624635492
transform 1 0 34500 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1390
timestamp 1624635492
transform 1 0 35236 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_384
timestamp 1624635492
transform 1 0 36432 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_408
timestamp 1624635492
transform 1 0 38640 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_396
timestamp 1624635492
transform 1 0 37536 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_282
timestamp 1624635492
transform 1 0 27048 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_286
timestamp 1624635492
transform 1 0 27416 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_277
timestamp 1624635492
transform 1 0 26588 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1401
timestamp 1624635492
transform 1 0 27324 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_306
timestamp 1624635492
transform 1 0 29256 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_294
timestamp 1624635492
transform 1 0 28152 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_310
timestamp 1624635492
transform 1 0 29624 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_298
timestamp 1624635492
transform 1 0 28520 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_327
timestamp 1624635492
transform 1 0 31188 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_315
timestamp 1624635492
transform 1 0 30084 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_322
timestamp 1624635492
transform 1 0 30728 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1414
timestamp 1624635492
transform 1 0 29992 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_351
timestamp 1624635492
transform 1 0 33396 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_339
timestamp 1624635492
transform 1 0 32292 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_343
timestamp 1624635492
transform 1 0 32660 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_334
timestamp 1624635492
transform 1 0 31832 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1402
timestamp 1624635492
transform 1 0 32568 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_372
timestamp 1624635492
transform 1 0 35328 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_363
timestamp 1624635492
transform 1 0 34500 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_367
timestamp 1624635492
transform 1 0 34868 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_355
timestamp 1624635492
transform 1 0 33764 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1415
timestamp 1624635492
transform 1 0 35236 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_384
timestamp 1624635492
transform 1 0 36432 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_391
timestamp 1624635492
transform 1 0 37076 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_387
timestamp 1624635492
transform 1 0 36708 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_379
timestamp 1624635492
transform 1 0 35972 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _162_
timestamp 1624635492
transform -1 0 37076 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_408
timestamp 1624635492
transform 1 0 38640 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_396
timestamp 1624635492
transform 1 0 37536 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_400
timestamp 1624635492
transform 1 0 37904 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1403
timestamp 1624635492
transform 1 0 37812 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_286
timestamp 1624635492
transform 1 0 27416 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_277
timestamp 1624635492
transform 1 0 26588 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1426
timestamp 1624635492
transform 1 0 27324 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_310
timestamp 1624635492
transform 1 0 29624 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_298
timestamp 1624635492
transform 1 0 28520 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_322
timestamp 1624635492
transform 1 0 30728 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_343
timestamp 1624635492
transform 1 0 32660 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_334
timestamp 1624635492
transform 1 0 31832 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1427
timestamp 1624635492
transform 1 0 32568 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_367
timestamp 1624635492
transform 1 0 34868 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_355
timestamp 1624635492
transform 1 0 33764 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_391
timestamp 1624635492
transform 1 0 37076 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_379
timestamp 1624635492
transform 1 0 35972 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_400
timestamp 1624635492
transform 1 0 37904 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1428
timestamp 1624635492
transform 1 0 37812 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_282
timestamp 1624635492
transform 1 0 27048 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_306
timestamp 1624635492
transform 1 0 29256 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_294
timestamp 1624635492
transform 1 0 28152 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_327
timestamp 1624635492
transform 1 0 31188 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_315
timestamp 1624635492
transform 1 0 30084 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1439
timestamp 1624635492
transform 1 0 29992 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_351
timestamp 1624635492
transform 1 0 33396 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_339
timestamp 1624635492
transform 1 0 32292 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_372
timestamp 1624635492
transform 1 0 35328 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_363
timestamp 1624635492
transform 1 0 34500 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1440
timestamp 1624635492
transform 1 0 35236 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_384
timestamp 1624635492
transform 1 0 36432 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_408
timestamp 1624635492
transform 1 0 38640 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_396
timestamp 1624635492
transform 1 0 37536 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_286
timestamp 1624635492
transform 1 0 27416 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_277
timestamp 1624635492
transform 1 0 26588 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1451
timestamp 1624635492
transform 1 0 27324 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_310
timestamp 1624635492
transform 1 0 29624 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_298
timestamp 1624635492
transform 1 0 28520 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_322
timestamp 1624635492
transform 1 0 30728 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_343
timestamp 1624635492
transform 1 0 32660 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_334
timestamp 1624635492
transform 1 0 31832 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1452
timestamp 1624635492
transform 1 0 32568 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_367
timestamp 1624635492
transform 1 0 34868 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_355
timestamp 1624635492
transform 1 0 33764 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_391
timestamp 1624635492
transform 1 0 37076 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_379
timestamp 1624635492
transform 1 0 35972 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_400
timestamp 1624635492
transform 1 0 37904 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1453
timestamp 1624635492
transform 1 0 37812 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_282
timestamp 1624635492
transform 1 0 27048 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_306
timestamp 1624635492
transform 1 0 29256 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_294
timestamp 1624635492
transform 1 0 28152 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_327
timestamp 1624635492
transform 1 0 31188 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_315
timestamp 1624635492
transform 1 0 30084 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1464
timestamp 1624635492
transform 1 0 29992 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_351
timestamp 1624635492
transform 1 0 33396 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_339
timestamp 1624635492
transform 1 0 32292 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_372
timestamp 1624635492
transform 1 0 35328 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_363
timestamp 1624635492
transform 1 0 34500 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1465
timestamp 1624635492
transform 1 0 35236 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_384
timestamp 1624635492
transform 1 0 36432 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_408
timestamp 1624635492
transform 1 0 38640 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_396
timestamp 1624635492
transform 1 0 37536 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_286
timestamp 1624635492
transform 1 0 27416 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_277
timestamp 1624635492
transform 1 0 26588 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1476
timestamp 1624635492
transform 1 0 27324 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_310
timestamp 1624635492
transform 1 0 29624 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_298
timestamp 1624635492
transform 1 0 28520 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_322
timestamp 1624635492
transform 1 0 30728 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_343
timestamp 1624635492
transform 1 0 32660 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_334
timestamp 1624635492
transform 1 0 31832 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1477
timestamp 1624635492
transform 1 0 32568 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_362
timestamp 1624635492
transform 1 0 34408 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_359
timestamp 1624635492
transform 1 0 34132 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_355
timestamp 1624635492
transform 1 0 33764 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__CLK
timestamp 1624635492
transform -1 0 34408 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _341_
timestamp 1624635492
transform -1 0 36524 0 1 65824
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_117_391
timestamp 1624635492
transform 1 0 37076 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_117_385
timestamp 1624635492
transform 1 0 36524 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__D
timestamp 1624635492
transform 1 0 36892 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_117_400
timestamp 1624635492
transform 1 0 37904 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1478
timestamp 1624635492
transform 1 0 37812 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_291
timestamp 1624635492
transform 1 0 27876 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_119_288
timestamp 1624635492
transform 1 0 27600 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_119_276
timestamp 1624635492
transform 1 0 26496 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_282
timestamp 1624635492
transform 1 0 27048 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1506
timestamp 1624635492
transform 1 0 27784 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_304
timestamp 1624635492
transform 1 0 29072 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_298
timestamp 1624635492
transform 1 0 28520 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_306
timestamp 1624635492
transform 1 0 29256 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_294
timestamp 1624635492
transform 1 0 28152 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 29072 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform -1 0 28520 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_332
timestamp 1624635492
transform 1 0 31648 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_320
timestamp 1624635492
transform 1 0 30544 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_316
timestamp 1624635492
transform 1 0 30176 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_322
timestamp 1624635492
transform 1 0 30728 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_315
timestamp 1624635492
transform 1 0 30084 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1507
timestamp 1624635492
transform 1 0 30452 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1489
timestamp 1624635492
transform 1 0 29992 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _178_
timestamp 1624635492
transform -1 0 30728 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_119_351
timestamp 1624635492
transform 1 0 33396 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_119_340
timestamp 1624635492
transform 1 0 32384 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_118_346
timestamp 1624635492
transform 1 0 32936 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_334
timestamp 1624635492
transform 1 0 31832 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output378_A
timestamp 1624635492
transform -1 0 33396 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output378
timestamp 1624635492
transform -1 0 32384 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1508
timestamp 1624635492
transform 1 0 33120 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_361
timestamp 1624635492
transform 1 0 34316 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_372
timestamp 1624635492
transform 1 0 35328 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_118_369
timestamp 1624635492
transform 1 0 35052 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_118_357
timestamp 1624635492
transform 1 0 33948 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_354
timestamp 1624635492
transform 1 0 33672 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output416_A
timestamp 1624635492
transform 1 0 33764 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output416
timestamp 1624635492
transform -1 0 34316 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1490
timestamp 1624635492
transform 1 0 35236 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_391
timestamp 1624635492
transform 1 0 37076 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_385
timestamp 1624635492
transform 1 0 36524 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_378
timestamp 1624635492
transform 1 0 35880 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_373
timestamp 1624635492
transform 1 0 35420 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_384
timestamp 1624635492
transform 1 0 36432 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 37076 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform -1 0 36524 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1509
timestamp 1624635492
transform 1 0 35788 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_407
timestamp 1624635492
transform 1 0 38548 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_119_403
timestamp 1624635492
transform 1 0 38180 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_408
timestamp 1624635492
transform 1 0 38640 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_396
timestamp 1624635492
transform 1 0 37536 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1510
timestamp 1624635492
transform 1 0 38456 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_424
timestamp 1624635492
transform 1 0 40112 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_412
timestamp 1624635492
transform 1 0 39008 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_448
timestamp 1624635492
transform 1 0 42320 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_436
timestamp 1624635492
transform 1 0 41216 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_469
timestamp 1624635492
transform 1 0 44252 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_457
timestamp 1624635492
transform 1 0 43148 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1354
timestamp 1624635492
transform 1 0 43056 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_493
timestamp 1624635492
transform 1 0 46460 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_481
timestamp 1624635492
transform 1 0 45356 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_514
timestamp 1624635492
transform 1 0 48392 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_505
timestamp 1624635492
transform 1 0 47564 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1355
timestamp 1624635492
transform 1 0 48300 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_538
timestamp 1624635492
transform 1 0 50600 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_526
timestamp 1624635492
transform 1 0 49496 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_546
timestamp 1624635492
transform 1 0 51336 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_429
timestamp 1624635492
transform 1 0 40572 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_420
timestamp 1624635492
transform 1 0 39744 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1366
timestamp 1624635492
transform 1 0 40480 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_453
timestamp 1624635492
transform 1 0 42780 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_441
timestamp 1624635492
transform 1 0 41676 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_465
timestamp 1624635492
transform 1 0 43884 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_486
timestamp 1624635492
transform 1 0 45816 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_477
timestamp 1624635492
transform 1 0 44988 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1367
timestamp 1624635492
transform 1 0 45724 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_510
timestamp 1624635492
transform 1 0 48024 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_498
timestamp 1624635492
transform 1 0 46920 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_534
timestamp 1624635492
transform 1 0 50232 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_522
timestamp 1624635492
transform 1 0 49128 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_543
timestamp 1624635492
transform 1 0 51060 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1368
timestamp 1624635492
transform 1 0 50968 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_424
timestamp 1624635492
transform 1 0 40112 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_412
timestamp 1624635492
transform 1 0 39008 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_448
timestamp 1624635492
transform 1 0 42320 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_436
timestamp 1624635492
transform 1 0 41216 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_469
timestamp 1624635492
transform 1 0 44252 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_457
timestamp 1624635492
transform 1 0 43148 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1379
timestamp 1624635492
transform 1 0 43056 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_493
timestamp 1624635492
transform 1 0 46460 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_481
timestamp 1624635492
transform 1 0 45356 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_514
timestamp 1624635492
transform 1 0 48392 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_505
timestamp 1624635492
transform 1 0 47564 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1380
timestamp 1624635492
transform 1 0 48300 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_538
timestamp 1624635492
transform 1 0 50600 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_526
timestamp 1624635492
transform 1 0 49496 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_429
timestamp 1624635492
transform 1 0 40572 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_420
timestamp 1624635492
transform 1 0 39744 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1391
timestamp 1624635492
transform 1 0 40480 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_453
timestamp 1624635492
transform 1 0 42780 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_441
timestamp 1624635492
transform 1 0 41676 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_465
timestamp 1624635492
transform 1 0 43884 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_486
timestamp 1624635492
transform 1 0 45816 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_477
timestamp 1624635492
transform 1 0 44988 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1392
timestamp 1624635492
transform 1 0 45724 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_110_518
timestamp 1624635492
transform 1 0 48760 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_110_510
timestamp 1624635492
transform 1 0 48024 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_498
timestamp 1624635492
transform 1 0 46920 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_534
timestamp 1624635492
transform 1 0 50232 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_522
timestamp 1624635492
transform 1 0 49128 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__CLK
timestamp 1624635492
transform 1 0 48944 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_110_543
timestamp 1624635492
transform 1 0 51060 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1393
timestamp 1624635492
transform 1 0 50968 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_429
timestamp 1624635492
transform 1 0 40572 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_420
timestamp 1624635492
transform 1 0 39744 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_424
timestamp 1624635492
transform 1 0 40112 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_412
timestamp 1624635492
transform 1 0 39008 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1416
timestamp 1624635492
transform 1 0 40480 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_453
timestamp 1624635492
transform 1 0 42780 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_441
timestamp 1624635492
transform 1 0 41676 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_448
timestamp 1624635492
transform 1 0 42320 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_436
timestamp 1624635492
transform 1 0 41216 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_465
timestamp 1624635492
transform 1 0 43884 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_469
timestamp 1624635492
transform 1 0 44252 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_457
timestamp 1624635492
transform 1 0 43148 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1404
timestamp 1624635492
transform 1 0 43056 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_486
timestamp 1624635492
transform 1 0 45816 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_477
timestamp 1624635492
transform 1 0 44988 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_111_493
timestamp 1624635492
transform 1 0 46460 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_481
timestamp 1624635492
transform 1 0 45356 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1417
timestamp 1624635492
transform 1 0 45724 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_510
timestamp 1624635492
transform 1 0 48024 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_498
timestamp 1624635492
transform 1 0 46920 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_514
timestamp 1624635492
transform 1 0 48392 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_512
timestamp 1624635492
transform 1 0 48208 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_504
timestamp 1624635492
transform 1 0 47472 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__RESET_B
timestamp 1624635492
transform -1 0 48944 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__D
timestamp 1624635492
transform 1 0 48760 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1405
timestamp 1624635492
transform 1 0 48300 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _244_
timestamp 1624635492
transform 1 0 47196 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_112_540
timestamp 1624635492
transform 1 0 50784 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_112_532
timestamp 1624635492
transform 1 0 50048 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_520
timestamp 1624635492
transform 1 0 48944 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_520
timestamp 1624635492
transform 1 0 48944 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _334_
timestamp 1624635492
transform 1 0 49312 0 1 62560
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_112_543
timestamp 1624635492
transform 1 0 51060 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_545
timestamp 1624635492
transform 1 0 51244 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1418
timestamp 1624635492
transform 1 0 50968 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_424
timestamp 1624635492
transform 1 0 40112 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_412
timestamp 1624635492
transform 1 0 39008 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_448
timestamp 1624635492
transform 1 0 42320 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_436
timestamp 1624635492
transform 1 0 41216 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_469
timestamp 1624635492
transform 1 0 44252 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_457
timestamp 1624635492
transform 1 0 43148 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1429
timestamp 1624635492
transform 1 0 43056 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_493
timestamp 1624635492
transform 1 0 46460 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_481
timestamp 1624635492
transform 1 0 45356 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_514
timestamp 1624635492
transform 1 0 48392 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_505
timestamp 1624635492
transform 1 0 47564 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1430
timestamp 1624635492
transform 1 0 48300 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_538
timestamp 1624635492
transform 1 0 50600 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_526
timestamp 1624635492
transform 1 0 49496 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_429
timestamp 1624635492
transform 1 0 40572 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_420
timestamp 1624635492
transform 1 0 39744 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1441
timestamp 1624635492
transform 1 0 40480 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_453
timestamp 1624635492
transform 1 0 42780 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_441
timestamp 1624635492
transform 1 0 41676 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_465
timestamp 1624635492
transform 1 0 43884 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_486
timestamp 1624635492
transform 1 0 45816 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_477
timestamp 1624635492
transform 1 0 44988 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1442
timestamp 1624635492
transform 1 0 45724 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_510
timestamp 1624635492
transform 1 0 48024 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_498
timestamp 1624635492
transform 1 0 46920 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_534
timestamp 1624635492
transform 1 0 50232 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_522
timestamp 1624635492
transform 1 0 49128 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_543
timestamp 1624635492
transform 1 0 51060 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1443
timestamp 1624635492
transform 1 0 50968 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_424
timestamp 1624635492
transform 1 0 40112 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_412
timestamp 1624635492
transform 1 0 39008 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_450
timestamp 1624635492
transform 1 0 42504 0 1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_115_438
timestamp 1624635492
transform 1 0 41400 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_432
timestamp 1624635492
transform 1 0 40848 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _260_
timestamp 1624635492
transform 1 0 41124 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_469
timestamp 1624635492
transform 1 0 44252 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_457
timestamp 1624635492
transform 1 0 43148 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1454
timestamp 1624635492
transform 1 0 43056 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_493
timestamp 1624635492
transform 1 0 46460 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_481
timestamp 1624635492
transform 1 0 45356 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_514
timestamp 1624635492
transform 1 0 48392 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_505
timestamp 1624635492
transform 1 0 47564 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1455
timestamp 1624635492
transform 1 0 48300 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_538
timestamp 1624635492
transform 1 0 50600 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_526
timestamp 1624635492
transform 1 0 49496 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_429
timestamp 1624635492
transform 1 0 40572 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_420
timestamp 1624635492
transform 1 0 39744 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1466
timestamp 1624635492
transform 1 0 40480 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_453
timestamp 1624635492
transform 1 0 42780 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_441
timestamp 1624635492
transform 1 0 41676 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_465
timestamp 1624635492
transform 1 0 43884 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _160_
timestamp 1624635492
transform -1 0 44896 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_486
timestamp 1624635492
transform 1 0 45816 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_484
timestamp 1624635492
transform 1 0 45632 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_476
timestamp 1624635492
transform 1 0 44896 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1467
timestamp 1624635492
transform 1 0 45724 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_518
timestamp 1624635492
transform 1 0 48760 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_514
timestamp 1624635492
transform 1 0 48392 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_510
timestamp 1624635492
transform 1 0 48024 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_498
timestamp 1624635492
transform 1 0 46920 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _271_
timestamp 1624635492
transform 1 0 48484 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_530
timestamp 1624635492
transform 1 0 49864 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_543
timestamp 1624635492
transform 1 0 51060 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1468
timestamp 1624635492
transform 1 0 50968 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_424
timestamp 1624635492
transform 1 0 40112 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_412
timestamp 1624635492
transform 1 0 39008 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_448
timestamp 1624635492
transform 1 0 42320 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_436
timestamp 1624635492
transform 1 0 41216 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_469
timestamp 1624635492
transform 1 0 44252 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_457
timestamp 1624635492
transform 1 0 43148 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1479
timestamp 1624635492
transform 1 0 43056 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_493
timestamp 1624635492
transform 1 0 46460 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_481
timestamp 1624635492
transform 1 0 45356 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_514
timestamp 1624635492
transform 1 0 48392 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_505
timestamp 1624635492
transform 1 0 47564 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1480
timestamp 1624635492
transform 1 0 48300 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_538
timestamp 1624635492
transform 1 0 50600 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_526
timestamp 1624635492
transform 1 0 49496 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_424
timestamp 1624635492
transform 1 0 40112 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_119_416
timestamp 1624635492
transform 1 0 39376 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_413
timestamp 1624635492
transform 1 0 39100 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_429
timestamp 1624635492
transform 1 0 40572 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_118_420
timestamp 1624635492
transform 1 0 39744 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output377_A
timestamp 1624635492
transform -1 0 39376 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output377
timestamp 1624635492
transform -1 0 40112 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1491
timestamp 1624635492
transform 1 0 40480 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1511
timestamp 1624635492
transform 1 0 41124 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output415
timestamp 1624635492
transform -1 0 42044 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output415_A
timestamp 1624635492
transform 1 0 41492 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_118_437
timestamp 1624635492
transform 1 0 41308 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_119_432
timestamp 1624635492
transform 1 0 40848 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_436
timestamp 1624635492
transform 1 0 41216 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_440
timestamp 1624635492
transform 1 0 41584 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_441
timestamp 1624635492
transform 1 0 41676 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_453
timestamp 1624635492
transform 1 0 42780 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_445
timestamp 1624635492
transform 1 0 42044 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_472
timestamp 1624635492
transform 1 0 44528 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_465
timestamp 1624635492
transform 1 0 43884 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_463
timestamp 1624635492
transform 1 0 43700 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_457
timestamp 1624635492
transform 1 0 43148 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_118_465
timestamp 1624635492
transform 1 0 43884 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1624635492
transform -1 0 44528 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1512
timestamp 1624635492
transform 1 0 43792 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_494
timestamp 1624635492
transform 1 0 46552 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_490
timestamp 1624635492
transform 1 0 46184 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_478
timestamp 1624635492
transform 1 0 45080 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_486
timestamp 1624635492
transform 1 0 45816 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_477
timestamp 1624635492
transform 1 0 44988 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 45080 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1513
timestamp 1624635492
transform 1 0 46460 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1492
timestamp 1624635492
transform 1 0 45724 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_509
timestamp 1624635492
transform 1 0 47932 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_502
timestamp 1624635492
transform 1 0 47288 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_510
timestamp 1624635492
transform 1 0 48024 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_498
timestamp 1624635492
transform 1 0 46920 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output376
timestamp 1624635492
transform -1 0 47932 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_537
timestamp 1624635492
transform 1 0 50508 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_531
timestamp 1624635492
transform 1 0 49956 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_523
timestamp 1624635492
transform 1 0 49220 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_521
timestamp 1624635492
transform 1 0 49036 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_534
timestamp 1624635492
transform 1 0 50232 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_522
timestamp 1624635492
transform 1 0 49128 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output414_A
timestamp 1624635492
transform -1 0 50508 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output414
timestamp 1624635492
transform -1 0 49956 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1514
timestamp 1624635492
transform 1 0 49128 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_543
timestamp 1624635492
transform 1 0 51060 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1493
timestamp 1624635492
transform 1 0 50968 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_549
timestamp 1624635492
transform 1 0 51612 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__B2
timestamp 1624635492
transform 1 0 51428 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_571
timestamp 1624635492
transform 1 0 53636 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_569
timestamp 1624635492
transform 1 0 53452 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_561
timestamp 1624635492
transform 1 0 52716 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1356
timestamp 1624635492
transform 1 0 53544 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_583
timestamp 1624635492
transform 1 0 54740 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_595
timestamp 1624635492
transform 1 0 55844 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_607
timestamp 1624635492
transform 1 0 56948 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_619
timestamp 1624635492
transform 1 0 58052 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_628
timestamp 1624635492
transform 1 0 58880 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1357
timestamp 1624635492
transform 1 0 58788 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_640
timestamp 1624635492
transform 1 0 59984 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_652
timestamp 1624635492
transform 1 0 61088 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_664
timestamp 1624635492
transform 1 0 62192 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_676
timestamp 1624635492
transform 1 0 63296 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_550
timestamp 1624635492
transform 1 0 51704 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_555
timestamp 1624635492
transform 1 0 52164 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_571
timestamp 1624635492
transform 1 0 53636 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_562
timestamp 1624635492
transform 1 0 52808 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_567
timestamp 1624635492
transform 1 0 53268 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1381
timestamp 1624635492
transform 1 0 53544 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_583
timestamp 1624635492
transform 1 0 54740 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_579
timestamp 1624635492
transform 1 0 54372 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_595
timestamp 1624635492
transform 1 0 55844 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_591
timestamp 1624635492
transform 1 0 55476 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_607
timestamp 1624635492
transform 1 0 56948 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_600
timestamp 1624635492
transform 1 0 56304 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1369
timestamp 1624635492
transform 1 0 56212 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_619
timestamp 1624635492
transform 1 0 58052 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_612
timestamp 1624635492
transform 1 0 57408 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_628
timestamp 1624635492
transform 1 0 58880 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_636
timestamp 1624635492
transform 1 0 59616 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_624
timestamp 1624635492
transform 1 0 58512 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1382
timestamp 1624635492
transform 1 0 58788 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_640
timestamp 1624635492
transform 1 0 59984 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_648
timestamp 1624635492
transform 1 0 60720 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_652
timestamp 1624635492
transform 1 0 61088 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_657
timestamp 1624635492
transform 1 0 61548 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1370
timestamp 1624635492
transform 1 0 61456 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_664
timestamp 1624635492
transform 1 0 62192 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_669
timestamp 1624635492
transform 1 0 62652 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_676
timestamp 1624635492
transform 1 0 63296 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_681
timestamp 1624635492
transform 1 0 63756 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_555
timestamp 1624635492
transform 1 0 52164 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_567
timestamp 1624635492
transform 1 0 53268 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_579
timestamp 1624635492
transform 1 0 54372 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_591
timestamp 1624635492
transform 1 0 55476 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_600
timestamp 1624635492
transform 1 0 56304 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1394
timestamp 1624635492
transform 1 0 56212 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_612
timestamp 1624635492
transform 1 0 57408 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_636
timestamp 1624635492
transform 1 0 59616 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_624
timestamp 1624635492
transform 1 0 58512 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_648
timestamp 1624635492
transform 1 0 60720 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_657
timestamp 1624635492
transform 1 0 61548 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1395
timestamp 1624635492
transform 1 0 61456 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_669
timestamp 1624635492
transform 1 0 62652 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_681
timestamp 1624635492
transform 1 0 63756 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_555
timestamp 1624635492
transform 1 0 52164 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_557
timestamp 1624635492
transform 1 0 52348 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_567
timestamp 1624635492
transform 1 0 53268 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_571
timestamp 1624635492
transform 1 0 53636 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_569
timestamp 1624635492
transform 1 0 53452 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1406
timestamp 1624635492
transform 1 0 53544 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_579
timestamp 1624635492
transform 1 0 54372 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_583
timestamp 1624635492
transform 1 0 54740 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_591
timestamp 1624635492
transform 1 0 55476 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_595
timestamp 1624635492
transform 1 0 55844 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_600
timestamp 1624635492
transform 1 0 56304 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_607
timestamp 1624635492
transform 1 0 56948 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1419
timestamp 1624635492
transform 1 0 56212 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_612
timestamp 1624635492
transform 1 0 57408 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_619
timestamp 1624635492
transform 1 0 58052 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_636
timestamp 1624635492
transform 1 0 59616 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_624
timestamp 1624635492
transform 1 0 58512 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_628
timestamp 1624635492
transform 1 0 58880 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1407
timestamp 1624635492
transform 1 0 58788 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_648
timestamp 1624635492
transform 1 0 60720 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_640
timestamp 1624635492
transform 1 0 59984 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_657
timestamp 1624635492
transform 1 0 61548 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_652
timestamp 1624635492
transform 1 0 61088 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1420
timestamp 1624635492
transform 1 0 61456 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_669
timestamp 1624635492
transform 1 0 62652 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_664
timestamp 1624635492
transform 1 0 62192 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_681
timestamp 1624635492
transform 1 0 63756 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_676
timestamp 1624635492
transform 1 0 63296 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_550
timestamp 1624635492
transform 1 0 51704 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_571
timestamp 1624635492
transform 1 0 53636 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_562
timestamp 1624635492
transform 1 0 52808 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1431
timestamp 1624635492
transform 1 0 53544 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_583
timestamp 1624635492
transform 1 0 54740 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_595
timestamp 1624635492
transform 1 0 55844 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_607
timestamp 1624635492
transform 1 0 56948 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_619
timestamp 1624635492
transform 1 0 58052 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_628
timestamp 1624635492
transform 1 0 58880 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1432
timestamp 1624635492
transform 1 0 58788 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_640
timestamp 1624635492
transform 1 0 59984 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_652
timestamp 1624635492
transform 1 0 61088 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_664
timestamp 1624635492
transform 1 0 62192 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_676
timestamp 1624635492
transform 1 0 63296 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_550
timestamp 1624635492
transform 1 0 51704 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_114_555
timestamp 1624635492
transform 1 0 52164 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _305_
timestamp 1624635492
transform -1 0 52716 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_571
timestamp 1624635492
transform 1 0 53636 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_562
timestamp 1624635492
transform 1 0 52808 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_561
timestamp 1624635492
transform 1 0 52716 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1456
timestamp 1624635492
transform 1 0 53544 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_583
timestamp 1624635492
transform 1 0 54740 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_573
timestamp 1624635492
transform 1 0 53820 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_595
timestamp 1624635492
transform 1 0 55844 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_114_597
timestamp 1624635492
transform 1 0 56028 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_585
timestamp 1624635492
transform 1 0 54924 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_607
timestamp 1624635492
transform 1 0 56948 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_600
timestamp 1624635492
transform 1 0 56304 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1444
timestamp 1624635492
transform 1 0 56212 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_619
timestamp 1624635492
transform 1 0 58052 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_612
timestamp 1624635492
transform 1 0 57408 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_628
timestamp 1624635492
transform 1 0 58880 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_636
timestamp 1624635492
transform 1 0 59616 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_624
timestamp 1624635492
transform 1 0 58512 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1457
timestamp 1624635492
transform 1 0 58788 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_640
timestamp 1624635492
transform 1 0 59984 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_648
timestamp 1624635492
transform 1 0 60720 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_652
timestamp 1624635492
transform 1 0 61088 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_657
timestamp 1624635492
transform 1 0 61548 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1445
timestamp 1624635492
transform 1 0 61456 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_664
timestamp 1624635492
transform 1 0 62192 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_669
timestamp 1624635492
transform 1 0 62652 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_676
timestamp 1624635492
transform 1 0 63296 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_681
timestamp 1624635492
transform 1 0 63756 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_555
timestamp 1624635492
transform 1 0 52164 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_567
timestamp 1624635492
transform 1 0 53268 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_579
timestamp 1624635492
transform 1 0 54372 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_591
timestamp 1624635492
transform 1 0 55476 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_600
timestamp 1624635492
transform 1 0 56304 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1469
timestamp 1624635492
transform 1 0 56212 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_612
timestamp 1624635492
transform 1 0 57408 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_636
timestamp 1624635492
transform 1 0 59616 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_624
timestamp 1624635492
transform 1 0 58512 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_648
timestamp 1624635492
transform 1 0 60720 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_657
timestamp 1624635492
transform 1 0 61548 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1470
timestamp 1624635492
transform 1 0 61456 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_669
timestamp 1624635492
transform 1 0 62652 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_681
timestamp 1624635492
transform 1 0 63756 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_555
timestamp 1624635492
transform 1 0 52164 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_550
timestamp 1624635492
transform 1 0 51704 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_567
timestamp 1624635492
transform 1 0 53268 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_571
timestamp 1624635492
transform 1 0 53636 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_562
timestamp 1624635492
transform 1 0 52808 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1481
timestamp 1624635492
transform 1 0 53544 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_579
timestamp 1624635492
transform 1 0 54372 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_583
timestamp 1624635492
transform 1 0 54740 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_591
timestamp 1624635492
transform 1 0 55476 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_595
timestamp 1624635492
transform 1 0 55844 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_600
timestamp 1624635492
transform 1 0 56304 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_607
timestamp 1624635492
transform 1 0 56948 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1494
timestamp 1624635492
transform 1 0 56212 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_614
timestamp 1624635492
transform 1 0 57592 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_619
timestamp 1624635492
transform 1 0 58052 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output413_A
timestamp 1624635492
transform 1 0 57408 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_118_626
timestamp 1624635492
transform 1 0 58696 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_628
timestamp 1624635492
transform 1 0 58880 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1482
timestamp 1624635492
transform 1 0 58788 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_638
timestamp 1624635492
transform 1 0 59800 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_640
timestamp 1624635492
transform 1 0 59984 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_657
timestamp 1624635492
transform 1 0 61548 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_650
timestamp 1624635492
transform 1 0 60904 0 -1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_117_652
timestamp 1624635492
transform 1 0 61088 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1495
timestamp 1624635492
transform 1 0 61456 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_669
timestamp 1624635492
transform 1 0 62652 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_664
timestamp 1624635492
transform 1 0 62192 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_681
timestamp 1624635492
transform 1 0 63756 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_676
timestamp 1624635492
transform 1 0 63296 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_119_559
timestamp 1624635492
transform 1 0 52532 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_552
timestamp 1624635492
transform 1 0 51888 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_119_549
timestamp 1624635492
transform 1 0 51612 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1624635492
transform -1 0 52532 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1515
timestamp 1624635492
transform 1 0 51796 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_565
timestamp 1624635492
transform 1 0 53084 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 53084 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_119_581
timestamp 1624635492
transform 1 0 54556 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_119_577
timestamp 1624635492
transform 1 0 54188 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output375_A
timestamp 1624635492
transform -1 0 54924 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1516
timestamp 1624635492
transform 1 0 54464 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_593
timestamp 1624635492
transform 1 0 55660 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_585
timestamp 1624635492
transform 1 0 54924 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output375
timestamp 1624635492
transform -1 0 55660 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_610
timestamp 1624635492
transform 1 0 57224 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_605
timestamp 1624635492
transform 1 0 56764 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1517
timestamp 1624635492
transform 1 0 57132 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_618
timestamp 1624635492
transform 1 0 57960 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output413
timestamp 1624635492
transform -1 0 57960 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_634
timestamp 1624635492
transform 1 0 59432 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_630
timestamp 1624635492
transform 1 0 59064 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1624635492
transform -1 0 59432 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_641
timestamp 1624635492
transform 1 0 60076 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 60076 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1518
timestamp 1624635492
transform 1 0 59800 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_653
timestamp 1624635492
transform 1 0 61180 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_670
timestamp 1624635492
transform 1 0 62744 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_119_665
timestamp 1624635492
transform 1 0 62284 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output374_A
timestamp 1624635492
transform -1 0 62744 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output374
timestamp 1624635492
transform -1 0 63480 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1519
timestamp 1624635492
transform 1 0 62468 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_678
timestamp 1624635492
transform 1 0 63480 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_693
timestamp 1624635492
transform 1 0 64860 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_697
timestamp 1624635492
transform 1 0 65228 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_685
timestamp 1624635492
transform 1 0 64124 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1358
timestamp 1624635492
transform 1 0 64032 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_705
timestamp 1624635492
transform 1 0 65964 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_709
timestamp 1624635492
transform 1 0 66332 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_722
timestamp 1624635492
transform 1 0 67528 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_108_714
timestamp 1624635492
transform 1 0 66792 0 -1 61472
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_107_721
timestamp 1624635492
transform 1 0 67436 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 67528 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1624635492
transform -1 0 68172 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1371
timestamp 1624635492
transform 1 0 66700 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_729
timestamp 1624635492
transform 1 0 68172 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1624635492
transform -1 0 68816 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1624635492
transform -1 0 68816 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_693
timestamp 1624635492
transform 1 0 64860 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_697
timestamp 1624635492
transform 1 0 65228 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_685
timestamp 1624635492
transform 1 0 64124 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1383
timestamp 1624635492
transform 1 0 64032 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_705
timestamp 1624635492
transform 1 0 65964 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_709
timestamp 1624635492
transform 1 0 66332 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_716
timestamp 1624635492
transform 1 0 66976 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_721
timestamp 1624635492
transform 1 0 67436 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1624635492
transform 1 0 66792 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1396
timestamp 1624635492
transform 1 0 66700 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_110_732
timestamp 1624635492
transform 1 0 68448 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_728
timestamp 1624635492
transform 1 0 68080 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1624635492
transform -1 0 68816 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1624635492
transform -1 0 68816 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_693
timestamp 1624635492
transform 1 0 64860 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_697
timestamp 1624635492
transform 1 0 65228 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_685
timestamp 1624635492
transform 1 0 64124 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1408
timestamp 1624635492
transform 1 0 64032 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_705
timestamp 1624635492
transform 1 0 65964 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_111_709
timestamp 1624635492
transform 1 0 66332 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__B
timestamp 1624635492
transform -1 0 66700 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_112_721
timestamp 1624635492
transform 1 0 67436 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_718
timestamp 1624635492
transform 1 0 67160 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_112_714
timestamp 1624635492
transform 1 0 66792 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_111_724
timestamp 1624635492
transform 1 0 67712 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_111_713
timestamp 1624635492
transform 1 0 66700 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output410_A
timestamp 1624635492
transform 1 0 67252 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output410
timestamp 1624635492
transform 1 0 67804 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1421
timestamp 1624635492
transform 1 0 66700 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 67068 0 1 62560
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_112_729
timestamp 1624635492
transform 1 0 68172 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_732
timestamp 1624635492
transform 1 0 68448 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1624635492
transform -1 0 68816 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1624635492
transform -1 0 68816 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_115_697
timestamp 1624635492
transform 1 0 65228 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_685
timestamp 1624635492
transform 1 0 64124 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_693
timestamp 1624635492
transform 1 0 64860 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_697
timestamp 1624635492
transform 1 0 65228 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_685
timestamp 1624635492
transform 1 0 64124 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1458
timestamp 1624635492
transform 1 0 64032 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1433
timestamp 1624635492
transform 1 0 64032 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_710
timestamp 1624635492
transform 1 0 66424 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_115_705
timestamp 1624635492
transform 1 0 65964 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_114_705
timestamp 1624635492
transform 1 0 65964 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_113_709
timestamp 1624635492
transform 1 0 66332 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B1
timestamp 1624635492
transform -1 0 66424 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1446
timestamp 1624635492
transform 1 0 66700 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A1
timestamp 1624635492
transform -1 0 66976 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A2
timestamp 1624635492
transform 1 0 66976 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output372_A
timestamp 1624635492
transform -1 0 67436 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_113_717
timestamp 1624635492
transform 1 0 67068 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_114_714
timestamp 1624635492
transform 1 0 66792 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_115_716
timestamp 1624635492
transform 1 0 66976 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output372
timestamp 1624635492
transform 1 0 67804 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_721
timestamp 1624635492
transform 1 0 67436 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_115_727
timestamp 1624635492
transform 1 0 67988 0 1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _083_
timestamp 1624635492
transform -1 0 67988 0 1 64736
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_114_718
timestamp 1624635492
transform 1 0 67160 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_114_730
timestamp 1624635492
transform 1 0 68264 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_113_729
timestamp 1624635492
transform 1 0 68172 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1624635492
transform -1 0 68816 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1624635492
transform -1 0 68816 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1624635492
transform -1 0 68816 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_693
timestamp 1624635492
transform 1 0 64860 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_117_685
timestamp 1624635492
transform 1 0 64124 0 1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1624635492
transform 1 0 64860 0 -1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__A1
timestamp 1624635492
transform -1 0 64860 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__A2
timestamp 1624635492
transform -1 0 65412 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1483
timestamp 1624635492
transform 1 0 64032 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_699
timestamp 1624635492
transform 1 0 65412 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_701
timestamp 1624635492
transform 1 0 65596 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__B2
timestamp 1624635492
transform 1 0 65412 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_4  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 67068 0 1 65824
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_117_725
timestamp 1624635492
transform 1 0 67804 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_717
timestamp 1624635492
transform 1 0 67068 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_116_724
timestamp 1624635492
transform 1 0 67712 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_116_716
timestamp 1624635492
transform 1 0 66976 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A3
timestamp 1624635492
transform -1 0 66976 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 68172 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1624635492
transform -1 0 68172 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1471
timestamp 1624635492
transform 1 0 66700 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_729
timestamp 1624635492
transform 1 0 68172 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_729
timestamp 1624635492
transform 1 0 68172 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1624635492
transform -1 0 68816 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1624635492
transform -1 0 68816 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_697
timestamp 1624635492
transform 1 0 65228 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_692
timestamp 1624635492
transform 1 0 64768 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_693
timestamp 1624635492
transform 1 0 64860 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output412_A
timestamp 1624635492
transform -1 0 64768 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__B1
timestamp 1624635492
transform -1 0 65412 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1520
timestamp 1624635492
transform 1 0 65136 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_119_709
timestamp 1624635492
transform 1 0 66332 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_705
timestamp 1624635492
transform 1 0 65964 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_709
timestamp 1624635492
transform 1 0 66332 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_699
timestamp 1624635492
transform 1 0 65412 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output411_A
timestamp 1624635492
transform 1 0 66148 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output412
timestamp 1624635492
transform -1 0 65964 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform -1 0 66700 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1496
timestamp 1624635492
transform 1 0 66700 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output373
timestamp 1624635492
transform 1 0 67068 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 66976 0 -1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_119_713
timestamp 1624635492
transform 1 0 66700 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1521
timestamp 1624635492
transform 1 0 67804 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output411
timestamp 1624635492
transform 1 0 67804 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output373_A
timestamp 1624635492
transform -1 0 68080 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_118_724
timestamp 1624635492
transform 1 0 67712 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_721
timestamp 1624635492
transform 1 0 67436 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_716
timestamp 1624635492
transform 1 0 66976 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_732
timestamp 1624635492
transform 1 0 68448 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_728
timestamp 1624635492
transform 1 0 68080 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_729
timestamp 1624635492
transform 1 0 68172 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1624635492
transform -1 0 68816 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1624635492
transform -1 0 68816 0 -1 66912
box -38 -48 314 592
<< labels >>
rlabel metal3 s 69200 28296 70000 28416 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 53378 69200 53434 70000 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 45650 69200 45706 70000 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 37830 69200 37886 70000 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 30102 69200 30158 70000 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 22282 69200 22338 70000 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 14462 69200 14518 70000 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 6734 69200 6790 70000 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s 0 69232 800 69352 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s 0 64064 800 64184 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s 0 58896 800 59016 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 69200 33464 70000 33584 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s 0 53728 800 53848 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s 0 48424 800 48544 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s 0 43256 800 43376 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s 0 38088 800 38208 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s 0 32920 800 33040 6 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s 0 27752 800 27872 6 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s 0 22584 800 22704 6 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s 0 17280 800 17400 6 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s 0 12112 800 12232 6 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 69200 38768 70000 38888 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 69200 44072 70000 44192 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 69200 49376 70000 49496 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 69200 54680 70000 54800 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 69200 59984 70000 60104 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 69200 65288 70000 65408 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 68926 69200 68982 70000 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 61198 69200 61254 70000 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 69200 552 70000 672 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 69200 45432 70000 45552 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 69200 50736 70000 50856 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 69200 56040 70000 56160 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 69200 61208 70000 61328 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 69200 66512 70000 66632 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 66994 69200 67050 70000 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 59266 69200 59322 70000 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 51446 69200 51502 70000 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 43718 69200 43774 70000 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 35898 69200 35954 70000 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 69200 4496 70000 4616 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 28078 69200 28134 70000 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 20350 69200 20406 70000 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 12530 69200 12586 70000 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 4802 69200 4858 70000 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 io_in[24]
port 45 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 io_in[25]
port 46 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 io_in[26]
port 47 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 io_in[27]
port 48 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 io_in[28]
port 49 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 io_in[29]
port 50 nsew signal input
rlabel metal3 s 69200 8440 70000 8560 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 io_in[30]
port 52 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 io_in[31]
port 53 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 io_in[32]
port 54 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 io_in[33]
port 55 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 io_in[34]
port 56 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[35]
port 57 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 io_in[36]
port 58 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 io_in[37]
port 59 nsew signal input
rlabel metal3 s 69200 12384 70000 12504 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 69200 16328 70000 16448 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 69200 20272 70000 20392 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 69200 24216 70000 24336 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 69200 29520 70000 29640 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 69200 34824 70000 34944 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 69200 40128 70000 40248 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 69200 3136 70000 3256 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 69200 48016 70000 48136 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 69200 53320 70000 53440 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 69200 58624 70000 58744 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 69200 63928 70000 64048 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 69200 69232 70000 69352 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 63130 69200 63186 70000 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 55310 69200 55366 70000 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 47582 69200 47638 70000 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 39762 69200 39818 70000 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 32034 69200 32090 70000 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 69200 7080 70000 7200 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 24214 69200 24270 70000 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 16486 69200 16542 70000 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 8666 69200 8722 70000 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 938 69200 994 70000 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s 0 65288 800 65408 6 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s 0 60120 800 60240 6 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s 0 54952 800 55072 6 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s 0 49784 800 49904 6 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s 0 44616 800 44736 6 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s 0 39448 800 39568 6 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 69200 11024 70000 11144 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s 0 34144 800 34264 6 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s 0 28976 800 29096 6 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s 0 23808 800 23928 6 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s 0 18640 800 18760 6 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s 0 8304 800 8424 6 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s 0 552 800 672 6 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 69200 14968 70000 15088 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 69200 19048 70000 19168 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 69200 22992 70000 23112 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 69200 26936 70000 27056 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 69200 32240 70000 32360 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 69200 37544 70000 37664 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 69200 42712 70000 42832 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 69200 1776 70000 1896 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 69200 46792 70000 46912 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 69200 51960 70000 52080 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 69200 57264 70000 57384 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 69200 62568 70000 62688 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 69200 67872 70000 67992 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 65062 69200 65118 70000 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 57334 69200 57390 70000 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 49514 69200 49570 70000 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 41694 69200 41750 70000 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 33966 69200 34022 70000 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 69200 5720 70000 5840 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 26146 69200 26202 70000 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 18418 69200 18474 70000 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 10598 69200 10654 70000 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 2870 69200 2926 70000 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s 0 66648 800 66768 6 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s 0 61480 800 61600 6 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s 0 56312 800 56432 6 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s 0 51008 800 51128 6 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s 0 45840 800 45960 6 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s 0 40672 800 40792 6 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 69200 9800 70000 9920 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s 0 35504 800 35624 6 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s 0 30336 800 30456 6 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s 0 25168 800 25288 6 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s 0 20000 800 20120 6 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s 0 14696 800 14816 6 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s 0 5720 800 5840 6 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 69200 13744 70000 13864 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 69200 17688 70000 17808 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 69200 21632 70000 21752 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 69200 25576 70000 25696 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 69200 30880 70000 31000 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 69200 36184 70000 36304 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 69200 41488 70000 41608 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 15014 0 15070 800 6 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 57610 0 57666 800 6 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 58070 0 58126 800 6 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 58530 0 58586 800 6 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 58898 0 58954 800 6 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 59358 0 59414 800 6 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 59818 0 59874 800 6 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 60186 0 60242 800 6 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 60646 0 60702 800 6 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 61014 0 61070 800 6 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 61474 0 61530 800 6 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 61934 0 61990 800 6 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 62302 0 62358 800 6 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 62762 0 62818 800 6 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 63222 0 63278 800 6 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 63590 0 63646 800 6 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 64050 0 64106 800 6 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 64418 0 64474 800 6 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 64878 0 64934 800 6 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 65338 0 65394 800 6 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 65706 0 65762 800 6 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 19798 0 19854 800 6 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 66166 0 66222 800 6 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 66626 0 66682 800 6 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 66994 0 67050 800 6 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 67454 0 67510 800 6 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 67822 0 67878 800 6 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 68282 0 68338 800 6 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 68742 0 68798 800 6 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 69110 0 69166 800 6 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 20258 0 20314 800 6 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 21086 0 21142 800 6 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 22374 0 22430 800 6 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 22834 0 22890 800 6 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 23202 0 23258 800 6 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 15566 0 15622 800 6 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 23662 0 23718 800 6 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 24030 0 24086 800 6 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 24490 0 24546 800 6 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 24950 0 25006 800 6 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 25778 0 25834 800 6 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 26146 0 26202 800 6 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 26606 0 26662 800 6 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 27066 0 27122 800 6 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 27434 0 27490 800 6 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 27894 0 27950 800 6 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 28354 0 28410 800 6 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 28722 0 28778 800 6 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 29182 0 29238 800 6 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 29550 0 29606 800 6 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 30010 0 30066 800 6 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 30470 0 30526 800 6 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 30838 0 30894 800 6 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 31298 0 31354 800 6 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 31758 0 31814 800 6 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 16394 0 16450 800 6 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 32126 0 32182 800 6 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 32586 0 32642 800 6 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 32954 0 33010 800 6 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 33414 0 33470 800 6 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 33874 0 33930 800 6 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 34242 0 34298 800 6 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 34702 0 34758 800 6 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 35162 0 35218 800 6 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 35530 0 35586 800 6 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 35990 0 36046 800 6 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 16854 0 16910 800 6 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 36358 0 36414 800 6 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 36818 0 36874 800 6 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 37278 0 37334 800 6 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 37646 0 37702 800 6 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 38106 0 38162 800 6 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 38566 0 38622 800 6 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 38934 0 38990 800 6 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 39394 0 39450 800 6 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 40222 0 40278 800 6 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 40682 0 40738 800 6 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 41050 0 41106 800 6 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 41510 0 41566 800 6 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 41878 0 41934 800 6 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 42338 0 42394 800 6 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 42798 0 42854 800 6 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 43166 0 43222 800 6 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 43626 0 43682 800 6 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 44086 0 44142 800 6 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 44454 0 44510 800 6 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 44914 0 44970 800 6 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 45282 0 45338 800 6 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 45742 0 45798 800 6 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 46202 0 46258 800 6 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 46570 0 46626 800 6 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 47030 0 47086 800 6 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 47490 0 47546 800 6 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 47858 0 47914 800 6 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 48318 0 48374 800 6 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 48686 0 48742 800 6 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 49146 0 49202 800 6 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 49606 0 49662 800 6 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 49974 0 50030 800 6 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 50434 0 50490 800 6 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 50894 0 50950 800 6 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 51262 0 51318 800 6 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 51722 0 51778 800 6 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 52090 0 52146 800 6 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 52550 0 52606 800 6 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 53010 0 53066 800 6 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 18510 0 18566 800 6 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 53378 0 53434 800 6 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 53838 0 53894 800 6 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 54298 0 54354 800 6 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 54666 0 54722 800 6 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 55126 0 55182 800 6 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 55494 0 55550 800 6 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 55954 0 56010 800 6 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 56414 0 56470 800 6 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 56782 0 56838 800 6 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 57242 0 57298 800 6 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 user_clock2
port 527 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 69662 0 69718 800 6 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 69846 0 69902 800 6 user_irq[2]
port 530 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 294 0 350 800 6 wbs_ack_o
port 533 nsew signal tristate
rlabel metal2 s 846 0 902 800 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 386 0 442 800 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_dat_o[0]
port 599 nsew signal tristate
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[10]
port 600 nsew signal tristate
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_o[11]
port 601 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[12]
port 602 nsew signal tristate
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[13]
port 603 nsew signal tristate
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_o[14]
port 604 nsew signal tristate
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[15]
port 605 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[16]
port 606 nsew signal tristate
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[17]
port 607 nsew signal tristate
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[18]
port 608 nsew signal tristate
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[19]
port 609 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[1]
port 610 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[20]
port 611 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[21]
port 612 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[22]
port 613 nsew signal tristate
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[23]
port 614 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[24]
port 615 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[25]
port 616 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[26]
port 617 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[27]
port 618 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[28]
port 619 nsew signal tristate
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[29]
port 620 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 wbs_dat_o[2]
port 621 nsew signal tristate
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[30]
port 622 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[31]
port 623 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_o[3]
port 624 nsew signal tristate
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[4]
port 625 nsew signal tristate
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_o[5]
port 626 nsew signal tristate
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_o[6]
port 627 nsew signal tristate
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_o[7]
port 628 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[8]
port 629 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[9]
port 630 nsew signal tristate
rlabel metal2 s 1214 0 1270 800 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 64208 2128 64528 67504 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 67504 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 67504 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 34208 2176 34528 67504 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 24208 2176 24528 67504 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 67504 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 67504 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 59208 2128 59528 67504 6 VGND
port 644 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 67504 6 VGND
port 645 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 67504 6 VGND
port 646 nsew ground bidirectional
rlabel metal4 s 29208 2176 29528 67504 6 VGND
port 647 nsew ground bidirectional
rlabel metal4 s 19208 2176 19528 67504 6 VGND
port 648 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 67504 6 VGND
port 649 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
<< end >>
