magic
tech sky130A
magscale 1 2
timestamp 1626693475
<< viali >>
rect 12415 7938 12449 7972
rect 12319 7716 12353 7750
rect 12031 7642 12065 7676
rect 12511 7494 12545 7528
rect 13375 7124 13409 7158
rect 11935 7050 11969 7084
rect 12319 6976 12353 7010
rect 12895 6902 12929 6936
rect 13087 6902 13121 6936
rect 13279 6902 13313 6936
rect 11935 6310 11969 6344
rect 13375 6310 13409 6344
rect 14047 6310 14081 6344
rect 13183 6088 13217 6122
rect 13279 6088 13313 6122
rect 11839 6014 11873 6048
rect 12895 6014 12929 6048
rect 11071 5866 11105 5900
rect 12415 5496 12449 5530
rect 13375 5496 13409 5530
rect 12207 5422 12241 5456
rect 12319 5422 12353 5456
rect 11167 5348 11201 5382
rect 11839 5348 11873 5382
rect 11359 5274 11393 5308
rect 12895 5274 12929 5308
rect 13087 5274 13121 5308
rect 13279 5274 13313 5308
rect 10687 5052 10721 5086
rect 13951 5052 13985 5086
rect 11839 4682 11873 4716
rect 12991 4682 13025 4716
rect 12319 4386 12353 4420
rect 11263 4312 11297 4346
rect 11935 4312 11969 4346
rect 12031 4312 12065 4346
rect 12607 3424 12641 3458
<< metal1 >>
rect 1152 16306 14784 16331
rect 1152 16254 3312 16306
rect 3364 16254 3376 16306
rect 3428 16254 3440 16306
rect 3492 16254 3504 16306
rect 3556 16254 7878 16306
rect 7930 16254 7942 16306
rect 7994 16254 8006 16306
rect 8058 16254 8070 16306
rect 8122 16254 12443 16306
rect 12495 16254 12507 16306
rect 12559 16254 12571 16306
rect 12623 16254 12635 16306
rect 12687 16254 14784 16306
rect 1152 16229 14784 16254
rect 1152 15492 14784 15517
rect 1152 15440 5595 15492
rect 5647 15440 5659 15492
rect 5711 15440 5723 15492
rect 5775 15440 5787 15492
rect 5839 15440 10160 15492
rect 10212 15440 10224 15492
rect 10276 15440 10288 15492
rect 10340 15440 10352 15492
rect 10404 15440 14784 15492
rect 1152 15415 14784 15440
rect 1152 14678 14784 14703
rect 1152 14626 3312 14678
rect 3364 14626 3376 14678
rect 3428 14626 3440 14678
rect 3492 14626 3504 14678
rect 3556 14626 7878 14678
rect 7930 14626 7942 14678
rect 7994 14626 8006 14678
rect 8058 14626 8070 14678
rect 8122 14626 12443 14678
rect 12495 14626 12507 14678
rect 12559 14626 12571 14678
rect 12623 14626 12635 14678
rect 12687 14626 14784 14678
rect 1152 14601 14784 14626
rect 1152 13864 14784 13889
rect 1152 13812 5595 13864
rect 5647 13812 5659 13864
rect 5711 13812 5723 13864
rect 5775 13812 5787 13864
rect 5839 13812 10160 13864
rect 10212 13812 10224 13864
rect 10276 13812 10288 13864
rect 10340 13812 10352 13864
rect 10404 13812 14784 13864
rect 1152 13787 14784 13812
rect 1152 13050 14784 13075
rect 1152 12998 3312 13050
rect 3364 12998 3376 13050
rect 3428 12998 3440 13050
rect 3492 12998 3504 13050
rect 3556 12998 7878 13050
rect 7930 12998 7942 13050
rect 7994 12998 8006 13050
rect 8058 12998 8070 13050
rect 8122 12998 12443 13050
rect 12495 12998 12507 13050
rect 12559 12998 12571 13050
rect 12623 12998 12635 13050
rect 12687 12998 14784 13050
rect 1152 12973 14784 12998
rect 1152 12236 14784 12261
rect 1152 12184 5595 12236
rect 5647 12184 5659 12236
rect 5711 12184 5723 12236
rect 5775 12184 5787 12236
rect 5839 12184 10160 12236
rect 10212 12184 10224 12236
rect 10276 12184 10288 12236
rect 10340 12184 10352 12236
rect 10404 12184 14784 12236
rect 1152 12159 14784 12184
rect 1152 11422 14784 11447
rect 1152 11370 3312 11422
rect 3364 11370 3376 11422
rect 3428 11370 3440 11422
rect 3492 11370 3504 11422
rect 3556 11370 7878 11422
rect 7930 11370 7942 11422
rect 7994 11370 8006 11422
rect 8058 11370 8070 11422
rect 8122 11370 12443 11422
rect 12495 11370 12507 11422
rect 12559 11370 12571 11422
rect 12623 11370 12635 11422
rect 12687 11370 14784 11422
rect 1152 11345 14784 11370
rect 1152 10608 14784 10633
rect 1152 10556 5595 10608
rect 5647 10556 5659 10608
rect 5711 10556 5723 10608
rect 5775 10556 5787 10608
rect 5839 10556 10160 10608
rect 10212 10556 10224 10608
rect 10276 10556 10288 10608
rect 10340 10556 10352 10608
rect 10404 10556 14784 10608
rect 1152 10531 14784 10556
rect 1152 9794 14784 9819
rect 1152 9742 3312 9794
rect 3364 9742 3376 9794
rect 3428 9742 3440 9794
rect 3492 9742 3504 9794
rect 3556 9742 7878 9794
rect 7930 9742 7942 9794
rect 7994 9742 8006 9794
rect 8058 9742 8070 9794
rect 8122 9742 12443 9794
rect 12495 9742 12507 9794
rect 12559 9742 12571 9794
rect 12623 9742 12635 9794
rect 12687 9742 14784 9794
rect 1152 9717 14784 9742
rect 1152 8980 14784 9005
rect 1152 8928 5595 8980
rect 5647 8928 5659 8980
rect 5711 8928 5723 8980
rect 5775 8928 5787 8980
rect 5839 8928 10160 8980
rect 10212 8928 10224 8980
rect 10276 8928 10288 8980
rect 10340 8928 10352 8980
rect 10404 8928 14784 8980
rect 1152 8903 14784 8928
rect 12880 8595 12886 8647
rect 12938 8635 12944 8647
rect 13360 8635 13366 8647
rect 12938 8607 13366 8635
rect 12938 8595 12944 8607
rect 13360 8595 13366 8607
rect 13418 8595 13424 8647
rect 1152 8166 14784 8191
rect 1152 8114 3312 8166
rect 3364 8114 3376 8166
rect 3428 8114 3440 8166
rect 3492 8114 3504 8166
rect 3556 8114 7878 8166
rect 7930 8114 7942 8166
rect 7994 8114 8006 8166
rect 8058 8114 8070 8166
rect 8122 8114 12443 8166
rect 12495 8114 12507 8166
rect 12559 8114 12571 8166
rect 12623 8114 12635 8166
rect 12687 8114 14784 8166
rect 1152 8089 14784 8114
rect 12403 7972 12461 7978
rect 12403 7938 12415 7972
rect 12449 7969 12461 7972
rect 13360 7969 13366 7981
rect 12449 7941 13366 7969
rect 12449 7938 12461 7941
rect 12403 7932 12461 7938
rect 13360 7929 13366 7941
rect 13418 7929 13424 7981
rect 12307 7750 12365 7756
rect 12307 7716 12319 7750
rect 12353 7716 12365 7750
rect 12307 7710 12365 7716
rect 12016 7673 12022 7685
rect 11977 7645 12022 7673
rect 12016 7633 12022 7645
rect 12074 7633 12080 7685
rect 12322 7673 12350 7710
rect 13168 7673 13174 7685
rect 12322 7645 13174 7673
rect 13168 7633 13174 7645
rect 13226 7633 13232 7685
rect 12499 7528 12557 7534
rect 12499 7494 12511 7528
rect 12545 7525 12557 7528
rect 13264 7525 13270 7537
rect 12545 7497 13270 7525
rect 12545 7494 12557 7497
rect 12499 7488 12557 7494
rect 13264 7485 13270 7497
rect 13322 7485 13328 7537
rect 1152 7352 14784 7377
rect 1152 7300 5595 7352
rect 5647 7300 5659 7352
rect 5711 7300 5723 7352
rect 5775 7300 5787 7352
rect 5839 7300 10160 7352
rect 10212 7300 10224 7352
rect 10276 7300 10288 7352
rect 10340 7300 10352 7352
rect 10404 7300 14784 7352
rect 1152 7275 14784 7300
rect 13360 7155 13366 7167
rect 13321 7127 13366 7155
rect 13360 7115 13366 7127
rect 13418 7115 13424 7167
rect 11923 7084 11981 7090
rect 11923 7050 11935 7084
rect 11969 7081 11981 7084
rect 12016 7081 12022 7093
rect 11969 7053 12022 7081
rect 11969 7050 11981 7053
rect 11923 7044 11981 7050
rect 12016 7041 12022 7053
rect 12074 7041 12080 7093
rect 12304 7007 12310 7019
rect 12265 6979 12310 7007
rect 12304 6967 12310 6979
rect 12362 6967 12368 7019
rect 12880 6933 12886 6945
rect 12841 6905 12886 6933
rect 12880 6893 12886 6905
rect 12938 6893 12944 6945
rect 13075 6936 13133 6942
rect 13075 6902 13087 6936
rect 13121 6902 13133 6936
rect 13264 6933 13270 6945
rect 13225 6905 13270 6933
rect 13075 6896 13133 6902
rect 13090 6859 13118 6896
rect 13264 6893 13270 6905
rect 13322 6893 13328 6945
rect 13360 6859 13366 6871
rect 13090 6831 13366 6859
rect 13360 6819 13366 6831
rect 13418 6819 13424 6871
rect 1152 6538 14784 6563
rect 1152 6486 3312 6538
rect 3364 6486 3376 6538
rect 3428 6486 3440 6538
rect 3492 6486 3504 6538
rect 3556 6486 7878 6538
rect 7930 6486 7942 6538
rect 7994 6486 8006 6538
rect 8058 6486 8070 6538
rect 8122 6486 12443 6538
rect 12495 6486 12507 6538
rect 12559 6486 12571 6538
rect 12623 6486 12635 6538
rect 12687 6486 14784 6538
rect 1152 6461 14784 6486
rect 11923 6344 11981 6350
rect 11923 6310 11935 6344
rect 11969 6341 11981 6344
rect 12880 6341 12886 6353
rect 11969 6313 12886 6341
rect 11969 6310 11981 6313
rect 11923 6304 11981 6310
rect 12880 6301 12886 6313
rect 12938 6301 12944 6353
rect 13168 6301 13174 6353
rect 13226 6341 13232 6353
rect 13363 6344 13421 6350
rect 13363 6341 13375 6344
rect 13226 6313 13375 6341
rect 13226 6301 13232 6313
rect 13363 6310 13375 6313
rect 13409 6310 13421 6344
rect 14032 6341 14038 6353
rect 13993 6313 14038 6341
rect 13363 6304 13421 6310
rect 14032 6301 14038 6313
rect 14090 6301 14096 6353
rect 14050 6193 14078 6301
rect 13186 6165 14078 6193
rect 12976 6079 12982 6131
rect 13034 6119 13040 6131
rect 13186 6128 13214 6165
rect 13171 6122 13229 6128
rect 13171 6119 13183 6122
rect 13034 6091 13183 6119
rect 13034 6079 13040 6091
rect 13171 6088 13183 6091
rect 13217 6088 13229 6122
rect 13171 6082 13229 6088
rect 13267 6122 13325 6128
rect 13267 6088 13279 6122
rect 13313 6119 13325 6122
rect 13360 6119 13366 6131
rect 13313 6091 13366 6119
rect 13313 6088 13325 6091
rect 13267 6082 13325 6088
rect 13360 6079 13366 6091
rect 13418 6079 13424 6131
rect 11824 6045 11830 6057
rect 11785 6017 11830 6045
rect 11824 6005 11830 6017
rect 11882 6005 11888 6057
rect 12880 6045 12886 6057
rect 12841 6017 12886 6045
rect 12880 6005 12886 6017
rect 12938 6005 12944 6057
rect 11056 5897 11062 5909
rect 11017 5869 11062 5897
rect 11056 5857 11062 5869
rect 11114 5857 11120 5909
rect 1152 5724 14784 5749
rect 1152 5672 5595 5724
rect 5647 5672 5659 5724
rect 5711 5672 5723 5724
rect 5775 5672 5787 5724
rect 5839 5672 10160 5724
rect 10212 5672 10224 5724
rect 10276 5672 10288 5724
rect 10340 5672 10352 5724
rect 10404 5672 14784 5724
rect 1152 5647 14784 5672
rect 12400 5527 12406 5539
rect 12361 5499 12406 5527
rect 12400 5487 12406 5499
rect 12458 5487 12464 5539
rect 13360 5527 13366 5539
rect 13321 5499 13366 5527
rect 13360 5487 13366 5499
rect 13418 5487 13424 5539
rect 12208 5462 12214 5465
rect 12195 5456 12214 5462
rect 12195 5422 12207 5456
rect 12195 5416 12214 5422
rect 12208 5413 12214 5416
rect 12266 5413 12272 5465
rect 12307 5456 12365 5462
rect 12307 5422 12319 5456
rect 12353 5453 12365 5456
rect 12496 5453 12502 5465
rect 12353 5425 12502 5453
rect 12353 5422 12365 5425
rect 12307 5416 12365 5422
rect 12496 5413 12502 5425
rect 12554 5413 12560 5465
rect 10672 5339 10678 5391
rect 10730 5379 10736 5391
rect 11056 5379 11062 5391
rect 10730 5351 11062 5379
rect 10730 5339 10736 5351
rect 11056 5339 11062 5351
rect 11114 5379 11120 5391
rect 11155 5382 11213 5388
rect 11155 5379 11167 5382
rect 11114 5351 11167 5379
rect 11114 5339 11120 5351
rect 11155 5348 11167 5351
rect 11201 5348 11213 5382
rect 11824 5379 11830 5391
rect 11785 5351 11830 5379
rect 11155 5342 11213 5348
rect 11170 5231 11198 5342
rect 11824 5339 11830 5351
rect 11882 5339 11888 5391
rect 11347 5308 11405 5314
rect 11347 5274 11359 5308
rect 11393 5305 11405 5308
rect 12880 5305 12886 5317
rect 11393 5277 12886 5305
rect 11393 5274 11405 5277
rect 11347 5268 11405 5274
rect 12880 5265 12886 5277
rect 12938 5265 12944 5317
rect 13075 5308 13133 5314
rect 13075 5274 13087 5308
rect 13121 5274 13133 5308
rect 13075 5268 13133 5274
rect 12496 5231 12502 5243
rect 11170 5203 12502 5231
rect 12496 5191 12502 5203
rect 12554 5191 12560 5243
rect 10672 5083 10678 5095
rect 10633 5055 10678 5083
rect 10672 5043 10678 5055
rect 10730 5043 10736 5095
rect 12208 5043 12214 5095
rect 12266 5083 12272 5095
rect 12880 5083 12886 5095
rect 12266 5055 12886 5083
rect 12266 5043 12272 5055
rect 12880 5043 12886 5055
rect 12938 5083 12944 5095
rect 13090 5083 13118 5268
rect 13168 5265 13174 5317
rect 13226 5305 13232 5317
rect 13267 5308 13325 5314
rect 13267 5305 13279 5308
rect 13226 5277 13279 5305
rect 13226 5265 13232 5277
rect 13267 5274 13279 5277
rect 13313 5274 13325 5308
rect 13267 5268 13325 5274
rect 13939 5086 13997 5092
rect 13939 5083 13951 5086
rect 12938 5055 13951 5083
rect 12938 5043 12944 5055
rect 13939 5052 13951 5055
rect 13985 5052 13997 5086
rect 13939 5046 13997 5052
rect 1152 4910 14784 4935
rect 1152 4858 3312 4910
rect 3364 4858 3376 4910
rect 3428 4858 3440 4910
rect 3492 4858 3504 4910
rect 3556 4858 7878 4910
rect 7930 4858 7942 4910
rect 7994 4858 8006 4910
rect 8058 4858 8070 4910
rect 8122 4858 12443 4910
rect 12495 4858 12507 4910
rect 12559 4858 12571 4910
rect 12623 4858 12635 4910
rect 12687 4858 14784 4910
rect 1152 4833 14784 4858
rect 11824 4713 11830 4725
rect 11785 4685 11830 4713
rect 11824 4673 11830 4685
rect 11882 4673 11888 4725
rect 12976 4713 12982 4725
rect 12937 4685 12982 4713
rect 12976 4673 12982 4685
rect 13034 4673 13040 4725
rect 12304 4417 12310 4429
rect 12265 4389 12310 4417
rect 12304 4377 12310 4389
rect 12362 4377 12368 4429
rect 11251 4346 11309 4352
rect 11251 4312 11263 4346
rect 11297 4343 11309 4346
rect 11923 4346 11981 4352
rect 11923 4343 11935 4346
rect 11297 4315 11935 4343
rect 11297 4312 11309 4315
rect 11251 4306 11309 4312
rect 11923 4312 11935 4315
rect 11969 4312 11981 4346
rect 11923 4306 11981 4312
rect 12019 4346 12077 4352
rect 12019 4312 12031 4346
rect 12065 4343 12077 4346
rect 12976 4343 12982 4355
rect 12065 4315 12982 4343
rect 12065 4312 12077 4315
rect 12019 4306 12077 4312
rect 8176 4229 8182 4281
rect 8234 4269 8240 4281
rect 10672 4269 10678 4281
rect 8234 4241 10678 4269
rect 8234 4229 8240 4241
rect 10672 4229 10678 4241
rect 10730 4269 10736 4281
rect 11266 4269 11294 4306
rect 12976 4303 12982 4315
rect 13034 4303 13040 4355
rect 10730 4241 11294 4269
rect 10730 4229 10736 4241
rect 1152 4096 14784 4121
rect 1152 4044 5595 4096
rect 5647 4044 5659 4096
rect 5711 4044 5723 4096
rect 5775 4044 5787 4096
rect 5839 4044 10160 4096
rect 10212 4044 10224 4096
rect 10276 4044 10288 4096
rect 10340 4044 10352 4096
rect 10404 4044 14784 4096
rect 1152 4019 14784 4044
rect 12595 3458 12653 3464
rect 12595 3424 12607 3458
rect 12641 3455 12653 3458
rect 12880 3455 12886 3467
rect 12641 3427 12886 3455
rect 12641 3424 12653 3427
rect 12595 3418 12653 3424
rect 12880 3415 12886 3427
rect 12938 3415 12944 3467
rect 1152 3282 14784 3307
rect 1152 3230 3312 3282
rect 3364 3230 3376 3282
rect 3428 3230 3440 3282
rect 3492 3230 3504 3282
rect 3556 3230 7878 3282
rect 7930 3230 7942 3282
rect 7994 3230 8006 3282
rect 8058 3230 8070 3282
rect 8122 3230 12443 3282
rect 12495 3230 12507 3282
rect 12559 3230 12571 3282
rect 12623 3230 12635 3282
rect 12687 3230 14784 3282
rect 1152 3205 14784 3230
<< via1 >>
rect 3312 16254 3364 16306
rect 3376 16254 3428 16306
rect 3440 16254 3492 16306
rect 3504 16254 3556 16306
rect 7878 16254 7930 16306
rect 7942 16254 7994 16306
rect 8006 16254 8058 16306
rect 8070 16254 8122 16306
rect 12443 16254 12495 16306
rect 12507 16254 12559 16306
rect 12571 16254 12623 16306
rect 12635 16254 12687 16306
rect 5595 15440 5647 15492
rect 5659 15440 5711 15492
rect 5723 15440 5775 15492
rect 5787 15440 5839 15492
rect 10160 15440 10212 15492
rect 10224 15440 10276 15492
rect 10288 15440 10340 15492
rect 10352 15440 10404 15492
rect 3312 14626 3364 14678
rect 3376 14626 3428 14678
rect 3440 14626 3492 14678
rect 3504 14626 3556 14678
rect 7878 14626 7930 14678
rect 7942 14626 7994 14678
rect 8006 14626 8058 14678
rect 8070 14626 8122 14678
rect 12443 14626 12495 14678
rect 12507 14626 12559 14678
rect 12571 14626 12623 14678
rect 12635 14626 12687 14678
rect 5595 13812 5647 13864
rect 5659 13812 5711 13864
rect 5723 13812 5775 13864
rect 5787 13812 5839 13864
rect 10160 13812 10212 13864
rect 10224 13812 10276 13864
rect 10288 13812 10340 13864
rect 10352 13812 10404 13864
rect 3312 12998 3364 13050
rect 3376 12998 3428 13050
rect 3440 12998 3492 13050
rect 3504 12998 3556 13050
rect 7878 12998 7930 13050
rect 7942 12998 7994 13050
rect 8006 12998 8058 13050
rect 8070 12998 8122 13050
rect 12443 12998 12495 13050
rect 12507 12998 12559 13050
rect 12571 12998 12623 13050
rect 12635 12998 12687 13050
rect 5595 12184 5647 12236
rect 5659 12184 5711 12236
rect 5723 12184 5775 12236
rect 5787 12184 5839 12236
rect 10160 12184 10212 12236
rect 10224 12184 10276 12236
rect 10288 12184 10340 12236
rect 10352 12184 10404 12236
rect 3312 11370 3364 11422
rect 3376 11370 3428 11422
rect 3440 11370 3492 11422
rect 3504 11370 3556 11422
rect 7878 11370 7930 11422
rect 7942 11370 7994 11422
rect 8006 11370 8058 11422
rect 8070 11370 8122 11422
rect 12443 11370 12495 11422
rect 12507 11370 12559 11422
rect 12571 11370 12623 11422
rect 12635 11370 12687 11422
rect 5595 10556 5647 10608
rect 5659 10556 5711 10608
rect 5723 10556 5775 10608
rect 5787 10556 5839 10608
rect 10160 10556 10212 10608
rect 10224 10556 10276 10608
rect 10288 10556 10340 10608
rect 10352 10556 10404 10608
rect 3312 9742 3364 9794
rect 3376 9742 3428 9794
rect 3440 9742 3492 9794
rect 3504 9742 3556 9794
rect 7878 9742 7930 9794
rect 7942 9742 7994 9794
rect 8006 9742 8058 9794
rect 8070 9742 8122 9794
rect 12443 9742 12495 9794
rect 12507 9742 12559 9794
rect 12571 9742 12623 9794
rect 12635 9742 12687 9794
rect 5595 8928 5647 8980
rect 5659 8928 5711 8980
rect 5723 8928 5775 8980
rect 5787 8928 5839 8980
rect 10160 8928 10212 8980
rect 10224 8928 10276 8980
rect 10288 8928 10340 8980
rect 10352 8928 10404 8980
rect 12886 8595 12938 8647
rect 13366 8595 13418 8647
rect 3312 8114 3364 8166
rect 3376 8114 3428 8166
rect 3440 8114 3492 8166
rect 3504 8114 3556 8166
rect 7878 8114 7930 8166
rect 7942 8114 7994 8166
rect 8006 8114 8058 8166
rect 8070 8114 8122 8166
rect 12443 8114 12495 8166
rect 12507 8114 12559 8166
rect 12571 8114 12623 8166
rect 12635 8114 12687 8166
rect 13366 7929 13418 7981
rect 12022 7676 12074 7685
rect 12022 7642 12031 7676
rect 12031 7642 12065 7676
rect 12065 7642 12074 7676
rect 12022 7633 12074 7642
rect 13174 7633 13226 7685
rect 13270 7485 13322 7537
rect 5595 7300 5647 7352
rect 5659 7300 5711 7352
rect 5723 7300 5775 7352
rect 5787 7300 5839 7352
rect 10160 7300 10212 7352
rect 10224 7300 10276 7352
rect 10288 7300 10340 7352
rect 10352 7300 10404 7352
rect 13366 7158 13418 7167
rect 13366 7124 13375 7158
rect 13375 7124 13409 7158
rect 13409 7124 13418 7158
rect 13366 7115 13418 7124
rect 12022 7041 12074 7093
rect 12310 7010 12362 7019
rect 12310 6976 12319 7010
rect 12319 6976 12353 7010
rect 12353 6976 12362 7010
rect 12310 6967 12362 6976
rect 12886 6936 12938 6945
rect 12886 6902 12895 6936
rect 12895 6902 12929 6936
rect 12929 6902 12938 6936
rect 12886 6893 12938 6902
rect 13270 6936 13322 6945
rect 13270 6902 13279 6936
rect 13279 6902 13313 6936
rect 13313 6902 13322 6936
rect 13270 6893 13322 6902
rect 13366 6819 13418 6871
rect 3312 6486 3364 6538
rect 3376 6486 3428 6538
rect 3440 6486 3492 6538
rect 3504 6486 3556 6538
rect 7878 6486 7930 6538
rect 7942 6486 7994 6538
rect 8006 6486 8058 6538
rect 8070 6486 8122 6538
rect 12443 6486 12495 6538
rect 12507 6486 12559 6538
rect 12571 6486 12623 6538
rect 12635 6486 12687 6538
rect 12886 6301 12938 6353
rect 13174 6301 13226 6353
rect 14038 6344 14090 6353
rect 14038 6310 14047 6344
rect 14047 6310 14081 6344
rect 14081 6310 14090 6344
rect 14038 6301 14090 6310
rect 12982 6079 13034 6131
rect 13366 6079 13418 6131
rect 11830 6048 11882 6057
rect 11830 6014 11839 6048
rect 11839 6014 11873 6048
rect 11873 6014 11882 6048
rect 11830 6005 11882 6014
rect 12886 6048 12938 6057
rect 12886 6014 12895 6048
rect 12895 6014 12929 6048
rect 12929 6014 12938 6048
rect 12886 6005 12938 6014
rect 11062 5900 11114 5909
rect 11062 5866 11071 5900
rect 11071 5866 11105 5900
rect 11105 5866 11114 5900
rect 11062 5857 11114 5866
rect 5595 5672 5647 5724
rect 5659 5672 5711 5724
rect 5723 5672 5775 5724
rect 5787 5672 5839 5724
rect 10160 5672 10212 5724
rect 10224 5672 10276 5724
rect 10288 5672 10340 5724
rect 10352 5672 10404 5724
rect 12406 5530 12458 5539
rect 12406 5496 12415 5530
rect 12415 5496 12449 5530
rect 12449 5496 12458 5530
rect 12406 5487 12458 5496
rect 13366 5530 13418 5539
rect 13366 5496 13375 5530
rect 13375 5496 13409 5530
rect 13409 5496 13418 5530
rect 13366 5487 13418 5496
rect 12214 5456 12266 5465
rect 12214 5422 12241 5456
rect 12241 5422 12266 5456
rect 12214 5413 12266 5422
rect 12502 5413 12554 5465
rect 10678 5339 10730 5391
rect 11062 5339 11114 5391
rect 11830 5382 11882 5391
rect 11830 5348 11839 5382
rect 11839 5348 11873 5382
rect 11873 5348 11882 5382
rect 11830 5339 11882 5348
rect 12886 5308 12938 5317
rect 12886 5274 12895 5308
rect 12895 5274 12929 5308
rect 12929 5274 12938 5308
rect 12886 5265 12938 5274
rect 12502 5191 12554 5243
rect 10678 5086 10730 5095
rect 10678 5052 10687 5086
rect 10687 5052 10721 5086
rect 10721 5052 10730 5086
rect 10678 5043 10730 5052
rect 12214 5043 12266 5095
rect 12886 5043 12938 5095
rect 13174 5265 13226 5317
rect 3312 4858 3364 4910
rect 3376 4858 3428 4910
rect 3440 4858 3492 4910
rect 3504 4858 3556 4910
rect 7878 4858 7930 4910
rect 7942 4858 7994 4910
rect 8006 4858 8058 4910
rect 8070 4858 8122 4910
rect 12443 4858 12495 4910
rect 12507 4858 12559 4910
rect 12571 4858 12623 4910
rect 12635 4858 12687 4910
rect 11830 4716 11882 4725
rect 11830 4682 11839 4716
rect 11839 4682 11873 4716
rect 11873 4682 11882 4716
rect 11830 4673 11882 4682
rect 12982 4716 13034 4725
rect 12982 4682 12991 4716
rect 12991 4682 13025 4716
rect 13025 4682 13034 4716
rect 12982 4673 13034 4682
rect 12310 4420 12362 4429
rect 12310 4386 12319 4420
rect 12319 4386 12353 4420
rect 12353 4386 12362 4420
rect 12310 4377 12362 4386
rect 8182 4229 8234 4281
rect 10678 4229 10730 4281
rect 12982 4303 13034 4355
rect 5595 4044 5647 4096
rect 5659 4044 5711 4096
rect 5723 4044 5775 4096
rect 5787 4044 5839 4096
rect 10160 4044 10212 4096
rect 10224 4044 10276 4096
rect 10288 4044 10340 4096
rect 10352 4044 10404 4096
rect 12886 3415 12938 3467
rect 3312 3230 3364 3282
rect 3376 3230 3428 3282
rect 3440 3230 3492 3282
rect 3504 3230 3556 3282
rect 7878 3230 7930 3282
rect 7942 3230 7994 3282
rect 8006 3230 8058 3282
rect 8070 3230 8122 3282
rect 12443 3230 12495 3282
rect 12507 3230 12559 3282
rect 12571 3230 12623 3282
rect 12635 3230 12687 3282
<< metal2 >>
rect 12884 16678 12940 16687
rect 12884 16613 12940 16622
rect 3286 16308 3582 16331
rect 3342 16306 3366 16308
rect 3422 16306 3446 16308
rect 3502 16306 3526 16308
rect 3364 16254 3366 16306
rect 3428 16254 3440 16306
rect 3502 16254 3504 16306
rect 3342 16252 3366 16254
rect 3422 16252 3446 16254
rect 3502 16252 3526 16254
rect 3286 16229 3582 16252
rect 7852 16308 8148 16331
rect 7908 16306 7932 16308
rect 7988 16306 8012 16308
rect 8068 16306 8092 16308
rect 7930 16254 7932 16306
rect 7994 16254 8006 16306
rect 8068 16254 8070 16306
rect 7908 16252 7932 16254
rect 7988 16252 8012 16254
rect 8068 16252 8092 16254
rect 7852 16229 8148 16252
rect 12417 16308 12713 16331
rect 12473 16306 12497 16308
rect 12553 16306 12577 16308
rect 12633 16306 12657 16308
rect 12495 16254 12497 16306
rect 12559 16254 12571 16306
rect 12633 16254 12635 16306
rect 12473 16252 12497 16254
rect 12553 16252 12577 16254
rect 12633 16252 12657 16254
rect 12417 16229 12713 16252
rect 5569 15494 5865 15517
rect 5625 15492 5649 15494
rect 5705 15492 5729 15494
rect 5785 15492 5809 15494
rect 5647 15440 5649 15492
rect 5711 15440 5723 15492
rect 5785 15440 5787 15492
rect 5625 15438 5649 15440
rect 5705 15438 5729 15440
rect 5785 15438 5809 15440
rect 5569 15415 5865 15438
rect 10134 15494 10430 15517
rect 10190 15492 10214 15494
rect 10270 15492 10294 15494
rect 10350 15492 10374 15494
rect 10212 15440 10214 15492
rect 10276 15440 10288 15492
rect 10350 15440 10352 15492
rect 10190 15438 10214 15440
rect 10270 15438 10294 15440
rect 10350 15438 10374 15440
rect 10134 15415 10430 15438
rect 3286 14680 3582 14703
rect 3342 14678 3366 14680
rect 3422 14678 3446 14680
rect 3502 14678 3526 14680
rect 3364 14626 3366 14678
rect 3428 14626 3440 14678
rect 3502 14626 3504 14678
rect 3342 14624 3366 14626
rect 3422 14624 3446 14626
rect 3502 14624 3526 14626
rect 3286 14601 3582 14624
rect 7852 14680 8148 14703
rect 7908 14678 7932 14680
rect 7988 14678 8012 14680
rect 8068 14678 8092 14680
rect 7930 14626 7932 14678
rect 7994 14626 8006 14678
rect 8068 14626 8070 14678
rect 7908 14624 7932 14626
rect 7988 14624 8012 14626
rect 8068 14624 8092 14626
rect 7852 14601 8148 14624
rect 12417 14680 12713 14703
rect 12473 14678 12497 14680
rect 12553 14678 12577 14680
rect 12633 14678 12657 14680
rect 12495 14626 12497 14678
rect 12559 14626 12571 14678
rect 12633 14626 12635 14678
rect 12473 14624 12497 14626
rect 12553 14624 12577 14626
rect 12633 14624 12657 14626
rect 12417 14601 12713 14624
rect 5569 13866 5865 13889
rect 5625 13864 5649 13866
rect 5705 13864 5729 13866
rect 5785 13864 5809 13866
rect 5647 13812 5649 13864
rect 5711 13812 5723 13864
rect 5785 13812 5787 13864
rect 5625 13810 5649 13812
rect 5705 13810 5729 13812
rect 5785 13810 5809 13812
rect 5569 13787 5865 13810
rect 10134 13866 10430 13889
rect 10190 13864 10214 13866
rect 10270 13864 10294 13866
rect 10350 13864 10374 13866
rect 10212 13812 10214 13864
rect 10276 13812 10288 13864
rect 10350 13812 10352 13864
rect 10190 13810 10214 13812
rect 10270 13810 10294 13812
rect 10350 13810 10374 13812
rect 10134 13787 10430 13810
rect 3286 13052 3582 13075
rect 3342 13050 3366 13052
rect 3422 13050 3446 13052
rect 3502 13050 3526 13052
rect 3364 12998 3366 13050
rect 3428 12998 3440 13050
rect 3502 12998 3504 13050
rect 3342 12996 3366 12998
rect 3422 12996 3446 12998
rect 3502 12996 3526 12998
rect 3286 12973 3582 12996
rect 7852 13052 8148 13075
rect 7908 13050 7932 13052
rect 7988 13050 8012 13052
rect 8068 13050 8092 13052
rect 7930 12998 7932 13050
rect 7994 12998 8006 13050
rect 8068 12998 8070 13050
rect 7908 12996 7932 12998
rect 7988 12996 8012 12998
rect 8068 12996 8092 12998
rect 7852 12973 8148 12996
rect 12417 13052 12713 13075
rect 12473 13050 12497 13052
rect 12553 13050 12577 13052
rect 12633 13050 12657 13052
rect 12495 12998 12497 13050
rect 12559 12998 12571 13050
rect 12633 12998 12635 13050
rect 12473 12996 12497 12998
rect 12553 12996 12577 12998
rect 12633 12996 12657 12998
rect 12417 12973 12713 12996
rect 5569 12238 5865 12261
rect 5625 12236 5649 12238
rect 5705 12236 5729 12238
rect 5785 12236 5809 12238
rect 5647 12184 5649 12236
rect 5711 12184 5723 12236
rect 5785 12184 5787 12236
rect 5625 12182 5649 12184
rect 5705 12182 5729 12184
rect 5785 12182 5809 12184
rect 5569 12159 5865 12182
rect 10134 12238 10430 12261
rect 10190 12236 10214 12238
rect 10270 12236 10294 12238
rect 10350 12236 10374 12238
rect 10212 12184 10214 12236
rect 10276 12184 10288 12236
rect 10350 12184 10352 12236
rect 10190 12182 10214 12184
rect 10270 12182 10294 12184
rect 10350 12182 10374 12184
rect 10134 12159 10430 12182
rect 3286 11424 3582 11447
rect 3342 11422 3366 11424
rect 3422 11422 3446 11424
rect 3502 11422 3526 11424
rect 3364 11370 3366 11422
rect 3428 11370 3440 11422
rect 3502 11370 3504 11422
rect 3342 11368 3366 11370
rect 3422 11368 3446 11370
rect 3502 11368 3526 11370
rect 3286 11345 3582 11368
rect 7852 11424 8148 11447
rect 7908 11422 7932 11424
rect 7988 11422 8012 11424
rect 8068 11422 8092 11424
rect 7930 11370 7932 11422
rect 7994 11370 8006 11422
rect 8068 11370 8070 11422
rect 7908 11368 7932 11370
rect 7988 11368 8012 11370
rect 8068 11368 8092 11370
rect 7852 11345 8148 11368
rect 12417 11424 12713 11447
rect 12473 11422 12497 11424
rect 12553 11422 12577 11424
rect 12633 11422 12657 11424
rect 12495 11370 12497 11422
rect 12559 11370 12571 11422
rect 12633 11370 12635 11422
rect 12473 11368 12497 11370
rect 12553 11368 12577 11370
rect 12633 11368 12657 11370
rect 12417 11345 12713 11368
rect 5569 10610 5865 10633
rect 5625 10608 5649 10610
rect 5705 10608 5729 10610
rect 5785 10608 5809 10610
rect 5647 10556 5649 10608
rect 5711 10556 5723 10608
rect 5785 10556 5787 10608
rect 5625 10554 5649 10556
rect 5705 10554 5729 10556
rect 5785 10554 5809 10556
rect 5569 10531 5865 10554
rect 10134 10610 10430 10633
rect 10190 10608 10214 10610
rect 10270 10608 10294 10610
rect 10350 10608 10374 10610
rect 10212 10556 10214 10608
rect 10276 10556 10288 10608
rect 10350 10556 10352 10608
rect 10190 10554 10214 10556
rect 10270 10554 10294 10556
rect 10350 10554 10374 10556
rect 10134 10531 10430 10554
rect 3286 9796 3582 9819
rect 3342 9794 3366 9796
rect 3422 9794 3446 9796
rect 3502 9794 3526 9796
rect 3364 9742 3366 9794
rect 3428 9742 3440 9794
rect 3502 9742 3504 9794
rect 3342 9740 3366 9742
rect 3422 9740 3446 9742
rect 3502 9740 3526 9742
rect 3286 9717 3582 9740
rect 7852 9796 8148 9819
rect 7908 9794 7932 9796
rect 7988 9794 8012 9796
rect 8068 9794 8092 9796
rect 7930 9742 7932 9794
rect 7994 9742 8006 9794
rect 8068 9742 8070 9794
rect 7908 9740 7932 9742
rect 7988 9740 8012 9742
rect 8068 9740 8092 9742
rect 7852 9717 8148 9740
rect 12417 9796 12713 9819
rect 12473 9794 12497 9796
rect 12553 9794 12577 9796
rect 12633 9794 12657 9796
rect 12495 9742 12497 9794
rect 12559 9742 12571 9794
rect 12633 9742 12635 9794
rect 12473 9740 12497 9742
rect 12553 9740 12577 9742
rect 12633 9740 12657 9742
rect 12417 9717 12713 9740
rect 5569 8982 5865 9005
rect 5625 8980 5649 8982
rect 5705 8980 5729 8982
rect 5785 8980 5809 8982
rect 5647 8928 5649 8980
rect 5711 8928 5723 8980
rect 5785 8928 5787 8980
rect 5625 8926 5649 8928
rect 5705 8926 5729 8928
rect 5785 8926 5809 8928
rect 5569 8903 5865 8926
rect 10134 8982 10430 9005
rect 10190 8980 10214 8982
rect 10270 8980 10294 8982
rect 10350 8980 10374 8982
rect 10212 8928 10214 8980
rect 10276 8928 10288 8980
rect 10350 8928 10352 8980
rect 10190 8926 10214 8928
rect 10270 8926 10294 8928
rect 10350 8926 10374 8928
rect 10134 8903 10430 8926
rect 12898 8653 12926 16613
rect 14036 10018 14092 10027
rect 14036 9953 14092 9962
rect 12886 8647 12938 8653
rect 12886 8589 12938 8595
rect 13366 8647 13418 8653
rect 13366 8589 13418 8595
rect 3286 8168 3582 8191
rect 3342 8166 3366 8168
rect 3422 8166 3446 8168
rect 3502 8166 3526 8168
rect 3364 8114 3366 8166
rect 3428 8114 3440 8166
rect 3502 8114 3504 8166
rect 3342 8112 3366 8114
rect 3422 8112 3446 8114
rect 3502 8112 3526 8114
rect 3286 8089 3582 8112
rect 7852 8168 8148 8191
rect 7908 8166 7932 8168
rect 7988 8166 8012 8168
rect 8068 8166 8092 8168
rect 7930 8114 7932 8166
rect 7994 8114 8006 8166
rect 8068 8114 8070 8166
rect 7908 8112 7932 8114
rect 7988 8112 8012 8114
rect 8068 8112 8092 8114
rect 7852 8089 8148 8112
rect 12417 8168 12713 8191
rect 12473 8166 12497 8168
rect 12553 8166 12577 8168
rect 12633 8166 12657 8168
rect 12495 8114 12497 8166
rect 12559 8114 12571 8166
rect 12633 8114 12635 8166
rect 12473 8112 12497 8114
rect 12553 8112 12577 8114
rect 12633 8112 12657 8114
rect 12417 8089 12713 8112
rect 13378 7987 13406 8589
rect 13366 7981 13418 7987
rect 13366 7923 13418 7929
rect 12022 7685 12074 7691
rect 12022 7627 12074 7633
rect 13174 7685 13226 7691
rect 13174 7627 13226 7633
rect 5569 7354 5865 7377
rect 5625 7352 5649 7354
rect 5705 7352 5729 7354
rect 5785 7352 5809 7354
rect 5647 7300 5649 7352
rect 5711 7300 5723 7352
rect 5785 7300 5787 7352
rect 5625 7298 5649 7300
rect 5705 7298 5729 7300
rect 5785 7298 5809 7300
rect 5569 7275 5865 7298
rect 10134 7354 10430 7377
rect 10190 7352 10214 7354
rect 10270 7352 10294 7354
rect 10350 7352 10374 7354
rect 10212 7300 10214 7352
rect 10276 7300 10288 7352
rect 10350 7300 10352 7352
rect 10190 7298 10214 7300
rect 10270 7298 10294 7300
rect 10350 7298 10374 7300
rect 10134 7275 10430 7298
rect 12034 7099 12062 7627
rect 12022 7093 12074 7099
rect 12022 7035 12074 7041
rect 12310 7019 12362 7025
rect 12310 6961 12362 6967
rect 3286 6540 3582 6563
rect 3342 6538 3366 6540
rect 3422 6538 3446 6540
rect 3502 6538 3526 6540
rect 3364 6486 3366 6538
rect 3428 6486 3440 6538
rect 3502 6486 3504 6538
rect 3342 6484 3366 6486
rect 3422 6484 3446 6486
rect 3502 6484 3526 6486
rect 3286 6461 3582 6484
rect 7852 6540 8148 6563
rect 7908 6538 7932 6540
rect 7988 6538 8012 6540
rect 8068 6538 8092 6540
rect 7930 6486 7932 6538
rect 7994 6486 8006 6538
rect 8068 6486 8070 6538
rect 7908 6484 7932 6486
rect 7988 6484 8012 6486
rect 8068 6484 8092 6486
rect 7852 6461 8148 6484
rect 11830 6057 11882 6063
rect 11830 5999 11882 6005
rect 11062 5909 11114 5915
rect 11062 5851 11114 5857
rect 5569 5726 5865 5749
rect 5625 5724 5649 5726
rect 5705 5724 5729 5726
rect 5785 5724 5809 5726
rect 5647 5672 5649 5724
rect 5711 5672 5723 5724
rect 5785 5672 5787 5724
rect 5625 5670 5649 5672
rect 5705 5670 5729 5672
rect 5785 5670 5809 5672
rect 5569 5647 5865 5670
rect 10134 5726 10430 5749
rect 10190 5724 10214 5726
rect 10270 5724 10294 5726
rect 10350 5724 10374 5726
rect 10212 5672 10214 5724
rect 10276 5672 10288 5724
rect 10350 5672 10352 5724
rect 10190 5670 10214 5672
rect 10270 5670 10294 5672
rect 10350 5670 10374 5672
rect 10134 5647 10430 5670
rect 11074 5397 11102 5851
rect 11842 5397 11870 5999
rect 12322 5564 12350 6961
rect 12886 6945 12938 6951
rect 12886 6887 12938 6893
rect 12417 6540 12713 6563
rect 12473 6538 12497 6540
rect 12553 6538 12577 6540
rect 12633 6538 12657 6540
rect 12495 6486 12497 6538
rect 12559 6486 12571 6538
rect 12633 6486 12635 6538
rect 12473 6484 12497 6486
rect 12553 6484 12577 6486
rect 12633 6484 12657 6486
rect 12417 6461 12713 6484
rect 12898 6359 12926 6887
rect 13186 6359 13214 7627
rect 13270 7537 13322 7543
rect 13270 7479 13322 7485
rect 13282 6951 13310 7479
rect 13378 7173 13406 7923
rect 13366 7167 13418 7173
rect 13366 7109 13418 7115
rect 13270 6945 13322 6951
rect 13270 6887 13322 6893
rect 13366 6871 13418 6877
rect 13366 6813 13418 6819
rect 12886 6353 12938 6359
rect 12886 6295 12938 6301
rect 13174 6353 13226 6359
rect 13174 6295 13226 6301
rect 12982 6131 13034 6137
rect 12982 6073 13034 6079
rect 12886 6057 12938 6063
rect 12886 5999 12938 6005
rect 12322 5545 12446 5564
rect 12322 5539 12458 5545
rect 12322 5536 12406 5539
rect 12214 5465 12266 5471
rect 12214 5407 12266 5413
rect 10678 5391 10730 5397
rect 10678 5333 10730 5339
rect 11062 5391 11114 5397
rect 11062 5333 11114 5339
rect 11830 5391 11882 5397
rect 11830 5333 11882 5339
rect 10690 5101 10718 5333
rect 10678 5095 10730 5101
rect 10678 5037 10730 5043
rect 3286 4912 3582 4935
rect 3342 4910 3366 4912
rect 3422 4910 3446 4912
rect 3502 4910 3526 4912
rect 3364 4858 3366 4910
rect 3428 4858 3440 4910
rect 3502 4858 3504 4910
rect 3342 4856 3366 4858
rect 3422 4856 3446 4858
rect 3502 4856 3526 4858
rect 3286 4833 3582 4856
rect 7852 4912 8148 4935
rect 7908 4910 7932 4912
rect 7988 4910 8012 4912
rect 8068 4910 8092 4912
rect 7930 4858 7932 4910
rect 7994 4858 8006 4910
rect 8068 4858 8070 4910
rect 7908 4856 7932 4858
rect 7988 4856 8012 4858
rect 8068 4856 8092 4858
rect 7852 4833 8148 4856
rect 10690 4287 10718 5037
rect 11842 4731 11870 5333
rect 12226 5101 12254 5407
rect 12214 5095 12266 5101
rect 12214 5037 12266 5043
rect 11830 4725 11882 4731
rect 11830 4667 11882 4673
rect 12322 4435 12350 5536
rect 12406 5481 12458 5487
rect 12502 5465 12554 5471
rect 12502 5407 12554 5413
rect 12514 5249 12542 5407
rect 12898 5323 12926 5999
rect 12886 5317 12938 5323
rect 12886 5259 12938 5265
rect 12502 5243 12554 5249
rect 12502 5185 12554 5191
rect 12886 5095 12938 5101
rect 12886 5037 12938 5043
rect 12417 4912 12713 4935
rect 12473 4910 12497 4912
rect 12553 4910 12577 4912
rect 12633 4910 12657 4912
rect 12495 4858 12497 4910
rect 12559 4858 12571 4910
rect 12633 4858 12635 4910
rect 12473 4856 12497 4858
rect 12553 4856 12577 4858
rect 12633 4856 12657 4858
rect 12417 4833 12713 4856
rect 12310 4429 12362 4435
rect 12310 4371 12362 4377
rect 8182 4281 8234 4287
rect 8182 4223 8234 4229
rect 10678 4281 10730 4287
rect 10678 4223 10730 4229
rect 5569 4098 5865 4121
rect 5625 4096 5649 4098
rect 5705 4096 5729 4098
rect 5785 4096 5809 4098
rect 5647 4044 5649 4096
rect 5711 4044 5723 4096
rect 5785 4044 5787 4096
rect 5625 4042 5649 4044
rect 5705 4042 5729 4044
rect 5785 4042 5809 4044
rect 5569 4019 5865 4042
rect 3286 3284 3582 3307
rect 3342 3282 3366 3284
rect 3422 3282 3446 3284
rect 3502 3282 3526 3284
rect 3364 3230 3366 3282
rect 3428 3230 3440 3282
rect 3502 3230 3504 3282
rect 3342 3228 3366 3230
rect 3422 3228 3446 3230
rect 3502 3228 3526 3230
rect 3286 3205 3582 3228
rect 7852 3284 8148 3307
rect 7908 3282 7932 3284
rect 7988 3282 8012 3284
rect 8068 3282 8092 3284
rect 7930 3230 7932 3282
rect 7994 3230 8006 3282
rect 8068 3230 8070 3282
rect 7908 3228 7932 3230
rect 7988 3228 8012 3230
rect 8068 3228 8092 3230
rect 7852 3205 8148 3228
rect 8194 3048 8222 4223
rect 10134 4098 10430 4121
rect 10190 4096 10214 4098
rect 10270 4096 10294 4098
rect 10350 4096 10374 4098
rect 10212 4044 10214 4096
rect 10276 4044 10288 4096
rect 10350 4044 10352 4096
rect 10190 4042 10214 4044
rect 10270 4042 10294 4044
rect 10350 4042 10374 4044
rect 10134 4019 10430 4042
rect 12898 3473 12926 5037
rect 12994 4731 13022 6073
rect 13186 5323 13214 6295
rect 13378 6137 13406 6813
rect 14050 6359 14078 9953
rect 14038 6353 14090 6359
rect 14038 6295 14090 6301
rect 13366 6131 13418 6137
rect 13366 6073 13418 6079
rect 13378 5545 13406 6073
rect 13366 5539 13418 5545
rect 13366 5481 13418 5487
rect 13174 5317 13226 5323
rect 13174 5259 13226 5265
rect 12982 4725 13034 4731
rect 12982 4667 13034 4673
rect 12994 4361 13022 4667
rect 12982 4355 13034 4361
rect 12982 4297 13034 4303
rect 12886 3467 12938 3473
rect 12886 3409 12938 3415
rect 12898 3367 12926 3409
rect 12884 3358 12940 3367
rect 12417 3284 12713 3307
rect 12884 3293 12940 3302
rect 12473 3282 12497 3284
rect 12553 3282 12577 3284
rect 12633 3282 12657 3284
rect 12495 3230 12497 3282
rect 12559 3230 12571 3282
rect 12633 3230 12635 3282
rect 12473 3228 12497 3230
rect 12553 3228 12577 3230
rect 12633 3228 12657 3230
rect 12417 3205 12713 3228
rect 8002 3020 8222 3048
rect 8002 800 8030 3020
rect 7988 0 8044 800
<< via2 >>
rect 12884 16622 12940 16678
rect 3286 16306 3342 16308
rect 3366 16306 3422 16308
rect 3446 16306 3502 16308
rect 3526 16306 3582 16308
rect 3286 16254 3312 16306
rect 3312 16254 3342 16306
rect 3366 16254 3376 16306
rect 3376 16254 3422 16306
rect 3446 16254 3492 16306
rect 3492 16254 3502 16306
rect 3526 16254 3556 16306
rect 3556 16254 3582 16306
rect 3286 16252 3342 16254
rect 3366 16252 3422 16254
rect 3446 16252 3502 16254
rect 3526 16252 3582 16254
rect 7852 16306 7908 16308
rect 7932 16306 7988 16308
rect 8012 16306 8068 16308
rect 8092 16306 8148 16308
rect 7852 16254 7878 16306
rect 7878 16254 7908 16306
rect 7932 16254 7942 16306
rect 7942 16254 7988 16306
rect 8012 16254 8058 16306
rect 8058 16254 8068 16306
rect 8092 16254 8122 16306
rect 8122 16254 8148 16306
rect 7852 16252 7908 16254
rect 7932 16252 7988 16254
rect 8012 16252 8068 16254
rect 8092 16252 8148 16254
rect 12417 16306 12473 16308
rect 12497 16306 12553 16308
rect 12577 16306 12633 16308
rect 12657 16306 12713 16308
rect 12417 16254 12443 16306
rect 12443 16254 12473 16306
rect 12497 16254 12507 16306
rect 12507 16254 12553 16306
rect 12577 16254 12623 16306
rect 12623 16254 12633 16306
rect 12657 16254 12687 16306
rect 12687 16254 12713 16306
rect 12417 16252 12473 16254
rect 12497 16252 12553 16254
rect 12577 16252 12633 16254
rect 12657 16252 12713 16254
rect 5569 15492 5625 15494
rect 5649 15492 5705 15494
rect 5729 15492 5785 15494
rect 5809 15492 5865 15494
rect 5569 15440 5595 15492
rect 5595 15440 5625 15492
rect 5649 15440 5659 15492
rect 5659 15440 5705 15492
rect 5729 15440 5775 15492
rect 5775 15440 5785 15492
rect 5809 15440 5839 15492
rect 5839 15440 5865 15492
rect 5569 15438 5625 15440
rect 5649 15438 5705 15440
rect 5729 15438 5785 15440
rect 5809 15438 5865 15440
rect 10134 15492 10190 15494
rect 10214 15492 10270 15494
rect 10294 15492 10350 15494
rect 10374 15492 10430 15494
rect 10134 15440 10160 15492
rect 10160 15440 10190 15492
rect 10214 15440 10224 15492
rect 10224 15440 10270 15492
rect 10294 15440 10340 15492
rect 10340 15440 10350 15492
rect 10374 15440 10404 15492
rect 10404 15440 10430 15492
rect 10134 15438 10190 15440
rect 10214 15438 10270 15440
rect 10294 15438 10350 15440
rect 10374 15438 10430 15440
rect 3286 14678 3342 14680
rect 3366 14678 3422 14680
rect 3446 14678 3502 14680
rect 3526 14678 3582 14680
rect 3286 14626 3312 14678
rect 3312 14626 3342 14678
rect 3366 14626 3376 14678
rect 3376 14626 3422 14678
rect 3446 14626 3492 14678
rect 3492 14626 3502 14678
rect 3526 14626 3556 14678
rect 3556 14626 3582 14678
rect 3286 14624 3342 14626
rect 3366 14624 3422 14626
rect 3446 14624 3502 14626
rect 3526 14624 3582 14626
rect 7852 14678 7908 14680
rect 7932 14678 7988 14680
rect 8012 14678 8068 14680
rect 8092 14678 8148 14680
rect 7852 14626 7878 14678
rect 7878 14626 7908 14678
rect 7932 14626 7942 14678
rect 7942 14626 7988 14678
rect 8012 14626 8058 14678
rect 8058 14626 8068 14678
rect 8092 14626 8122 14678
rect 8122 14626 8148 14678
rect 7852 14624 7908 14626
rect 7932 14624 7988 14626
rect 8012 14624 8068 14626
rect 8092 14624 8148 14626
rect 12417 14678 12473 14680
rect 12497 14678 12553 14680
rect 12577 14678 12633 14680
rect 12657 14678 12713 14680
rect 12417 14626 12443 14678
rect 12443 14626 12473 14678
rect 12497 14626 12507 14678
rect 12507 14626 12553 14678
rect 12577 14626 12623 14678
rect 12623 14626 12633 14678
rect 12657 14626 12687 14678
rect 12687 14626 12713 14678
rect 12417 14624 12473 14626
rect 12497 14624 12553 14626
rect 12577 14624 12633 14626
rect 12657 14624 12713 14626
rect 5569 13864 5625 13866
rect 5649 13864 5705 13866
rect 5729 13864 5785 13866
rect 5809 13864 5865 13866
rect 5569 13812 5595 13864
rect 5595 13812 5625 13864
rect 5649 13812 5659 13864
rect 5659 13812 5705 13864
rect 5729 13812 5775 13864
rect 5775 13812 5785 13864
rect 5809 13812 5839 13864
rect 5839 13812 5865 13864
rect 5569 13810 5625 13812
rect 5649 13810 5705 13812
rect 5729 13810 5785 13812
rect 5809 13810 5865 13812
rect 10134 13864 10190 13866
rect 10214 13864 10270 13866
rect 10294 13864 10350 13866
rect 10374 13864 10430 13866
rect 10134 13812 10160 13864
rect 10160 13812 10190 13864
rect 10214 13812 10224 13864
rect 10224 13812 10270 13864
rect 10294 13812 10340 13864
rect 10340 13812 10350 13864
rect 10374 13812 10404 13864
rect 10404 13812 10430 13864
rect 10134 13810 10190 13812
rect 10214 13810 10270 13812
rect 10294 13810 10350 13812
rect 10374 13810 10430 13812
rect 3286 13050 3342 13052
rect 3366 13050 3422 13052
rect 3446 13050 3502 13052
rect 3526 13050 3582 13052
rect 3286 12998 3312 13050
rect 3312 12998 3342 13050
rect 3366 12998 3376 13050
rect 3376 12998 3422 13050
rect 3446 12998 3492 13050
rect 3492 12998 3502 13050
rect 3526 12998 3556 13050
rect 3556 12998 3582 13050
rect 3286 12996 3342 12998
rect 3366 12996 3422 12998
rect 3446 12996 3502 12998
rect 3526 12996 3582 12998
rect 7852 13050 7908 13052
rect 7932 13050 7988 13052
rect 8012 13050 8068 13052
rect 8092 13050 8148 13052
rect 7852 12998 7878 13050
rect 7878 12998 7908 13050
rect 7932 12998 7942 13050
rect 7942 12998 7988 13050
rect 8012 12998 8058 13050
rect 8058 12998 8068 13050
rect 8092 12998 8122 13050
rect 8122 12998 8148 13050
rect 7852 12996 7908 12998
rect 7932 12996 7988 12998
rect 8012 12996 8068 12998
rect 8092 12996 8148 12998
rect 12417 13050 12473 13052
rect 12497 13050 12553 13052
rect 12577 13050 12633 13052
rect 12657 13050 12713 13052
rect 12417 12998 12443 13050
rect 12443 12998 12473 13050
rect 12497 12998 12507 13050
rect 12507 12998 12553 13050
rect 12577 12998 12623 13050
rect 12623 12998 12633 13050
rect 12657 12998 12687 13050
rect 12687 12998 12713 13050
rect 12417 12996 12473 12998
rect 12497 12996 12553 12998
rect 12577 12996 12633 12998
rect 12657 12996 12713 12998
rect 5569 12236 5625 12238
rect 5649 12236 5705 12238
rect 5729 12236 5785 12238
rect 5809 12236 5865 12238
rect 5569 12184 5595 12236
rect 5595 12184 5625 12236
rect 5649 12184 5659 12236
rect 5659 12184 5705 12236
rect 5729 12184 5775 12236
rect 5775 12184 5785 12236
rect 5809 12184 5839 12236
rect 5839 12184 5865 12236
rect 5569 12182 5625 12184
rect 5649 12182 5705 12184
rect 5729 12182 5785 12184
rect 5809 12182 5865 12184
rect 10134 12236 10190 12238
rect 10214 12236 10270 12238
rect 10294 12236 10350 12238
rect 10374 12236 10430 12238
rect 10134 12184 10160 12236
rect 10160 12184 10190 12236
rect 10214 12184 10224 12236
rect 10224 12184 10270 12236
rect 10294 12184 10340 12236
rect 10340 12184 10350 12236
rect 10374 12184 10404 12236
rect 10404 12184 10430 12236
rect 10134 12182 10190 12184
rect 10214 12182 10270 12184
rect 10294 12182 10350 12184
rect 10374 12182 10430 12184
rect 3286 11422 3342 11424
rect 3366 11422 3422 11424
rect 3446 11422 3502 11424
rect 3526 11422 3582 11424
rect 3286 11370 3312 11422
rect 3312 11370 3342 11422
rect 3366 11370 3376 11422
rect 3376 11370 3422 11422
rect 3446 11370 3492 11422
rect 3492 11370 3502 11422
rect 3526 11370 3556 11422
rect 3556 11370 3582 11422
rect 3286 11368 3342 11370
rect 3366 11368 3422 11370
rect 3446 11368 3502 11370
rect 3526 11368 3582 11370
rect 7852 11422 7908 11424
rect 7932 11422 7988 11424
rect 8012 11422 8068 11424
rect 8092 11422 8148 11424
rect 7852 11370 7878 11422
rect 7878 11370 7908 11422
rect 7932 11370 7942 11422
rect 7942 11370 7988 11422
rect 8012 11370 8058 11422
rect 8058 11370 8068 11422
rect 8092 11370 8122 11422
rect 8122 11370 8148 11422
rect 7852 11368 7908 11370
rect 7932 11368 7988 11370
rect 8012 11368 8068 11370
rect 8092 11368 8148 11370
rect 12417 11422 12473 11424
rect 12497 11422 12553 11424
rect 12577 11422 12633 11424
rect 12657 11422 12713 11424
rect 12417 11370 12443 11422
rect 12443 11370 12473 11422
rect 12497 11370 12507 11422
rect 12507 11370 12553 11422
rect 12577 11370 12623 11422
rect 12623 11370 12633 11422
rect 12657 11370 12687 11422
rect 12687 11370 12713 11422
rect 12417 11368 12473 11370
rect 12497 11368 12553 11370
rect 12577 11368 12633 11370
rect 12657 11368 12713 11370
rect 5569 10608 5625 10610
rect 5649 10608 5705 10610
rect 5729 10608 5785 10610
rect 5809 10608 5865 10610
rect 5569 10556 5595 10608
rect 5595 10556 5625 10608
rect 5649 10556 5659 10608
rect 5659 10556 5705 10608
rect 5729 10556 5775 10608
rect 5775 10556 5785 10608
rect 5809 10556 5839 10608
rect 5839 10556 5865 10608
rect 5569 10554 5625 10556
rect 5649 10554 5705 10556
rect 5729 10554 5785 10556
rect 5809 10554 5865 10556
rect 10134 10608 10190 10610
rect 10214 10608 10270 10610
rect 10294 10608 10350 10610
rect 10374 10608 10430 10610
rect 10134 10556 10160 10608
rect 10160 10556 10190 10608
rect 10214 10556 10224 10608
rect 10224 10556 10270 10608
rect 10294 10556 10340 10608
rect 10340 10556 10350 10608
rect 10374 10556 10404 10608
rect 10404 10556 10430 10608
rect 10134 10554 10190 10556
rect 10214 10554 10270 10556
rect 10294 10554 10350 10556
rect 10374 10554 10430 10556
rect 3286 9794 3342 9796
rect 3366 9794 3422 9796
rect 3446 9794 3502 9796
rect 3526 9794 3582 9796
rect 3286 9742 3312 9794
rect 3312 9742 3342 9794
rect 3366 9742 3376 9794
rect 3376 9742 3422 9794
rect 3446 9742 3492 9794
rect 3492 9742 3502 9794
rect 3526 9742 3556 9794
rect 3556 9742 3582 9794
rect 3286 9740 3342 9742
rect 3366 9740 3422 9742
rect 3446 9740 3502 9742
rect 3526 9740 3582 9742
rect 7852 9794 7908 9796
rect 7932 9794 7988 9796
rect 8012 9794 8068 9796
rect 8092 9794 8148 9796
rect 7852 9742 7878 9794
rect 7878 9742 7908 9794
rect 7932 9742 7942 9794
rect 7942 9742 7988 9794
rect 8012 9742 8058 9794
rect 8058 9742 8068 9794
rect 8092 9742 8122 9794
rect 8122 9742 8148 9794
rect 7852 9740 7908 9742
rect 7932 9740 7988 9742
rect 8012 9740 8068 9742
rect 8092 9740 8148 9742
rect 12417 9794 12473 9796
rect 12497 9794 12553 9796
rect 12577 9794 12633 9796
rect 12657 9794 12713 9796
rect 12417 9742 12443 9794
rect 12443 9742 12473 9794
rect 12497 9742 12507 9794
rect 12507 9742 12553 9794
rect 12577 9742 12623 9794
rect 12623 9742 12633 9794
rect 12657 9742 12687 9794
rect 12687 9742 12713 9794
rect 12417 9740 12473 9742
rect 12497 9740 12553 9742
rect 12577 9740 12633 9742
rect 12657 9740 12713 9742
rect 5569 8980 5625 8982
rect 5649 8980 5705 8982
rect 5729 8980 5785 8982
rect 5809 8980 5865 8982
rect 5569 8928 5595 8980
rect 5595 8928 5625 8980
rect 5649 8928 5659 8980
rect 5659 8928 5705 8980
rect 5729 8928 5775 8980
rect 5775 8928 5785 8980
rect 5809 8928 5839 8980
rect 5839 8928 5865 8980
rect 5569 8926 5625 8928
rect 5649 8926 5705 8928
rect 5729 8926 5785 8928
rect 5809 8926 5865 8928
rect 10134 8980 10190 8982
rect 10214 8980 10270 8982
rect 10294 8980 10350 8982
rect 10374 8980 10430 8982
rect 10134 8928 10160 8980
rect 10160 8928 10190 8980
rect 10214 8928 10224 8980
rect 10224 8928 10270 8980
rect 10294 8928 10340 8980
rect 10340 8928 10350 8980
rect 10374 8928 10404 8980
rect 10404 8928 10430 8980
rect 10134 8926 10190 8928
rect 10214 8926 10270 8928
rect 10294 8926 10350 8928
rect 10374 8926 10430 8928
rect 14036 9962 14092 10018
rect 3286 8166 3342 8168
rect 3366 8166 3422 8168
rect 3446 8166 3502 8168
rect 3526 8166 3582 8168
rect 3286 8114 3312 8166
rect 3312 8114 3342 8166
rect 3366 8114 3376 8166
rect 3376 8114 3422 8166
rect 3446 8114 3492 8166
rect 3492 8114 3502 8166
rect 3526 8114 3556 8166
rect 3556 8114 3582 8166
rect 3286 8112 3342 8114
rect 3366 8112 3422 8114
rect 3446 8112 3502 8114
rect 3526 8112 3582 8114
rect 7852 8166 7908 8168
rect 7932 8166 7988 8168
rect 8012 8166 8068 8168
rect 8092 8166 8148 8168
rect 7852 8114 7878 8166
rect 7878 8114 7908 8166
rect 7932 8114 7942 8166
rect 7942 8114 7988 8166
rect 8012 8114 8058 8166
rect 8058 8114 8068 8166
rect 8092 8114 8122 8166
rect 8122 8114 8148 8166
rect 7852 8112 7908 8114
rect 7932 8112 7988 8114
rect 8012 8112 8068 8114
rect 8092 8112 8148 8114
rect 12417 8166 12473 8168
rect 12497 8166 12553 8168
rect 12577 8166 12633 8168
rect 12657 8166 12713 8168
rect 12417 8114 12443 8166
rect 12443 8114 12473 8166
rect 12497 8114 12507 8166
rect 12507 8114 12553 8166
rect 12577 8114 12623 8166
rect 12623 8114 12633 8166
rect 12657 8114 12687 8166
rect 12687 8114 12713 8166
rect 12417 8112 12473 8114
rect 12497 8112 12553 8114
rect 12577 8112 12633 8114
rect 12657 8112 12713 8114
rect 5569 7352 5625 7354
rect 5649 7352 5705 7354
rect 5729 7352 5785 7354
rect 5809 7352 5865 7354
rect 5569 7300 5595 7352
rect 5595 7300 5625 7352
rect 5649 7300 5659 7352
rect 5659 7300 5705 7352
rect 5729 7300 5775 7352
rect 5775 7300 5785 7352
rect 5809 7300 5839 7352
rect 5839 7300 5865 7352
rect 5569 7298 5625 7300
rect 5649 7298 5705 7300
rect 5729 7298 5785 7300
rect 5809 7298 5865 7300
rect 10134 7352 10190 7354
rect 10214 7352 10270 7354
rect 10294 7352 10350 7354
rect 10374 7352 10430 7354
rect 10134 7300 10160 7352
rect 10160 7300 10190 7352
rect 10214 7300 10224 7352
rect 10224 7300 10270 7352
rect 10294 7300 10340 7352
rect 10340 7300 10350 7352
rect 10374 7300 10404 7352
rect 10404 7300 10430 7352
rect 10134 7298 10190 7300
rect 10214 7298 10270 7300
rect 10294 7298 10350 7300
rect 10374 7298 10430 7300
rect 3286 6538 3342 6540
rect 3366 6538 3422 6540
rect 3446 6538 3502 6540
rect 3526 6538 3582 6540
rect 3286 6486 3312 6538
rect 3312 6486 3342 6538
rect 3366 6486 3376 6538
rect 3376 6486 3422 6538
rect 3446 6486 3492 6538
rect 3492 6486 3502 6538
rect 3526 6486 3556 6538
rect 3556 6486 3582 6538
rect 3286 6484 3342 6486
rect 3366 6484 3422 6486
rect 3446 6484 3502 6486
rect 3526 6484 3582 6486
rect 7852 6538 7908 6540
rect 7932 6538 7988 6540
rect 8012 6538 8068 6540
rect 8092 6538 8148 6540
rect 7852 6486 7878 6538
rect 7878 6486 7908 6538
rect 7932 6486 7942 6538
rect 7942 6486 7988 6538
rect 8012 6486 8058 6538
rect 8058 6486 8068 6538
rect 8092 6486 8122 6538
rect 8122 6486 8148 6538
rect 7852 6484 7908 6486
rect 7932 6484 7988 6486
rect 8012 6484 8068 6486
rect 8092 6484 8148 6486
rect 5569 5724 5625 5726
rect 5649 5724 5705 5726
rect 5729 5724 5785 5726
rect 5809 5724 5865 5726
rect 5569 5672 5595 5724
rect 5595 5672 5625 5724
rect 5649 5672 5659 5724
rect 5659 5672 5705 5724
rect 5729 5672 5775 5724
rect 5775 5672 5785 5724
rect 5809 5672 5839 5724
rect 5839 5672 5865 5724
rect 5569 5670 5625 5672
rect 5649 5670 5705 5672
rect 5729 5670 5785 5672
rect 5809 5670 5865 5672
rect 10134 5724 10190 5726
rect 10214 5724 10270 5726
rect 10294 5724 10350 5726
rect 10374 5724 10430 5726
rect 10134 5672 10160 5724
rect 10160 5672 10190 5724
rect 10214 5672 10224 5724
rect 10224 5672 10270 5724
rect 10294 5672 10340 5724
rect 10340 5672 10350 5724
rect 10374 5672 10404 5724
rect 10404 5672 10430 5724
rect 10134 5670 10190 5672
rect 10214 5670 10270 5672
rect 10294 5670 10350 5672
rect 10374 5670 10430 5672
rect 12417 6538 12473 6540
rect 12497 6538 12553 6540
rect 12577 6538 12633 6540
rect 12657 6538 12713 6540
rect 12417 6486 12443 6538
rect 12443 6486 12473 6538
rect 12497 6486 12507 6538
rect 12507 6486 12553 6538
rect 12577 6486 12623 6538
rect 12623 6486 12633 6538
rect 12657 6486 12687 6538
rect 12687 6486 12713 6538
rect 12417 6484 12473 6486
rect 12497 6484 12553 6486
rect 12577 6484 12633 6486
rect 12657 6484 12713 6486
rect 3286 4910 3342 4912
rect 3366 4910 3422 4912
rect 3446 4910 3502 4912
rect 3526 4910 3582 4912
rect 3286 4858 3312 4910
rect 3312 4858 3342 4910
rect 3366 4858 3376 4910
rect 3376 4858 3422 4910
rect 3446 4858 3492 4910
rect 3492 4858 3502 4910
rect 3526 4858 3556 4910
rect 3556 4858 3582 4910
rect 3286 4856 3342 4858
rect 3366 4856 3422 4858
rect 3446 4856 3502 4858
rect 3526 4856 3582 4858
rect 7852 4910 7908 4912
rect 7932 4910 7988 4912
rect 8012 4910 8068 4912
rect 8092 4910 8148 4912
rect 7852 4858 7878 4910
rect 7878 4858 7908 4910
rect 7932 4858 7942 4910
rect 7942 4858 7988 4910
rect 8012 4858 8058 4910
rect 8058 4858 8068 4910
rect 8092 4858 8122 4910
rect 8122 4858 8148 4910
rect 7852 4856 7908 4858
rect 7932 4856 7988 4858
rect 8012 4856 8068 4858
rect 8092 4856 8148 4858
rect 12417 4910 12473 4912
rect 12497 4910 12553 4912
rect 12577 4910 12633 4912
rect 12657 4910 12713 4912
rect 12417 4858 12443 4910
rect 12443 4858 12473 4910
rect 12497 4858 12507 4910
rect 12507 4858 12553 4910
rect 12577 4858 12623 4910
rect 12623 4858 12633 4910
rect 12657 4858 12687 4910
rect 12687 4858 12713 4910
rect 12417 4856 12473 4858
rect 12497 4856 12553 4858
rect 12577 4856 12633 4858
rect 12657 4856 12713 4858
rect 5569 4096 5625 4098
rect 5649 4096 5705 4098
rect 5729 4096 5785 4098
rect 5809 4096 5865 4098
rect 5569 4044 5595 4096
rect 5595 4044 5625 4096
rect 5649 4044 5659 4096
rect 5659 4044 5705 4096
rect 5729 4044 5775 4096
rect 5775 4044 5785 4096
rect 5809 4044 5839 4096
rect 5839 4044 5865 4096
rect 5569 4042 5625 4044
rect 5649 4042 5705 4044
rect 5729 4042 5785 4044
rect 5809 4042 5865 4044
rect 3286 3282 3342 3284
rect 3366 3282 3422 3284
rect 3446 3282 3502 3284
rect 3526 3282 3582 3284
rect 3286 3230 3312 3282
rect 3312 3230 3342 3282
rect 3366 3230 3376 3282
rect 3376 3230 3422 3282
rect 3446 3230 3492 3282
rect 3492 3230 3502 3282
rect 3526 3230 3556 3282
rect 3556 3230 3582 3282
rect 3286 3228 3342 3230
rect 3366 3228 3422 3230
rect 3446 3228 3502 3230
rect 3526 3228 3582 3230
rect 7852 3282 7908 3284
rect 7932 3282 7988 3284
rect 8012 3282 8068 3284
rect 8092 3282 8148 3284
rect 7852 3230 7878 3282
rect 7878 3230 7908 3282
rect 7932 3230 7942 3282
rect 7942 3230 7988 3282
rect 8012 3230 8058 3282
rect 8058 3230 8068 3282
rect 8092 3230 8122 3282
rect 8122 3230 8148 3282
rect 7852 3228 7908 3230
rect 7932 3228 7988 3230
rect 8012 3228 8068 3230
rect 8092 3228 8148 3230
rect 10134 4096 10190 4098
rect 10214 4096 10270 4098
rect 10294 4096 10350 4098
rect 10374 4096 10430 4098
rect 10134 4044 10160 4096
rect 10160 4044 10190 4096
rect 10214 4044 10224 4096
rect 10224 4044 10270 4096
rect 10294 4044 10340 4096
rect 10340 4044 10350 4096
rect 10374 4044 10404 4096
rect 10404 4044 10430 4096
rect 10134 4042 10190 4044
rect 10214 4042 10270 4044
rect 10294 4042 10350 4044
rect 10374 4042 10430 4044
rect 12884 3302 12940 3358
rect 12417 3282 12473 3284
rect 12497 3282 12553 3284
rect 12577 3282 12633 3284
rect 12657 3282 12713 3284
rect 12417 3230 12443 3282
rect 12443 3230 12473 3282
rect 12497 3230 12507 3282
rect 12507 3230 12553 3282
rect 12577 3230 12623 3282
rect 12623 3230 12633 3282
rect 12657 3230 12687 3282
rect 12687 3230 12713 3282
rect 12417 3228 12473 3230
rect 12497 3228 12553 3230
rect 12577 3228 12633 3230
rect 12657 3228 12713 3230
<< metal3 >>
rect 12879 16680 12945 16683
rect 15200 16680 16000 16710
rect 12879 16678 16000 16680
rect 12879 16622 12884 16678
rect 12940 16622 16000 16678
rect 12879 16620 16000 16622
rect 12879 16617 12945 16620
rect 15200 16590 16000 16620
rect 3274 16312 3594 16313
rect 3274 16248 3282 16312
rect 3346 16248 3362 16312
rect 3426 16248 3442 16312
rect 3506 16248 3522 16312
rect 3586 16248 3594 16312
rect 3274 16247 3594 16248
rect 7840 16312 8160 16313
rect 7840 16248 7848 16312
rect 7912 16248 7928 16312
rect 7992 16248 8008 16312
rect 8072 16248 8088 16312
rect 8152 16248 8160 16312
rect 7840 16247 8160 16248
rect 12405 16312 12725 16313
rect 12405 16248 12413 16312
rect 12477 16248 12493 16312
rect 12557 16248 12573 16312
rect 12637 16248 12653 16312
rect 12717 16248 12725 16312
rect 12405 16247 12725 16248
rect 5557 15498 5877 15499
rect 5557 15434 5565 15498
rect 5629 15434 5645 15498
rect 5709 15434 5725 15498
rect 5789 15434 5805 15498
rect 5869 15434 5877 15498
rect 5557 15433 5877 15434
rect 10122 15498 10442 15499
rect 10122 15434 10130 15498
rect 10194 15434 10210 15498
rect 10274 15434 10290 15498
rect 10354 15434 10370 15498
rect 10434 15434 10442 15498
rect 10122 15433 10442 15434
rect 3274 14684 3594 14685
rect 3274 14620 3282 14684
rect 3346 14620 3362 14684
rect 3426 14620 3442 14684
rect 3506 14620 3522 14684
rect 3586 14620 3594 14684
rect 3274 14619 3594 14620
rect 7840 14684 8160 14685
rect 7840 14620 7848 14684
rect 7912 14620 7928 14684
rect 7992 14620 8008 14684
rect 8072 14620 8088 14684
rect 8152 14620 8160 14684
rect 7840 14619 8160 14620
rect 12405 14684 12725 14685
rect 12405 14620 12413 14684
rect 12477 14620 12493 14684
rect 12557 14620 12573 14684
rect 12637 14620 12653 14684
rect 12717 14620 12725 14684
rect 12405 14619 12725 14620
rect 5557 13870 5877 13871
rect 5557 13806 5565 13870
rect 5629 13806 5645 13870
rect 5709 13806 5725 13870
rect 5789 13806 5805 13870
rect 5869 13806 5877 13870
rect 5557 13805 5877 13806
rect 10122 13870 10442 13871
rect 10122 13806 10130 13870
rect 10194 13806 10210 13870
rect 10274 13806 10290 13870
rect 10354 13806 10370 13870
rect 10434 13806 10442 13870
rect 10122 13805 10442 13806
rect 3274 13056 3594 13057
rect 3274 12992 3282 13056
rect 3346 12992 3362 13056
rect 3426 12992 3442 13056
rect 3506 12992 3522 13056
rect 3586 12992 3594 13056
rect 3274 12991 3594 12992
rect 7840 13056 8160 13057
rect 7840 12992 7848 13056
rect 7912 12992 7928 13056
rect 7992 12992 8008 13056
rect 8072 12992 8088 13056
rect 8152 12992 8160 13056
rect 7840 12991 8160 12992
rect 12405 13056 12725 13057
rect 12405 12992 12413 13056
rect 12477 12992 12493 13056
rect 12557 12992 12573 13056
rect 12637 12992 12653 13056
rect 12717 12992 12725 13056
rect 12405 12991 12725 12992
rect 5557 12242 5877 12243
rect 5557 12178 5565 12242
rect 5629 12178 5645 12242
rect 5709 12178 5725 12242
rect 5789 12178 5805 12242
rect 5869 12178 5877 12242
rect 5557 12177 5877 12178
rect 10122 12242 10442 12243
rect 10122 12178 10130 12242
rect 10194 12178 10210 12242
rect 10274 12178 10290 12242
rect 10354 12178 10370 12242
rect 10434 12178 10442 12242
rect 10122 12177 10442 12178
rect 3274 11428 3594 11429
rect 3274 11364 3282 11428
rect 3346 11364 3362 11428
rect 3426 11364 3442 11428
rect 3506 11364 3522 11428
rect 3586 11364 3594 11428
rect 3274 11363 3594 11364
rect 7840 11428 8160 11429
rect 7840 11364 7848 11428
rect 7912 11364 7928 11428
rect 7992 11364 8008 11428
rect 8072 11364 8088 11428
rect 8152 11364 8160 11428
rect 7840 11363 8160 11364
rect 12405 11428 12725 11429
rect 12405 11364 12413 11428
rect 12477 11364 12493 11428
rect 12557 11364 12573 11428
rect 12637 11364 12653 11428
rect 12717 11364 12725 11428
rect 12405 11363 12725 11364
rect 5557 10614 5877 10615
rect 5557 10550 5565 10614
rect 5629 10550 5645 10614
rect 5709 10550 5725 10614
rect 5789 10550 5805 10614
rect 5869 10550 5877 10614
rect 5557 10549 5877 10550
rect 10122 10614 10442 10615
rect 10122 10550 10130 10614
rect 10194 10550 10210 10614
rect 10274 10550 10290 10614
rect 10354 10550 10370 10614
rect 10434 10550 10442 10614
rect 10122 10549 10442 10550
rect 14031 10020 14097 10023
rect 15200 10020 16000 10050
rect 14031 10018 16000 10020
rect 14031 9962 14036 10018
rect 14092 9962 16000 10018
rect 14031 9960 16000 9962
rect 14031 9957 14097 9960
rect 15200 9930 16000 9960
rect 3274 9800 3594 9801
rect 3274 9736 3282 9800
rect 3346 9736 3362 9800
rect 3426 9736 3442 9800
rect 3506 9736 3522 9800
rect 3586 9736 3594 9800
rect 3274 9735 3594 9736
rect 7840 9800 8160 9801
rect 7840 9736 7848 9800
rect 7912 9736 7928 9800
rect 7992 9736 8008 9800
rect 8072 9736 8088 9800
rect 8152 9736 8160 9800
rect 7840 9735 8160 9736
rect 12405 9800 12725 9801
rect 12405 9736 12413 9800
rect 12477 9736 12493 9800
rect 12557 9736 12573 9800
rect 12637 9736 12653 9800
rect 12717 9736 12725 9800
rect 12405 9735 12725 9736
rect 5557 8986 5877 8987
rect 5557 8922 5565 8986
rect 5629 8922 5645 8986
rect 5709 8922 5725 8986
rect 5789 8922 5805 8986
rect 5869 8922 5877 8986
rect 5557 8921 5877 8922
rect 10122 8986 10442 8987
rect 10122 8922 10130 8986
rect 10194 8922 10210 8986
rect 10274 8922 10290 8986
rect 10354 8922 10370 8986
rect 10434 8922 10442 8986
rect 10122 8921 10442 8922
rect 3274 8172 3594 8173
rect 3274 8108 3282 8172
rect 3346 8108 3362 8172
rect 3426 8108 3442 8172
rect 3506 8108 3522 8172
rect 3586 8108 3594 8172
rect 3274 8107 3594 8108
rect 7840 8172 8160 8173
rect 7840 8108 7848 8172
rect 7912 8108 7928 8172
rect 7992 8108 8008 8172
rect 8072 8108 8088 8172
rect 8152 8108 8160 8172
rect 7840 8107 8160 8108
rect 12405 8172 12725 8173
rect 12405 8108 12413 8172
rect 12477 8108 12493 8172
rect 12557 8108 12573 8172
rect 12637 8108 12653 8172
rect 12717 8108 12725 8172
rect 12405 8107 12725 8108
rect 5557 7358 5877 7359
rect 5557 7294 5565 7358
rect 5629 7294 5645 7358
rect 5709 7294 5725 7358
rect 5789 7294 5805 7358
rect 5869 7294 5877 7358
rect 5557 7293 5877 7294
rect 10122 7358 10442 7359
rect 10122 7294 10130 7358
rect 10194 7294 10210 7358
rect 10274 7294 10290 7358
rect 10354 7294 10370 7358
rect 10434 7294 10442 7358
rect 10122 7293 10442 7294
rect 3274 6544 3594 6545
rect 3274 6480 3282 6544
rect 3346 6480 3362 6544
rect 3426 6480 3442 6544
rect 3506 6480 3522 6544
rect 3586 6480 3594 6544
rect 3274 6479 3594 6480
rect 7840 6544 8160 6545
rect 7840 6480 7848 6544
rect 7912 6480 7928 6544
rect 7992 6480 8008 6544
rect 8072 6480 8088 6544
rect 8152 6480 8160 6544
rect 7840 6479 8160 6480
rect 12405 6544 12725 6545
rect 12405 6480 12413 6544
rect 12477 6480 12493 6544
rect 12557 6480 12573 6544
rect 12637 6480 12653 6544
rect 12717 6480 12725 6544
rect 12405 6479 12725 6480
rect 5557 5730 5877 5731
rect 5557 5666 5565 5730
rect 5629 5666 5645 5730
rect 5709 5666 5725 5730
rect 5789 5666 5805 5730
rect 5869 5666 5877 5730
rect 5557 5665 5877 5666
rect 10122 5730 10442 5731
rect 10122 5666 10130 5730
rect 10194 5666 10210 5730
rect 10274 5666 10290 5730
rect 10354 5666 10370 5730
rect 10434 5666 10442 5730
rect 10122 5665 10442 5666
rect 3274 4916 3594 4917
rect 3274 4852 3282 4916
rect 3346 4852 3362 4916
rect 3426 4852 3442 4916
rect 3506 4852 3522 4916
rect 3586 4852 3594 4916
rect 3274 4851 3594 4852
rect 7840 4916 8160 4917
rect 7840 4852 7848 4916
rect 7912 4852 7928 4916
rect 7992 4852 8008 4916
rect 8072 4852 8088 4916
rect 8152 4852 8160 4916
rect 7840 4851 8160 4852
rect 12405 4916 12725 4917
rect 12405 4852 12413 4916
rect 12477 4852 12493 4916
rect 12557 4852 12573 4916
rect 12637 4852 12653 4916
rect 12717 4852 12725 4916
rect 12405 4851 12725 4852
rect 5557 4102 5877 4103
rect 5557 4038 5565 4102
rect 5629 4038 5645 4102
rect 5709 4038 5725 4102
rect 5789 4038 5805 4102
rect 5869 4038 5877 4102
rect 5557 4037 5877 4038
rect 10122 4102 10442 4103
rect 10122 4038 10130 4102
rect 10194 4038 10210 4102
rect 10274 4038 10290 4102
rect 10354 4038 10370 4102
rect 10434 4038 10442 4102
rect 10122 4037 10442 4038
rect 12879 3360 12945 3363
rect 15200 3360 16000 3390
rect 12879 3358 16000 3360
rect 12879 3302 12884 3358
rect 12940 3302 16000 3358
rect 12879 3300 16000 3302
rect 12879 3297 12945 3300
rect 3274 3288 3594 3289
rect 3274 3224 3282 3288
rect 3346 3224 3362 3288
rect 3426 3224 3442 3288
rect 3506 3224 3522 3288
rect 3586 3224 3594 3288
rect 3274 3223 3594 3224
rect 7840 3288 8160 3289
rect 7840 3224 7848 3288
rect 7912 3224 7928 3288
rect 7992 3224 8008 3288
rect 8072 3224 8088 3288
rect 8152 3224 8160 3288
rect 7840 3223 8160 3224
rect 12405 3288 12725 3289
rect 12405 3224 12413 3288
rect 12477 3224 12493 3288
rect 12557 3224 12573 3288
rect 12637 3224 12653 3288
rect 12717 3224 12725 3288
rect 15200 3270 16000 3300
rect 12405 3223 12725 3224
<< via3 >>
rect 3282 16308 3346 16312
rect 3282 16252 3286 16308
rect 3286 16252 3342 16308
rect 3342 16252 3346 16308
rect 3282 16248 3346 16252
rect 3362 16308 3426 16312
rect 3362 16252 3366 16308
rect 3366 16252 3422 16308
rect 3422 16252 3426 16308
rect 3362 16248 3426 16252
rect 3442 16308 3506 16312
rect 3442 16252 3446 16308
rect 3446 16252 3502 16308
rect 3502 16252 3506 16308
rect 3442 16248 3506 16252
rect 3522 16308 3586 16312
rect 3522 16252 3526 16308
rect 3526 16252 3582 16308
rect 3582 16252 3586 16308
rect 3522 16248 3586 16252
rect 7848 16308 7912 16312
rect 7848 16252 7852 16308
rect 7852 16252 7908 16308
rect 7908 16252 7912 16308
rect 7848 16248 7912 16252
rect 7928 16308 7992 16312
rect 7928 16252 7932 16308
rect 7932 16252 7988 16308
rect 7988 16252 7992 16308
rect 7928 16248 7992 16252
rect 8008 16308 8072 16312
rect 8008 16252 8012 16308
rect 8012 16252 8068 16308
rect 8068 16252 8072 16308
rect 8008 16248 8072 16252
rect 8088 16308 8152 16312
rect 8088 16252 8092 16308
rect 8092 16252 8148 16308
rect 8148 16252 8152 16308
rect 8088 16248 8152 16252
rect 12413 16308 12477 16312
rect 12413 16252 12417 16308
rect 12417 16252 12473 16308
rect 12473 16252 12477 16308
rect 12413 16248 12477 16252
rect 12493 16308 12557 16312
rect 12493 16252 12497 16308
rect 12497 16252 12553 16308
rect 12553 16252 12557 16308
rect 12493 16248 12557 16252
rect 12573 16308 12637 16312
rect 12573 16252 12577 16308
rect 12577 16252 12633 16308
rect 12633 16252 12637 16308
rect 12573 16248 12637 16252
rect 12653 16308 12717 16312
rect 12653 16252 12657 16308
rect 12657 16252 12713 16308
rect 12713 16252 12717 16308
rect 12653 16248 12717 16252
rect 5565 15494 5629 15498
rect 5565 15438 5569 15494
rect 5569 15438 5625 15494
rect 5625 15438 5629 15494
rect 5565 15434 5629 15438
rect 5645 15494 5709 15498
rect 5645 15438 5649 15494
rect 5649 15438 5705 15494
rect 5705 15438 5709 15494
rect 5645 15434 5709 15438
rect 5725 15494 5789 15498
rect 5725 15438 5729 15494
rect 5729 15438 5785 15494
rect 5785 15438 5789 15494
rect 5725 15434 5789 15438
rect 5805 15494 5869 15498
rect 5805 15438 5809 15494
rect 5809 15438 5865 15494
rect 5865 15438 5869 15494
rect 5805 15434 5869 15438
rect 10130 15494 10194 15498
rect 10130 15438 10134 15494
rect 10134 15438 10190 15494
rect 10190 15438 10194 15494
rect 10130 15434 10194 15438
rect 10210 15494 10274 15498
rect 10210 15438 10214 15494
rect 10214 15438 10270 15494
rect 10270 15438 10274 15494
rect 10210 15434 10274 15438
rect 10290 15494 10354 15498
rect 10290 15438 10294 15494
rect 10294 15438 10350 15494
rect 10350 15438 10354 15494
rect 10290 15434 10354 15438
rect 10370 15494 10434 15498
rect 10370 15438 10374 15494
rect 10374 15438 10430 15494
rect 10430 15438 10434 15494
rect 10370 15434 10434 15438
rect 3282 14680 3346 14684
rect 3282 14624 3286 14680
rect 3286 14624 3342 14680
rect 3342 14624 3346 14680
rect 3282 14620 3346 14624
rect 3362 14680 3426 14684
rect 3362 14624 3366 14680
rect 3366 14624 3422 14680
rect 3422 14624 3426 14680
rect 3362 14620 3426 14624
rect 3442 14680 3506 14684
rect 3442 14624 3446 14680
rect 3446 14624 3502 14680
rect 3502 14624 3506 14680
rect 3442 14620 3506 14624
rect 3522 14680 3586 14684
rect 3522 14624 3526 14680
rect 3526 14624 3582 14680
rect 3582 14624 3586 14680
rect 3522 14620 3586 14624
rect 7848 14680 7912 14684
rect 7848 14624 7852 14680
rect 7852 14624 7908 14680
rect 7908 14624 7912 14680
rect 7848 14620 7912 14624
rect 7928 14680 7992 14684
rect 7928 14624 7932 14680
rect 7932 14624 7988 14680
rect 7988 14624 7992 14680
rect 7928 14620 7992 14624
rect 8008 14680 8072 14684
rect 8008 14624 8012 14680
rect 8012 14624 8068 14680
rect 8068 14624 8072 14680
rect 8008 14620 8072 14624
rect 8088 14680 8152 14684
rect 8088 14624 8092 14680
rect 8092 14624 8148 14680
rect 8148 14624 8152 14680
rect 8088 14620 8152 14624
rect 12413 14680 12477 14684
rect 12413 14624 12417 14680
rect 12417 14624 12473 14680
rect 12473 14624 12477 14680
rect 12413 14620 12477 14624
rect 12493 14680 12557 14684
rect 12493 14624 12497 14680
rect 12497 14624 12553 14680
rect 12553 14624 12557 14680
rect 12493 14620 12557 14624
rect 12573 14680 12637 14684
rect 12573 14624 12577 14680
rect 12577 14624 12633 14680
rect 12633 14624 12637 14680
rect 12573 14620 12637 14624
rect 12653 14680 12717 14684
rect 12653 14624 12657 14680
rect 12657 14624 12713 14680
rect 12713 14624 12717 14680
rect 12653 14620 12717 14624
rect 5565 13866 5629 13870
rect 5565 13810 5569 13866
rect 5569 13810 5625 13866
rect 5625 13810 5629 13866
rect 5565 13806 5629 13810
rect 5645 13866 5709 13870
rect 5645 13810 5649 13866
rect 5649 13810 5705 13866
rect 5705 13810 5709 13866
rect 5645 13806 5709 13810
rect 5725 13866 5789 13870
rect 5725 13810 5729 13866
rect 5729 13810 5785 13866
rect 5785 13810 5789 13866
rect 5725 13806 5789 13810
rect 5805 13866 5869 13870
rect 5805 13810 5809 13866
rect 5809 13810 5865 13866
rect 5865 13810 5869 13866
rect 5805 13806 5869 13810
rect 10130 13866 10194 13870
rect 10130 13810 10134 13866
rect 10134 13810 10190 13866
rect 10190 13810 10194 13866
rect 10130 13806 10194 13810
rect 10210 13866 10274 13870
rect 10210 13810 10214 13866
rect 10214 13810 10270 13866
rect 10270 13810 10274 13866
rect 10210 13806 10274 13810
rect 10290 13866 10354 13870
rect 10290 13810 10294 13866
rect 10294 13810 10350 13866
rect 10350 13810 10354 13866
rect 10290 13806 10354 13810
rect 10370 13866 10434 13870
rect 10370 13810 10374 13866
rect 10374 13810 10430 13866
rect 10430 13810 10434 13866
rect 10370 13806 10434 13810
rect 3282 13052 3346 13056
rect 3282 12996 3286 13052
rect 3286 12996 3342 13052
rect 3342 12996 3346 13052
rect 3282 12992 3346 12996
rect 3362 13052 3426 13056
rect 3362 12996 3366 13052
rect 3366 12996 3422 13052
rect 3422 12996 3426 13052
rect 3362 12992 3426 12996
rect 3442 13052 3506 13056
rect 3442 12996 3446 13052
rect 3446 12996 3502 13052
rect 3502 12996 3506 13052
rect 3442 12992 3506 12996
rect 3522 13052 3586 13056
rect 3522 12996 3526 13052
rect 3526 12996 3582 13052
rect 3582 12996 3586 13052
rect 3522 12992 3586 12996
rect 7848 13052 7912 13056
rect 7848 12996 7852 13052
rect 7852 12996 7908 13052
rect 7908 12996 7912 13052
rect 7848 12992 7912 12996
rect 7928 13052 7992 13056
rect 7928 12996 7932 13052
rect 7932 12996 7988 13052
rect 7988 12996 7992 13052
rect 7928 12992 7992 12996
rect 8008 13052 8072 13056
rect 8008 12996 8012 13052
rect 8012 12996 8068 13052
rect 8068 12996 8072 13052
rect 8008 12992 8072 12996
rect 8088 13052 8152 13056
rect 8088 12996 8092 13052
rect 8092 12996 8148 13052
rect 8148 12996 8152 13052
rect 8088 12992 8152 12996
rect 12413 13052 12477 13056
rect 12413 12996 12417 13052
rect 12417 12996 12473 13052
rect 12473 12996 12477 13052
rect 12413 12992 12477 12996
rect 12493 13052 12557 13056
rect 12493 12996 12497 13052
rect 12497 12996 12553 13052
rect 12553 12996 12557 13052
rect 12493 12992 12557 12996
rect 12573 13052 12637 13056
rect 12573 12996 12577 13052
rect 12577 12996 12633 13052
rect 12633 12996 12637 13052
rect 12573 12992 12637 12996
rect 12653 13052 12717 13056
rect 12653 12996 12657 13052
rect 12657 12996 12713 13052
rect 12713 12996 12717 13052
rect 12653 12992 12717 12996
rect 5565 12238 5629 12242
rect 5565 12182 5569 12238
rect 5569 12182 5625 12238
rect 5625 12182 5629 12238
rect 5565 12178 5629 12182
rect 5645 12238 5709 12242
rect 5645 12182 5649 12238
rect 5649 12182 5705 12238
rect 5705 12182 5709 12238
rect 5645 12178 5709 12182
rect 5725 12238 5789 12242
rect 5725 12182 5729 12238
rect 5729 12182 5785 12238
rect 5785 12182 5789 12238
rect 5725 12178 5789 12182
rect 5805 12238 5869 12242
rect 5805 12182 5809 12238
rect 5809 12182 5865 12238
rect 5865 12182 5869 12238
rect 5805 12178 5869 12182
rect 10130 12238 10194 12242
rect 10130 12182 10134 12238
rect 10134 12182 10190 12238
rect 10190 12182 10194 12238
rect 10130 12178 10194 12182
rect 10210 12238 10274 12242
rect 10210 12182 10214 12238
rect 10214 12182 10270 12238
rect 10270 12182 10274 12238
rect 10210 12178 10274 12182
rect 10290 12238 10354 12242
rect 10290 12182 10294 12238
rect 10294 12182 10350 12238
rect 10350 12182 10354 12238
rect 10290 12178 10354 12182
rect 10370 12238 10434 12242
rect 10370 12182 10374 12238
rect 10374 12182 10430 12238
rect 10430 12182 10434 12238
rect 10370 12178 10434 12182
rect 3282 11424 3346 11428
rect 3282 11368 3286 11424
rect 3286 11368 3342 11424
rect 3342 11368 3346 11424
rect 3282 11364 3346 11368
rect 3362 11424 3426 11428
rect 3362 11368 3366 11424
rect 3366 11368 3422 11424
rect 3422 11368 3426 11424
rect 3362 11364 3426 11368
rect 3442 11424 3506 11428
rect 3442 11368 3446 11424
rect 3446 11368 3502 11424
rect 3502 11368 3506 11424
rect 3442 11364 3506 11368
rect 3522 11424 3586 11428
rect 3522 11368 3526 11424
rect 3526 11368 3582 11424
rect 3582 11368 3586 11424
rect 3522 11364 3586 11368
rect 7848 11424 7912 11428
rect 7848 11368 7852 11424
rect 7852 11368 7908 11424
rect 7908 11368 7912 11424
rect 7848 11364 7912 11368
rect 7928 11424 7992 11428
rect 7928 11368 7932 11424
rect 7932 11368 7988 11424
rect 7988 11368 7992 11424
rect 7928 11364 7992 11368
rect 8008 11424 8072 11428
rect 8008 11368 8012 11424
rect 8012 11368 8068 11424
rect 8068 11368 8072 11424
rect 8008 11364 8072 11368
rect 8088 11424 8152 11428
rect 8088 11368 8092 11424
rect 8092 11368 8148 11424
rect 8148 11368 8152 11424
rect 8088 11364 8152 11368
rect 12413 11424 12477 11428
rect 12413 11368 12417 11424
rect 12417 11368 12473 11424
rect 12473 11368 12477 11424
rect 12413 11364 12477 11368
rect 12493 11424 12557 11428
rect 12493 11368 12497 11424
rect 12497 11368 12553 11424
rect 12553 11368 12557 11424
rect 12493 11364 12557 11368
rect 12573 11424 12637 11428
rect 12573 11368 12577 11424
rect 12577 11368 12633 11424
rect 12633 11368 12637 11424
rect 12573 11364 12637 11368
rect 12653 11424 12717 11428
rect 12653 11368 12657 11424
rect 12657 11368 12713 11424
rect 12713 11368 12717 11424
rect 12653 11364 12717 11368
rect 5565 10610 5629 10614
rect 5565 10554 5569 10610
rect 5569 10554 5625 10610
rect 5625 10554 5629 10610
rect 5565 10550 5629 10554
rect 5645 10610 5709 10614
rect 5645 10554 5649 10610
rect 5649 10554 5705 10610
rect 5705 10554 5709 10610
rect 5645 10550 5709 10554
rect 5725 10610 5789 10614
rect 5725 10554 5729 10610
rect 5729 10554 5785 10610
rect 5785 10554 5789 10610
rect 5725 10550 5789 10554
rect 5805 10610 5869 10614
rect 5805 10554 5809 10610
rect 5809 10554 5865 10610
rect 5865 10554 5869 10610
rect 5805 10550 5869 10554
rect 10130 10610 10194 10614
rect 10130 10554 10134 10610
rect 10134 10554 10190 10610
rect 10190 10554 10194 10610
rect 10130 10550 10194 10554
rect 10210 10610 10274 10614
rect 10210 10554 10214 10610
rect 10214 10554 10270 10610
rect 10270 10554 10274 10610
rect 10210 10550 10274 10554
rect 10290 10610 10354 10614
rect 10290 10554 10294 10610
rect 10294 10554 10350 10610
rect 10350 10554 10354 10610
rect 10290 10550 10354 10554
rect 10370 10610 10434 10614
rect 10370 10554 10374 10610
rect 10374 10554 10430 10610
rect 10430 10554 10434 10610
rect 10370 10550 10434 10554
rect 3282 9796 3346 9800
rect 3282 9740 3286 9796
rect 3286 9740 3342 9796
rect 3342 9740 3346 9796
rect 3282 9736 3346 9740
rect 3362 9796 3426 9800
rect 3362 9740 3366 9796
rect 3366 9740 3422 9796
rect 3422 9740 3426 9796
rect 3362 9736 3426 9740
rect 3442 9796 3506 9800
rect 3442 9740 3446 9796
rect 3446 9740 3502 9796
rect 3502 9740 3506 9796
rect 3442 9736 3506 9740
rect 3522 9796 3586 9800
rect 3522 9740 3526 9796
rect 3526 9740 3582 9796
rect 3582 9740 3586 9796
rect 3522 9736 3586 9740
rect 7848 9796 7912 9800
rect 7848 9740 7852 9796
rect 7852 9740 7908 9796
rect 7908 9740 7912 9796
rect 7848 9736 7912 9740
rect 7928 9796 7992 9800
rect 7928 9740 7932 9796
rect 7932 9740 7988 9796
rect 7988 9740 7992 9796
rect 7928 9736 7992 9740
rect 8008 9796 8072 9800
rect 8008 9740 8012 9796
rect 8012 9740 8068 9796
rect 8068 9740 8072 9796
rect 8008 9736 8072 9740
rect 8088 9796 8152 9800
rect 8088 9740 8092 9796
rect 8092 9740 8148 9796
rect 8148 9740 8152 9796
rect 8088 9736 8152 9740
rect 12413 9796 12477 9800
rect 12413 9740 12417 9796
rect 12417 9740 12473 9796
rect 12473 9740 12477 9796
rect 12413 9736 12477 9740
rect 12493 9796 12557 9800
rect 12493 9740 12497 9796
rect 12497 9740 12553 9796
rect 12553 9740 12557 9796
rect 12493 9736 12557 9740
rect 12573 9796 12637 9800
rect 12573 9740 12577 9796
rect 12577 9740 12633 9796
rect 12633 9740 12637 9796
rect 12573 9736 12637 9740
rect 12653 9796 12717 9800
rect 12653 9740 12657 9796
rect 12657 9740 12713 9796
rect 12713 9740 12717 9796
rect 12653 9736 12717 9740
rect 5565 8982 5629 8986
rect 5565 8926 5569 8982
rect 5569 8926 5625 8982
rect 5625 8926 5629 8982
rect 5565 8922 5629 8926
rect 5645 8982 5709 8986
rect 5645 8926 5649 8982
rect 5649 8926 5705 8982
rect 5705 8926 5709 8982
rect 5645 8922 5709 8926
rect 5725 8982 5789 8986
rect 5725 8926 5729 8982
rect 5729 8926 5785 8982
rect 5785 8926 5789 8982
rect 5725 8922 5789 8926
rect 5805 8982 5869 8986
rect 5805 8926 5809 8982
rect 5809 8926 5865 8982
rect 5865 8926 5869 8982
rect 5805 8922 5869 8926
rect 10130 8982 10194 8986
rect 10130 8926 10134 8982
rect 10134 8926 10190 8982
rect 10190 8926 10194 8982
rect 10130 8922 10194 8926
rect 10210 8982 10274 8986
rect 10210 8926 10214 8982
rect 10214 8926 10270 8982
rect 10270 8926 10274 8982
rect 10210 8922 10274 8926
rect 10290 8982 10354 8986
rect 10290 8926 10294 8982
rect 10294 8926 10350 8982
rect 10350 8926 10354 8982
rect 10290 8922 10354 8926
rect 10370 8982 10434 8986
rect 10370 8926 10374 8982
rect 10374 8926 10430 8982
rect 10430 8926 10434 8982
rect 10370 8922 10434 8926
rect 3282 8168 3346 8172
rect 3282 8112 3286 8168
rect 3286 8112 3342 8168
rect 3342 8112 3346 8168
rect 3282 8108 3346 8112
rect 3362 8168 3426 8172
rect 3362 8112 3366 8168
rect 3366 8112 3422 8168
rect 3422 8112 3426 8168
rect 3362 8108 3426 8112
rect 3442 8168 3506 8172
rect 3442 8112 3446 8168
rect 3446 8112 3502 8168
rect 3502 8112 3506 8168
rect 3442 8108 3506 8112
rect 3522 8168 3586 8172
rect 3522 8112 3526 8168
rect 3526 8112 3582 8168
rect 3582 8112 3586 8168
rect 3522 8108 3586 8112
rect 7848 8168 7912 8172
rect 7848 8112 7852 8168
rect 7852 8112 7908 8168
rect 7908 8112 7912 8168
rect 7848 8108 7912 8112
rect 7928 8168 7992 8172
rect 7928 8112 7932 8168
rect 7932 8112 7988 8168
rect 7988 8112 7992 8168
rect 7928 8108 7992 8112
rect 8008 8168 8072 8172
rect 8008 8112 8012 8168
rect 8012 8112 8068 8168
rect 8068 8112 8072 8168
rect 8008 8108 8072 8112
rect 8088 8168 8152 8172
rect 8088 8112 8092 8168
rect 8092 8112 8148 8168
rect 8148 8112 8152 8168
rect 8088 8108 8152 8112
rect 12413 8168 12477 8172
rect 12413 8112 12417 8168
rect 12417 8112 12473 8168
rect 12473 8112 12477 8168
rect 12413 8108 12477 8112
rect 12493 8168 12557 8172
rect 12493 8112 12497 8168
rect 12497 8112 12553 8168
rect 12553 8112 12557 8168
rect 12493 8108 12557 8112
rect 12573 8168 12637 8172
rect 12573 8112 12577 8168
rect 12577 8112 12633 8168
rect 12633 8112 12637 8168
rect 12573 8108 12637 8112
rect 12653 8168 12717 8172
rect 12653 8112 12657 8168
rect 12657 8112 12713 8168
rect 12713 8112 12717 8168
rect 12653 8108 12717 8112
rect 5565 7354 5629 7358
rect 5565 7298 5569 7354
rect 5569 7298 5625 7354
rect 5625 7298 5629 7354
rect 5565 7294 5629 7298
rect 5645 7354 5709 7358
rect 5645 7298 5649 7354
rect 5649 7298 5705 7354
rect 5705 7298 5709 7354
rect 5645 7294 5709 7298
rect 5725 7354 5789 7358
rect 5725 7298 5729 7354
rect 5729 7298 5785 7354
rect 5785 7298 5789 7354
rect 5725 7294 5789 7298
rect 5805 7354 5869 7358
rect 5805 7298 5809 7354
rect 5809 7298 5865 7354
rect 5865 7298 5869 7354
rect 5805 7294 5869 7298
rect 10130 7354 10194 7358
rect 10130 7298 10134 7354
rect 10134 7298 10190 7354
rect 10190 7298 10194 7354
rect 10130 7294 10194 7298
rect 10210 7354 10274 7358
rect 10210 7298 10214 7354
rect 10214 7298 10270 7354
rect 10270 7298 10274 7354
rect 10210 7294 10274 7298
rect 10290 7354 10354 7358
rect 10290 7298 10294 7354
rect 10294 7298 10350 7354
rect 10350 7298 10354 7354
rect 10290 7294 10354 7298
rect 10370 7354 10434 7358
rect 10370 7298 10374 7354
rect 10374 7298 10430 7354
rect 10430 7298 10434 7354
rect 10370 7294 10434 7298
rect 3282 6540 3346 6544
rect 3282 6484 3286 6540
rect 3286 6484 3342 6540
rect 3342 6484 3346 6540
rect 3282 6480 3346 6484
rect 3362 6540 3426 6544
rect 3362 6484 3366 6540
rect 3366 6484 3422 6540
rect 3422 6484 3426 6540
rect 3362 6480 3426 6484
rect 3442 6540 3506 6544
rect 3442 6484 3446 6540
rect 3446 6484 3502 6540
rect 3502 6484 3506 6540
rect 3442 6480 3506 6484
rect 3522 6540 3586 6544
rect 3522 6484 3526 6540
rect 3526 6484 3582 6540
rect 3582 6484 3586 6540
rect 3522 6480 3586 6484
rect 7848 6540 7912 6544
rect 7848 6484 7852 6540
rect 7852 6484 7908 6540
rect 7908 6484 7912 6540
rect 7848 6480 7912 6484
rect 7928 6540 7992 6544
rect 7928 6484 7932 6540
rect 7932 6484 7988 6540
rect 7988 6484 7992 6540
rect 7928 6480 7992 6484
rect 8008 6540 8072 6544
rect 8008 6484 8012 6540
rect 8012 6484 8068 6540
rect 8068 6484 8072 6540
rect 8008 6480 8072 6484
rect 8088 6540 8152 6544
rect 8088 6484 8092 6540
rect 8092 6484 8148 6540
rect 8148 6484 8152 6540
rect 8088 6480 8152 6484
rect 12413 6540 12477 6544
rect 12413 6484 12417 6540
rect 12417 6484 12473 6540
rect 12473 6484 12477 6540
rect 12413 6480 12477 6484
rect 12493 6540 12557 6544
rect 12493 6484 12497 6540
rect 12497 6484 12553 6540
rect 12553 6484 12557 6540
rect 12493 6480 12557 6484
rect 12573 6540 12637 6544
rect 12573 6484 12577 6540
rect 12577 6484 12633 6540
rect 12633 6484 12637 6540
rect 12573 6480 12637 6484
rect 12653 6540 12717 6544
rect 12653 6484 12657 6540
rect 12657 6484 12713 6540
rect 12713 6484 12717 6540
rect 12653 6480 12717 6484
rect 5565 5726 5629 5730
rect 5565 5670 5569 5726
rect 5569 5670 5625 5726
rect 5625 5670 5629 5726
rect 5565 5666 5629 5670
rect 5645 5726 5709 5730
rect 5645 5670 5649 5726
rect 5649 5670 5705 5726
rect 5705 5670 5709 5726
rect 5645 5666 5709 5670
rect 5725 5726 5789 5730
rect 5725 5670 5729 5726
rect 5729 5670 5785 5726
rect 5785 5670 5789 5726
rect 5725 5666 5789 5670
rect 5805 5726 5869 5730
rect 5805 5670 5809 5726
rect 5809 5670 5865 5726
rect 5865 5670 5869 5726
rect 5805 5666 5869 5670
rect 10130 5726 10194 5730
rect 10130 5670 10134 5726
rect 10134 5670 10190 5726
rect 10190 5670 10194 5726
rect 10130 5666 10194 5670
rect 10210 5726 10274 5730
rect 10210 5670 10214 5726
rect 10214 5670 10270 5726
rect 10270 5670 10274 5726
rect 10210 5666 10274 5670
rect 10290 5726 10354 5730
rect 10290 5670 10294 5726
rect 10294 5670 10350 5726
rect 10350 5670 10354 5726
rect 10290 5666 10354 5670
rect 10370 5726 10434 5730
rect 10370 5670 10374 5726
rect 10374 5670 10430 5726
rect 10430 5670 10434 5726
rect 10370 5666 10434 5670
rect 3282 4912 3346 4916
rect 3282 4856 3286 4912
rect 3286 4856 3342 4912
rect 3342 4856 3346 4912
rect 3282 4852 3346 4856
rect 3362 4912 3426 4916
rect 3362 4856 3366 4912
rect 3366 4856 3422 4912
rect 3422 4856 3426 4912
rect 3362 4852 3426 4856
rect 3442 4912 3506 4916
rect 3442 4856 3446 4912
rect 3446 4856 3502 4912
rect 3502 4856 3506 4912
rect 3442 4852 3506 4856
rect 3522 4912 3586 4916
rect 3522 4856 3526 4912
rect 3526 4856 3582 4912
rect 3582 4856 3586 4912
rect 3522 4852 3586 4856
rect 7848 4912 7912 4916
rect 7848 4856 7852 4912
rect 7852 4856 7908 4912
rect 7908 4856 7912 4912
rect 7848 4852 7912 4856
rect 7928 4912 7992 4916
rect 7928 4856 7932 4912
rect 7932 4856 7988 4912
rect 7988 4856 7992 4912
rect 7928 4852 7992 4856
rect 8008 4912 8072 4916
rect 8008 4856 8012 4912
rect 8012 4856 8068 4912
rect 8068 4856 8072 4912
rect 8008 4852 8072 4856
rect 8088 4912 8152 4916
rect 8088 4856 8092 4912
rect 8092 4856 8148 4912
rect 8148 4856 8152 4912
rect 8088 4852 8152 4856
rect 12413 4912 12477 4916
rect 12413 4856 12417 4912
rect 12417 4856 12473 4912
rect 12473 4856 12477 4912
rect 12413 4852 12477 4856
rect 12493 4912 12557 4916
rect 12493 4856 12497 4912
rect 12497 4856 12553 4912
rect 12553 4856 12557 4912
rect 12493 4852 12557 4856
rect 12573 4912 12637 4916
rect 12573 4856 12577 4912
rect 12577 4856 12633 4912
rect 12633 4856 12637 4912
rect 12573 4852 12637 4856
rect 12653 4912 12717 4916
rect 12653 4856 12657 4912
rect 12657 4856 12713 4912
rect 12713 4856 12717 4912
rect 12653 4852 12717 4856
rect 5565 4098 5629 4102
rect 5565 4042 5569 4098
rect 5569 4042 5625 4098
rect 5625 4042 5629 4098
rect 5565 4038 5629 4042
rect 5645 4098 5709 4102
rect 5645 4042 5649 4098
rect 5649 4042 5705 4098
rect 5705 4042 5709 4098
rect 5645 4038 5709 4042
rect 5725 4098 5789 4102
rect 5725 4042 5729 4098
rect 5729 4042 5785 4098
rect 5785 4042 5789 4098
rect 5725 4038 5789 4042
rect 5805 4098 5869 4102
rect 5805 4042 5809 4098
rect 5809 4042 5865 4098
rect 5865 4042 5869 4098
rect 5805 4038 5869 4042
rect 10130 4098 10194 4102
rect 10130 4042 10134 4098
rect 10134 4042 10190 4098
rect 10190 4042 10194 4098
rect 10130 4038 10194 4042
rect 10210 4098 10274 4102
rect 10210 4042 10214 4098
rect 10214 4042 10270 4098
rect 10270 4042 10274 4098
rect 10210 4038 10274 4042
rect 10290 4098 10354 4102
rect 10290 4042 10294 4098
rect 10294 4042 10350 4098
rect 10350 4042 10354 4098
rect 10290 4038 10354 4042
rect 10370 4098 10434 4102
rect 10370 4042 10374 4098
rect 10374 4042 10430 4098
rect 10430 4042 10434 4098
rect 10370 4038 10434 4042
rect 3282 3284 3346 3288
rect 3282 3228 3286 3284
rect 3286 3228 3342 3284
rect 3342 3228 3346 3284
rect 3282 3224 3346 3228
rect 3362 3284 3426 3288
rect 3362 3228 3366 3284
rect 3366 3228 3422 3284
rect 3422 3228 3426 3284
rect 3362 3224 3426 3228
rect 3442 3284 3506 3288
rect 3442 3228 3446 3284
rect 3446 3228 3502 3284
rect 3502 3228 3506 3284
rect 3442 3224 3506 3228
rect 3522 3284 3586 3288
rect 3522 3228 3526 3284
rect 3526 3228 3582 3284
rect 3582 3228 3586 3284
rect 3522 3224 3586 3228
rect 7848 3284 7912 3288
rect 7848 3228 7852 3284
rect 7852 3228 7908 3284
rect 7908 3228 7912 3284
rect 7848 3224 7912 3228
rect 7928 3284 7992 3288
rect 7928 3228 7932 3284
rect 7932 3228 7988 3284
rect 7988 3228 7992 3284
rect 7928 3224 7992 3228
rect 8008 3284 8072 3288
rect 8008 3228 8012 3284
rect 8012 3228 8068 3284
rect 8068 3228 8072 3284
rect 8008 3224 8072 3228
rect 8088 3284 8152 3288
rect 8088 3228 8092 3284
rect 8092 3228 8148 3284
rect 8148 3228 8152 3284
rect 8088 3224 8152 3228
rect 12413 3284 12477 3288
rect 12413 3228 12417 3284
rect 12417 3228 12473 3284
rect 12473 3228 12477 3284
rect 12413 3224 12477 3228
rect 12493 3284 12557 3288
rect 12493 3228 12497 3284
rect 12497 3228 12553 3284
rect 12553 3228 12557 3284
rect 12493 3224 12557 3228
rect 12573 3284 12637 3288
rect 12573 3228 12577 3284
rect 12577 3228 12633 3284
rect 12633 3228 12637 3284
rect 12573 3224 12637 3228
rect 12653 3284 12717 3288
rect 12653 3228 12657 3284
rect 12657 3228 12713 3284
rect 12713 3228 12717 3284
rect 12653 3224 12717 3228
<< metal4 >>
rect 3274 16312 3595 16331
rect 3274 16248 3282 16312
rect 3346 16248 3362 16312
rect 3426 16248 3442 16312
rect 3506 16248 3522 16312
rect 3586 16248 3595 16312
rect 3274 14684 3595 16248
rect 3274 14620 3282 14684
rect 3346 14620 3362 14684
rect 3426 14620 3442 14684
rect 3506 14620 3522 14684
rect 3586 14620 3595 14684
rect 3274 13056 3595 14620
rect 3274 12992 3282 13056
rect 3346 12992 3362 13056
rect 3426 12992 3442 13056
rect 3506 12992 3522 13056
rect 3586 12992 3595 13056
rect 3274 11428 3595 12992
rect 3274 11364 3282 11428
rect 3346 11364 3362 11428
rect 3426 11364 3442 11428
rect 3506 11364 3522 11428
rect 3586 11364 3595 11428
rect 3274 9800 3595 11364
rect 3274 9736 3282 9800
rect 3346 9736 3362 9800
rect 3426 9736 3442 9800
rect 3506 9736 3522 9800
rect 3586 9736 3595 9800
rect 3274 8172 3595 9736
rect 3274 8108 3282 8172
rect 3346 8108 3362 8172
rect 3426 8108 3442 8172
rect 3506 8108 3522 8172
rect 3586 8108 3595 8172
rect 3274 6544 3595 8108
rect 3274 6480 3282 6544
rect 3346 6480 3362 6544
rect 3426 6480 3442 6544
rect 3506 6480 3522 6544
rect 3586 6480 3595 6544
rect 3274 4916 3595 6480
rect 3274 4852 3282 4916
rect 3346 4852 3362 4916
rect 3426 4852 3442 4916
rect 3506 4852 3522 4916
rect 3586 4852 3595 4916
rect 3274 3288 3595 4852
rect 3274 3224 3282 3288
rect 3346 3224 3362 3288
rect 3426 3224 3442 3288
rect 3506 3224 3522 3288
rect 3586 3224 3595 3288
rect 3274 3205 3595 3224
rect 5557 15498 5877 16331
rect 5557 15434 5565 15498
rect 5629 15434 5645 15498
rect 5709 15434 5725 15498
rect 5789 15434 5805 15498
rect 5869 15434 5877 15498
rect 5557 13870 5877 15434
rect 5557 13806 5565 13870
rect 5629 13806 5645 13870
rect 5709 13806 5725 13870
rect 5789 13806 5805 13870
rect 5869 13806 5877 13870
rect 5557 12242 5877 13806
rect 5557 12178 5565 12242
rect 5629 12178 5645 12242
rect 5709 12178 5725 12242
rect 5789 12178 5805 12242
rect 5869 12178 5877 12242
rect 5557 10614 5877 12178
rect 5557 10550 5565 10614
rect 5629 10550 5645 10614
rect 5709 10550 5725 10614
rect 5789 10550 5805 10614
rect 5869 10550 5877 10614
rect 5557 8986 5877 10550
rect 5557 8922 5565 8986
rect 5629 8922 5645 8986
rect 5709 8922 5725 8986
rect 5789 8922 5805 8986
rect 5869 8922 5877 8986
rect 5557 7358 5877 8922
rect 5557 7294 5565 7358
rect 5629 7294 5645 7358
rect 5709 7294 5725 7358
rect 5789 7294 5805 7358
rect 5869 7294 5877 7358
rect 5557 5730 5877 7294
rect 5557 5666 5565 5730
rect 5629 5666 5645 5730
rect 5709 5666 5725 5730
rect 5789 5666 5805 5730
rect 5869 5666 5877 5730
rect 5557 4102 5877 5666
rect 5557 4038 5565 4102
rect 5629 4038 5645 4102
rect 5709 4038 5725 4102
rect 5789 4038 5805 4102
rect 5869 4038 5877 4102
rect 5557 3205 5877 4038
rect 7840 16312 8160 16331
rect 7840 16248 7848 16312
rect 7912 16248 7928 16312
rect 7992 16248 8008 16312
rect 8072 16248 8088 16312
rect 8152 16248 8160 16312
rect 7840 14684 8160 16248
rect 7840 14620 7848 14684
rect 7912 14620 7928 14684
rect 7992 14620 8008 14684
rect 8072 14620 8088 14684
rect 8152 14620 8160 14684
rect 7840 13056 8160 14620
rect 7840 12992 7848 13056
rect 7912 12992 7928 13056
rect 7992 12992 8008 13056
rect 8072 12992 8088 13056
rect 8152 12992 8160 13056
rect 7840 11428 8160 12992
rect 7840 11364 7848 11428
rect 7912 11364 7928 11428
rect 7992 11364 8008 11428
rect 8072 11364 8088 11428
rect 8152 11364 8160 11428
rect 7840 9800 8160 11364
rect 7840 9736 7848 9800
rect 7912 9736 7928 9800
rect 7992 9736 8008 9800
rect 8072 9736 8088 9800
rect 8152 9736 8160 9800
rect 7840 8172 8160 9736
rect 7840 8108 7848 8172
rect 7912 8108 7928 8172
rect 7992 8108 8008 8172
rect 8072 8108 8088 8172
rect 8152 8108 8160 8172
rect 7840 6544 8160 8108
rect 7840 6480 7848 6544
rect 7912 6480 7928 6544
rect 7992 6480 8008 6544
rect 8072 6480 8088 6544
rect 8152 6480 8160 6544
rect 7840 4916 8160 6480
rect 7840 4852 7848 4916
rect 7912 4852 7928 4916
rect 7992 4852 8008 4916
rect 8072 4852 8088 4916
rect 8152 4852 8160 4916
rect 7840 3288 8160 4852
rect 7840 3224 7848 3288
rect 7912 3224 7928 3288
rect 7992 3224 8008 3288
rect 8072 3224 8088 3288
rect 8152 3224 8160 3288
rect 7840 3205 8160 3224
rect 10122 15498 10443 16331
rect 10122 15434 10130 15498
rect 10194 15434 10210 15498
rect 10274 15434 10290 15498
rect 10354 15434 10370 15498
rect 10434 15434 10443 15498
rect 10122 13870 10443 15434
rect 10122 13806 10130 13870
rect 10194 13806 10210 13870
rect 10274 13806 10290 13870
rect 10354 13806 10370 13870
rect 10434 13806 10443 13870
rect 10122 12242 10443 13806
rect 10122 12178 10130 12242
rect 10194 12178 10210 12242
rect 10274 12178 10290 12242
rect 10354 12178 10370 12242
rect 10434 12178 10443 12242
rect 10122 10614 10443 12178
rect 10122 10550 10130 10614
rect 10194 10550 10210 10614
rect 10274 10550 10290 10614
rect 10354 10550 10370 10614
rect 10434 10550 10443 10614
rect 10122 8986 10443 10550
rect 10122 8922 10130 8986
rect 10194 8922 10210 8986
rect 10274 8922 10290 8986
rect 10354 8922 10370 8986
rect 10434 8922 10443 8986
rect 10122 7358 10443 8922
rect 10122 7294 10130 7358
rect 10194 7294 10210 7358
rect 10274 7294 10290 7358
rect 10354 7294 10370 7358
rect 10434 7294 10443 7358
rect 10122 5730 10443 7294
rect 10122 5666 10130 5730
rect 10194 5666 10210 5730
rect 10274 5666 10290 5730
rect 10354 5666 10370 5730
rect 10434 5666 10443 5730
rect 10122 4102 10443 5666
rect 10122 4038 10130 4102
rect 10194 4038 10210 4102
rect 10274 4038 10290 4102
rect 10354 4038 10370 4102
rect 10434 4038 10443 4102
rect 10122 3205 10443 4038
rect 12405 16312 12725 16331
rect 12405 16248 12413 16312
rect 12477 16248 12493 16312
rect 12557 16248 12573 16312
rect 12637 16248 12653 16312
rect 12717 16248 12725 16312
rect 12405 14684 12725 16248
rect 12405 14620 12413 14684
rect 12477 14620 12493 14684
rect 12557 14620 12573 14684
rect 12637 14620 12653 14684
rect 12717 14620 12725 14684
rect 12405 13056 12725 14620
rect 12405 12992 12413 13056
rect 12477 12992 12493 13056
rect 12557 12992 12573 13056
rect 12637 12992 12653 13056
rect 12717 12992 12725 13056
rect 12405 11428 12725 12992
rect 12405 11364 12413 11428
rect 12477 11364 12493 11428
rect 12557 11364 12573 11428
rect 12637 11364 12653 11428
rect 12717 11364 12725 11428
rect 12405 9800 12725 11364
rect 12405 9736 12413 9800
rect 12477 9736 12493 9800
rect 12557 9736 12573 9800
rect 12637 9736 12653 9800
rect 12717 9736 12725 9800
rect 12405 8172 12725 9736
rect 12405 8108 12413 8172
rect 12477 8108 12493 8172
rect 12557 8108 12573 8172
rect 12637 8108 12653 8172
rect 12717 8108 12725 8172
rect 12405 6544 12725 8108
rect 12405 6480 12413 6544
rect 12477 6480 12493 6544
rect 12557 6480 12573 6544
rect 12637 6480 12653 6544
rect 12717 6480 12725 6544
rect 12405 4916 12725 6480
rect 12405 4852 12413 4916
rect 12477 4852 12493 4916
rect 12557 4852 12573 4916
rect 12637 4852 12653 4916
rect 12717 4852 12725 4916
rect 12405 3288 12725 4852
rect 12405 3224 12413 3288
rect 12477 3224 12493 3288
rect 12557 3224 12573 3288
rect 12637 3224 12653 3288
rect 12717 3224 12725 3288
rect 12405 3205 12725 3224
use sky130_fd_sc_hvl__decap_8  FILLER_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 1152 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_8
timestamp 1624635493
transform 1 0 1920 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_0
timestamp 1624635493
transform 1 0 1152 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_8
timestamp 1624635493
transform 1 0 1920 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_16
timestamp 1624635493
transform 1 0 2688 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_16
timestamp 1624635493
transform 1 0 2688 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_24
timestamp 1624635493
transform 1 0 3456 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_24
timestamp 1624635493
transform 1 0 3456 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_32
timestamp 1624635493
transform 1 0 4224 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_32
timestamp 1624635493
transform 1 0 4224 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_40
timestamp 1624635493
transform 1 0 4992 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_40
timestamp 1624635493
transform 1 0 4992 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_48
timestamp 1624635493
transform 1 0 5760 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_56
timestamp 1624635493
transform 1 0 6528 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_48
timestamp 1624635493
transform 1 0 5760 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_56
timestamp 1624635493
transform 1 0 6528 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_64
timestamp 1624635493
transform 1 0 7296 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_64
timestamp 1624635493
transform 1 0 7296 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_72
timestamp 1624635493
transform 1 0 8064 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_72
timestamp 1624635493
transform 1 0 8064 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_80
timestamp 1624635493
transform 1 0 8832 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_80
timestamp 1624635493
transform 1 0 8832 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_88
timestamp 1624635493
transform 1 0 9600 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_88
timestamp 1624635493
transform 1 0 9600 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_96
timestamp 1624635493
transform 1 0 10368 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_96
timestamp 1624635493
transform 1 0 10368 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__nand3_1  x1.x2 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform -1 0 12480 0 1 4070
box -66 -43 738 897
use sky130_fd_sc_hvl__diode_2  ANTENNA_x1.x2_A $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 11232 0 1 4070
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_104
timestamp 1624635493
transform 1 0 11136 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_112 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 11904 0 -1 4070
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_104 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 11136 0 1 4070
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_107
timestamp 1624635493
transform 1 0 11424 0 1 4070
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  ANTENNA_x1.x2_B
timestamp 1624635493
transform 1 0 12864 0 1 4070
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  ANTENNA_x1.x1_B
timestamp 1624635493
transform 1 0 12480 0 -1 4070
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_116 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 12288 0 -1 4070
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_120
timestamp 1624635493
transform 1 0 12672 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_118
timestamp 1624635493
transform 1 0 12480 0 1 4070
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_128
timestamp 1624635493
transform 1 0 13440 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_124
timestamp 1624635493
transform 1 0 13056 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_136
timestamp 1624635493
transform 1 0 14208 0 -1 4070
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_140
timestamp 1624635493
transform 1 0 14592 0 -1 4070
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_132
timestamp 1624635493
transform 1 0 13824 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__fill_2  FILLER_1_140
timestamp 1624635493
transform 1 0 14592 0 1 4070
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_0
timestamp 1624635493
transform 1 0 1152 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_8
timestamp 1624635493
transform 1 0 1920 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_16
timestamp 1624635493
transform 1 0 2688 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_24
timestamp 1624635493
transform 1 0 3456 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_32
timestamp 1624635493
transform 1 0 4224 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_40
timestamp 1624635493
transform 1 0 4992 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_48
timestamp 1624635493
transform 1 0 5760 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_56
timestamp 1624635493
transform 1 0 6528 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_64
timestamp 1624635493
transform 1 0 7296 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_72
timestamp 1624635493
transform 1 0 8064 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_80
timestamp 1624635493
transform 1 0 8832 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_88
timestamp 1624635493
transform 1 0 9600 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__diode_2  ANTENNA_x1.x1_A
timestamp 1624635493
transform 1 0 10560 0 -1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  FILLER_2_96
timestamp 1624635493
transform 1 0 10368 0 -1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_100
timestamp 1624635493
transform 1 0 10752 0 -1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__inv_1  x0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 11136 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__nand3_1  x1.x1
timestamp 1624635493
transform 1 0 11808 0 -1 5698
box -66 -43 738 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_107
timestamp 1624635493
transform 1 0 11424 0 -1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__nor3_1  x2.x1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 12864 0 -1 5698
box -66 -43 738 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_118
timestamp 1624635493
transform 1 0 12480 0 -1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_129
timestamp 1624635493
transform 1 0 13536 0 -1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  ANTENNA_x2.x1_B
timestamp 1624635493
transform 1 0 13920 0 -1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_135
timestamp 1624635493
transform 1 0 14112 0 -1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_2_139
timestamp 1624635493
transform 1 0 14496 0 -1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_141
timestamp 1624635493
transform 1 0 14688 0 -1 5698
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_0
timestamp 1624635493
transform 1 0 1152 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_8
timestamp 1624635493
transform 1 0 1920 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_16
timestamp 1624635493
transform 1 0 2688 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_24
timestamp 1624635493
transform 1 0 3456 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_32
timestamp 1624635493
transform 1 0 4224 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_40
timestamp 1624635493
transform 1 0 4992 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_48
timestamp 1624635493
transform 1 0 5760 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_56
timestamp 1624635493
transform 1 0 6528 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_64
timestamp 1624635493
transform 1 0 7296 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_72
timestamp 1624635493
transform 1 0 8064 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_80
timestamp 1624635493
transform 1 0 8832 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_88
timestamp 1624635493
transform 1 0 9600 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__diode_2  ANTENNA_x0_A
timestamp 1624635493
transform -1 0 11136 0 1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_4  FILLER_3_96
timestamp 1624635493
transform 1 0 10368 0 1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_3_100
timestamp 1624635493
transform 1 0 10752 0 1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__inv_4  x1.x3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624635493
transform 1 0 11712 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_3_104
timestamp 1624635493
transform 1 0 11136 0 1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_3_108
timestamp 1624635493
transform 1 0 11520 0 1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__nor3_1  x2.x2
timestamp 1624635493
transform 1 0 12864 0 1 5698
box -66 -43 738 897
use sky130_fd_sc_hvl__decap_4  FILLER_3_118
timestamp 1624635493
transform 1 0 12480 0 1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  FILLER_3_129
timestamp 1624635493
transform 1 0 13536 0 1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  ANTENNA_x2.x2_B
timestamp 1624635493
transform 1 0 13920 0 1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_4  FILLER_3_135
timestamp 1624635493
transform 1 0 14112 0 1 5698
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_3_139
timestamp 1624635493
transform 1 0 14496 0 1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_3_141
timestamp 1624635493
transform 1 0 14688 0 1 5698
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_0
timestamp 1624635493
transform 1 0 1152 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_8
timestamp 1624635493
transform 1 0 1920 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_16
timestamp 1624635493
transform 1 0 2688 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_24
timestamp 1624635493
transform 1 0 3456 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_32
timestamp 1624635493
transform 1 0 4224 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_40
timestamp 1624635493
transform 1 0 4992 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_48
timestamp 1624635493
transform 1 0 5760 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_56
timestamp 1624635493
transform 1 0 6528 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_64
timestamp 1624635493
transform 1 0 7296 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_72
timestamp 1624635493
transform 1 0 8064 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_80
timestamp 1624635493
transform 1 0 8832 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_88
timestamp 1624635493
transform 1 0 9600 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_96
timestamp 1624635493
transform 1 0 10368 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_4  x1.x4
timestamp 1624635493
transform -1 0 12480 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_4_104
timestamp 1624635493
transform 1 0 11136 0 -1 7326
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_4_108
timestamp 1624635493
transform 1 0 11520 0 -1 7326
box -66 -43 258 897
use sky130_fd_sc_hvl__nor3_1  x5
timestamp 1624635493
transform 1 0 12864 0 -1 7326
box -66 -43 738 897
use sky130_fd_sc_hvl__decap_4  FILLER_4_118
timestamp 1624635493
transform 1 0 12480 0 -1 7326
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_4_129
timestamp 1624635493
transform 1 0 13536 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_4_137
timestamp 1624635493
transform 1 0 14304 0 -1 7326
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  FILLER_4_141
timestamp 1624635493
transform 1 0 14688 0 -1 7326
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_0
timestamp 1624635493
transform 1 0 1152 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_8
timestamp 1624635493
transform 1 0 1920 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_16
timestamp 1624635493
transform 1 0 2688 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_24
timestamp 1624635493
transform 1 0 3456 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_32
timestamp 1624635493
transform 1 0 4224 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_40
timestamp 1624635493
transform 1 0 4992 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_48
timestamp 1624635493
transform 1 0 5760 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_56
timestamp 1624635493
transform 1 0 6528 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_64
timestamp 1624635493
transform 1 0 7296 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_72
timestamp 1624635493
transform 1 0 8064 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_80
timestamp 1624635493
transform 1 0 8832 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_88
timestamp 1624635493
transform 1 0 9600 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_96
timestamp 1624635493
transform 1 0 10368 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_104
timestamp 1624635493
transform 1 0 11136 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__fill_1  FILLER_5_112
timestamp 1624635493
transform 1 0 11904 0 1 7326
box -66 -43 162 897
use sky130_fd_sc_hvl__nor3_1  x6
timestamp 1624635493
transform 1 0 12000 0 1 7326
box -66 -43 738 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_120
timestamp 1624635493
transform 1 0 12672 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_5_128
timestamp 1624635493
transform 1 0 13440 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_5_136
timestamp 1624635493
transform 1 0 14208 0 1 7326
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_5_140
timestamp 1624635493
transform 1 0 14592 0 1 7326
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_0
timestamp 1624635493
transform 1 0 1152 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_8
timestamp 1624635493
transform 1 0 1920 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_16
timestamp 1624635493
transform 1 0 2688 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_24
timestamp 1624635493
transform 1 0 3456 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_32
timestamp 1624635493
transform 1 0 4224 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_40
timestamp 1624635493
transform 1 0 4992 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_48
timestamp 1624635493
transform 1 0 5760 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_56
timestamp 1624635493
transform 1 0 6528 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_64
timestamp 1624635493
transform 1 0 7296 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_72
timestamp 1624635493
transform 1 0 8064 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_80
timestamp 1624635493
transform 1 0 8832 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_88
timestamp 1624635493
transform 1 0 9600 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_96
timestamp 1624635493
transform 1 0 10368 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_104
timestamp 1624635493
transform 1 0 11136 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_112
timestamp 1624635493
transform 1 0 11904 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_120
timestamp 1624635493
transform 1 0 12672 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_6_128
timestamp 1624635493
transform 1 0 13440 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_6_136
timestamp 1624635493
transform 1 0 14208 0 -1 8954
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_6_140
timestamp 1624635493
transform 1 0 14592 0 -1 8954
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_0
timestamp 1624635493
transform 1 0 1152 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_8
timestamp 1624635493
transform 1 0 1920 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_0
timestamp 1624635493
transform 1 0 1152 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_8
timestamp 1624635493
transform 1 0 1920 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_16
timestamp 1624635493
transform 1 0 2688 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_16
timestamp 1624635493
transform 1 0 2688 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_24
timestamp 1624635493
transform 1 0 3456 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_24
timestamp 1624635493
transform 1 0 3456 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_32
timestamp 1624635493
transform 1 0 4224 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_32
timestamp 1624635493
transform 1 0 4224 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_40
timestamp 1624635493
transform 1 0 4992 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_40
timestamp 1624635493
transform 1 0 4992 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_48
timestamp 1624635493
transform 1 0 5760 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_56
timestamp 1624635493
transform 1 0 6528 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_48
timestamp 1624635493
transform 1 0 5760 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_56
timestamp 1624635493
transform 1 0 6528 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_64
timestamp 1624635493
transform 1 0 7296 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_64
timestamp 1624635493
transform 1 0 7296 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_72
timestamp 1624635493
transform 1 0 8064 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_72
timestamp 1624635493
transform 1 0 8064 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_80
timestamp 1624635493
transform 1 0 8832 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_80
timestamp 1624635493
transform 1 0 8832 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_88
timestamp 1624635493
transform 1 0 9600 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_88
timestamp 1624635493
transform 1 0 9600 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_96
timestamp 1624635493
transform 1 0 10368 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_96
timestamp 1624635493
transform 1 0 10368 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_104
timestamp 1624635493
transform 1 0 11136 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_112
timestamp 1624635493
transform 1 0 11904 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_104
timestamp 1624635493
transform 1 0 11136 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_112
timestamp 1624635493
transform 1 0 11904 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_120
timestamp 1624635493
transform 1 0 12672 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_120
timestamp 1624635493
transform 1 0 12672 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_7_128
timestamp 1624635493
transform 1 0 13440 0 1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_8_128
timestamp 1624635493
transform 1 0 13440 0 -1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_7_136
timestamp 1624635493
transform 1 0 14208 0 1 8954
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_7_140
timestamp 1624635493
transform 1 0 14592 0 1 8954
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_4  FILLER_8_136
timestamp 1624635493
transform 1 0 14208 0 -1 10582
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_8_140
timestamp 1624635493
transform 1 0 14592 0 -1 10582
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_0
timestamp 1624635493
transform 1 0 1152 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_8
timestamp 1624635493
transform 1 0 1920 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_16
timestamp 1624635493
transform 1 0 2688 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_24
timestamp 1624635493
transform 1 0 3456 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_32
timestamp 1624635493
transform 1 0 4224 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_40
timestamp 1624635493
transform 1 0 4992 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_48
timestamp 1624635493
transform 1 0 5760 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_56
timestamp 1624635493
transform 1 0 6528 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_64
timestamp 1624635493
transform 1 0 7296 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_72
timestamp 1624635493
transform 1 0 8064 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_80
timestamp 1624635493
transform 1 0 8832 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_88
timestamp 1624635493
transform 1 0 9600 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_96
timestamp 1624635493
transform 1 0 10368 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_104
timestamp 1624635493
transform 1 0 11136 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_112
timestamp 1624635493
transform 1 0 11904 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_120
timestamp 1624635493
transform 1 0 12672 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_9_128
timestamp 1624635493
transform 1 0 13440 0 1 10582
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_9_136
timestamp 1624635493
transform 1 0 14208 0 1 10582
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_9_140
timestamp 1624635493
transform 1 0 14592 0 1 10582
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_0
timestamp 1624635493
transform 1 0 1152 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_8
timestamp 1624635493
transform 1 0 1920 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_16
timestamp 1624635493
transform 1 0 2688 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_24
timestamp 1624635493
transform 1 0 3456 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_32
timestamp 1624635493
transform 1 0 4224 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_40
timestamp 1624635493
transform 1 0 4992 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_48
timestamp 1624635493
transform 1 0 5760 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_56
timestamp 1624635493
transform 1 0 6528 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_64
timestamp 1624635493
transform 1 0 7296 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_72
timestamp 1624635493
transform 1 0 8064 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_80
timestamp 1624635493
transform 1 0 8832 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_88
timestamp 1624635493
transform 1 0 9600 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_96
timestamp 1624635493
transform 1 0 10368 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_104
timestamp 1624635493
transform 1 0 11136 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_112
timestamp 1624635493
transform 1 0 11904 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_120
timestamp 1624635493
transform 1 0 12672 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_10_128
timestamp 1624635493
transform 1 0 13440 0 -1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_10_136
timestamp 1624635493
transform 1 0 14208 0 -1 12210
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_10_140
timestamp 1624635493
transform 1 0 14592 0 -1 12210
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_0
timestamp 1624635493
transform 1 0 1152 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_8
timestamp 1624635493
transform 1 0 1920 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_16
timestamp 1624635493
transform 1 0 2688 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_24
timestamp 1624635493
transform 1 0 3456 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_32
timestamp 1624635493
transform 1 0 4224 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_40
timestamp 1624635493
transform 1 0 4992 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_48
timestamp 1624635493
transform 1 0 5760 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_56
timestamp 1624635493
transform 1 0 6528 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_64
timestamp 1624635493
transform 1 0 7296 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_72
timestamp 1624635493
transform 1 0 8064 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_80
timestamp 1624635493
transform 1 0 8832 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_88
timestamp 1624635493
transform 1 0 9600 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_96
timestamp 1624635493
transform 1 0 10368 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_104
timestamp 1624635493
transform 1 0 11136 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_112
timestamp 1624635493
transform 1 0 11904 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_120
timestamp 1624635493
transform 1 0 12672 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_11_128
timestamp 1624635493
transform 1 0 13440 0 1 12210
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_11_136
timestamp 1624635493
transform 1 0 14208 0 1 12210
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_11_140
timestamp 1624635493
transform 1 0 14592 0 1 12210
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_0
timestamp 1624635493
transform 1 0 1152 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_8
timestamp 1624635493
transform 1 0 1920 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_16
timestamp 1624635493
transform 1 0 2688 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_24
timestamp 1624635493
transform 1 0 3456 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_32
timestamp 1624635493
transform 1 0 4224 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_40
timestamp 1624635493
transform 1 0 4992 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_48
timestamp 1624635493
transform 1 0 5760 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_56
timestamp 1624635493
transform 1 0 6528 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_64
timestamp 1624635493
transform 1 0 7296 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_72
timestamp 1624635493
transform 1 0 8064 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_80
timestamp 1624635493
transform 1 0 8832 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_88
timestamp 1624635493
transform 1 0 9600 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_96
timestamp 1624635493
transform 1 0 10368 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_104
timestamp 1624635493
transform 1 0 11136 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_112
timestamp 1624635493
transform 1 0 11904 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_120
timestamp 1624635493
transform 1 0 12672 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_12_128
timestamp 1624635493
transform 1 0 13440 0 -1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_12_136
timestamp 1624635493
transform 1 0 14208 0 -1 13838
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_12_140
timestamp 1624635493
transform 1 0 14592 0 -1 13838
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_0
timestamp 1624635493
transform 1 0 1152 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_8
timestamp 1624635493
transform 1 0 1920 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_16
timestamp 1624635493
transform 1 0 2688 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_24
timestamp 1624635493
transform 1 0 3456 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_32
timestamp 1624635493
transform 1 0 4224 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_40
timestamp 1624635493
transform 1 0 4992 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_48
timestamp 1624635493
transform 1 0 5760 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_56
timestamp 1624635493
transform 1 0 6528 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_64
timestamp 1624635493
transform 1 0 7296 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_72
timestamp 1624635493
transform 1 0 8064 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_80
timestamp 1624635493
transform 1 0 8832 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_88
timestamp 1624635493
transform 1 0 9600 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_96
timestamp 1624635493
transform 1 0 10368 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_104
timestamp 1624635493
transform 1 0 11136 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_112
timestamp 1624635493
transform 1 0 11904 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_120
timestamp 1624635493
transform 1 0 12672 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_13_128
timestamp 1624635493
transform 1 0 13440 0 1 13838
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_13_136
timestamp 1624635493
transform 1 0 14208 0 1 13838
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_13_140
timestamp 1624635493
transform 1 0 14592 0 1 13838
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_0
timestamp 1624635493
transform 1 0 1152 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_8
timestamp 1624635493
transform 1 0 1920 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_16
timestamp 1624635493
transform 1 0 2688 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_24
timestamp 1624635493
transform 1 0 3456 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_32
timestamp 1624635493
transform 1 0 4224 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_40
timestamp 1624635493
transform 1 0 4992 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_48
timestamp 1624635493
transform 1 0 5760 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_56
timestamp 1624635493
transform 1 0 6528 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_64
timestamp 1624635493
transform 1 0 7296 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_72
timestamp 1624635493
transform 1 0 8064 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_80
timestamp 1624635493
transform 1 0 8832 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_88
timestamp 1624635493
transform 1 0 9600 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_96
timestamp 1624635493
transform 1 0 10368 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_104
timestamp 1624635493
transform 1 0 11136 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_112
timestamp 1624635493
transform 1 0 11904 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_120
timestamp 1624635493
transform 1 0 12672 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_14_128
timestamp 1624635493
transform 1 0 13440 0 -1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_14_136
timestamp 1624635493
transform 1 0 14208 0 -1 15466
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_14_140
timestamp 1624635493
transform 1 0 14592 0 -1 15466
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_0
timestamp 1624635493
transform 1 0 1152 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_8
timestamp 1624635493
transform 1 0 1920 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_16
timestamp 1624635493
transform 1 0 2688 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_24
timestamp 1624635493
transform 1 0 3456 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_32
timestamp 1624635493
transform 1 0 4224 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_40
timestamp 1624635493
transform 1 0 4992 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_48
timestamp 1624635493
transform 1 0 5760 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_56
timestamp 1624635493
transform 1 0 6528 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_64
timestamp 1624635493
transform 1 0 7296 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_72
timestamp 1624635493
transform 1 0 8064 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_80
timestamp 1624635493
transform 1 0 8832 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_88
timestamp 1624635493
transform 1 0 9600 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_96
timestamp 1624635493
transform 1 0 10368 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_104
timestamp 1624635493
transform 1 0 11136 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_112
timestamp 1624635493
transform 1 0 11904 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_120
timestamp 1624635493
transform 1 0 12672 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_15_128
timestamp 1624635493
transform 1 0 13440 0 1 15466
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_15_136
timestamp 1624635493
transform 1 0 14208 0 1 15466
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_15_140
timestamp 1624635493
transform 1 0 14592 0 1 15466
box -66 -43 258 897
<< labels >>
rlabel metal3 s 15200 9930 16000 10050 6 INN
port 0 nsew signal input
rlabel metal3 s 15200 3270 16000 3390 6 INP
port 1 nsew signal input
rlabel metal3 s 15200 16590 16000 16710 6 Q
port 2 nsew signal tristate
rlabel metal2 s 7988 0 8044 800 6 clk
port 3 nsew signal input
rlabel metal4 s 12405 3205 12725 16331 6 vccd2
port 4 nsew power bidirectional
rlabel metal4 s 7840 3205 8160 16331 6 vccd2
port 5 nsew power bidirectional
rlabel metal4 s 3275 3205 3595 16331 6 vccd2
port 6 nsew power bidirectional
rlabel metal4 s 10123 3205 10443 16331 6 vssd2
port 7 nsew ground bidirectional
rlabel metal4 s 5557 3205 5877 16331 6 vssd2
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 20000
<< end >>
