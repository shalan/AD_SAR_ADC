magic
tech sky130A
magscale 1 2
timestamp 1626105910
<< checkpaint >>
rect -1260 -1260 51260 48852
<< locali >>
rect 19073 14535 19107 15045
rect 27721 13991 27755 16541
rect 37473 12767 37507 13413
<< viali >>
rect 1869 47209 1903 47243
rect 1961 47073 1995 47107
rect 2605 47073 2639 47107
rect 22753 45441 22787 45475
rect 24869 45441 24903 45475
rect 23029 45373 23063 45407
rect 24409 45305 24443 45339
rect 22201 45237 22235 45271
rect 1961 42721 1995 42755
rect 39635 42721 39669 42755
rect 43617 42721 43651 42755
rect 39037 42653 39071 42687
rect 40693 42653 40727 42687
rect 43361 42653 43395 42687
rect 1869 42517 1903 42551
rect 2605 42517 2639 42551
rect 42809 42517 42843 42551
rect 44741 42517 44775 42551
rect 43177 41973 43211 42007
rect 7573 41701 7607 41735
rect 7021 41633 7055 41667
rect 13001 41633 13035 41667
rect 13369 41633 13403 41667
rect 47961 41633 47995 41667
rect 48145 41633 48179 41667
rect 13645 41565 13679 41599
rect 14381 41497 14415 41531
rect 6745 41429 6779 41463
rect 47317 41429 47351 41463
rect 13921 40885 13955 40919
rect 16681 39593 16715 39627
rect 15485 39525 15519 39559
rect 16037 39457 16071 39491
rect 22661 39457 22695 39491
rect 22937 39457 22971 39491
rect 23121 39457 23155 39491
rect 21925 39389 21959 39423
rect 22845 39389 22879 39423
rect 22753 39321 22787 39355
rect 22477 39253 22511 39287
rect 23673 39253 23707 39287
rect 24225 39253 24259 39287
rect 24685 38845 24719 38879
rect 25145 38845 25179 38879
rect 33517 38845 33551 38879
rect 33241 38777 33275 38811
rect 23581 38709 23615 38743
rect 24593 38709 24627 38743
rect 29101 38709 29135 38743
rect 32873 38505 32907 38539
rect 10057 38437 10091 38471
rect 5181 38369 5215 38403
rect 6101 38369 6135 38403
rect 9965 38369 9999 38403
rect 28365 38369 28399 38403
rect 28825 38369 28859 38403
rect 5457 38301 5491 38335
rect 10609 38301 10643 38335
rect 27997 38301 28031 38335
rect 28227 38233 28261 38267
rect 27721 38165 27755 38199
rect 28089 38165 28123 38199
rect 29377 38165 29411 38199
rect 28917 37621 28951 37655
rect 1869 37417 1903 37451
rect 1961 37281 1995 37315
rect 2605 37281 2639 37315
rect 17601 36873 17635 36907
rect 15025 36805 15059 36839
rect 16405 36737 16439 36771
rect 16160 36601 16194 36635
rect 13369 36533 13403 36567
rect 17049 36533 17083 36567
rect 11713 36329 11747 36363
rect 12449 36261 12483 36295
rect 12265 36193 12299 36227
rect 12541 36193 12575 36227
rect 12685 36193 12719 36227
rect 13461 36125 13495 36159
rect 12817 36057 12851 36091
rect 47225 35581 47259 35615
rect 47685 35581 47719 35615
rect 47777 35513 47811 35547
rect 13277 35445 13311 35479
rect 10425 34017 10459 34051
rect 10885 34017 10919 34051
rect 10241 33949 10275 33983
rect 38209 33813 38243 33847
rect 39129 33541 39163 33575
rect 38833 33405 38867 33439
rect 38577 33337 38611 33371
rect 38743 33337 38777 33371
rect 38945 33337 38979 33371
rect 38117 33269 38151 33303
rect 39589 33269 39623 33303
rect 40141 33269 40175 33303
rect 47041 33269 47075 33303
rect 37933 33065 37967 33099
rect 47041 32997 47075 33031
rect 47961 32997 47995 33031
rect 30481 32929 30515 32963
rect 38491 32929 38525 32963
rect 38761 32929 38795 32963
rect 47731 32929 47765 32963
rect 47869 32929 47903 32963
rect 48145 32929 48179 32963
rect 38577 32861 38611 32895
rect 38679 32861 38713 32895
rect 39497 32861 39531 32895
rect 38945 32793 38979 32827
rect 30665 32725 30699 32759
rect 40049 32725 40083 32759
rect 46581 32725 46615 32759
rect 47593 32725 47627 32759
rect 47225 32521 47259 32555
rect 1777 32385 1811 32419
rect 40693 32385 40727 32419
rect 1961 32249 1995 32283
rect 2605 32249 2639 32283
rect 40426 32249 40460 32283
rect 38025 32181 38059 32215
rect 38669 32181 38703 32215
rect 39313 32181 39347 32215
rect 21557 31977 21591 32011
rect 20913 31909 20947 31943
rect 20821 31841 20855 31875
rect 38945 31841 38979 31875
rect 39221 31841 39255 31875
rect 39865 31841 39899 31875
rect 3157 31773 3191 31807
rect 38301 31773 38335 31807
rect 39037 31773 39071 31807
rect 39129 31773 39163 31807
rect 39405 31773 39439 31807
rect 1777 31433 1811 31467
rect 39681 31433 39715 31467
rect 39129 31365 39163 31399
rect 2145 31297 2179 31331
rect 3525 31297 3559 31331
rect 1961 31229 1995 31263
rect 2053 31229 2087 31263
rect 2237 31229 2271 31263
rect 2421 31229 2455 31263
rect 2973 31161 3007 31195
rect 38577 31161 38611 31195
rect 4077 31093 4111 31127
rect 15669 30821 15703 30855
rect 15945 30753 15979 30787
rect 16405 30753 16439 30787
rect 34345 30753 34379 30787
rect 32505 30685 32539 30719
rect 34621 30685 34655 30719
rect 2973 30549 3007 30583
rect 33241 30549 33275 30583
rect 35081 30277 35115 30311
rect 35357 30277 35391 30311
rect 36185 30277 36219 30311
rect 33517 30209 33551 30243
rect 45385 30209 45419 30243
rect 35241 30141 35275 30175
rect 35449 30141 35483 30175
rect 35586 30141 35620 30175
rect 35725 30141 35759 30175
rect 45017 30141 45051 30175
rect 45477 30141 45511 30175
rect 33977 30073 34011 30107
rect 34529 30005 34563 30039
rect 44465 30005 44499 30039
rect 44005 29801 44039 29835
rect 25973 29665 26007 29699
rect 25605 29597 25639 29631
rect 25789 29597 25823 29631
rect 25881 29597 25915 29631
rect 26065 29597 26099 29631
rect 44649 29597 44683 29631
rect 25145 29529 25179 29563
rect 26709 29529 26743 29563
rect 27261 29461 27295 29495
rect 34713 29461 34747 29495
rect 44097 29257 44131 29291
rect 44925 29189 44959 29223
rect 44833 29121 44867 29155
rect 44741 29053 44775 29087
rect 45017 29053 45051 29087
rect 45201 29053 45235 29087
rect 25237 28985 25271 29019
rect 44557 28917 44591 28951
rect 22201 28713 22235 28747
rect 31033 28713 31067 28747
rect 36277 28713 36311 28747
rect 44189 28713 44223 28747
rect 38117 28509 38151 28543
rect 38393 28509 38427 28543
rect 37013 28373 37047 28407
rect 38853 28373 38887 28407
rect 24225 28169 24259 28203
rect 32781 28169 32815 28203
rect 23121 28101 23155 28135
rect 23765 28033 23799 28067
rect 31861 28033 31895 28067
rect 22569 27965 22603 27999
rect 22845 27965 22879 27999
rect 22989 27965 23023 27999
rect 31677 27965 31711 27999
rect 31769 27965 31803 27999
rect 31953 27965 31987 27999
rect 32137 27965 32171 27999
rect 22753 27897 22787 27931
rect 30941 27829 30975 27863
rect 31493 27829 31527 27863
rect 33333 27829 33367 27863
rect 1777 27557 1811 27591
rect 22477 27557 22511 27591
rect 1961 27489 1995 27523
rect 2605 27489 2639 27523
rect 31125 27421 31159 27455
rect 34437 27081 34471 27115
rect 4077 26877 4111 26911
rect 30021 26877 30055 26911
rect 34345 26877 34379 26911
rect 30297 26809 30331 26843
rect 29469 26741 29503 26775
rect 31769 26741 31803 26775
rect 32689 26741 32723 26775
rect 35081 26741 35115 26775
rect 32229 26537 32263 26571
rect 2968 26401 3002 26435
rect 3065 26401 3099 26435
rect 3157 26401 3191 26435
rect 3341 26401 3375 26435
rect 3985 26333 4019 26367
rect 2789 26265 2823 26299
rect 4537 26265 4571 26299
rect 3893 25653 3927 25687
rect 45937 25653 45971 25687
rect 46489 25381 46523 25415
rect 46397 25313 46431 25347
rect 46581 25313 46615 25347
rect 46765 25313 46799 25347
rect 47501 25313 47535 25347
rect 48145 25313 48179 25347
rect 45201 25109 45235 25143
rect 46213 25109 46247 25143
rect 47961 25109 47995 25143
rect 46121 24905 46155 24939
rect 39773 24701 39807 24735
rect 40601 24701 40635 24735
rect 45569 24701 45603 24735
rect 28549 24633 28583 24667
rect 40233 24633 40267 24667
rect 27997 24565 28031 24599
rect 29837 24565 29871 24599
rect 19717 24361 19751 24395
rect 36093 24293 36127 24327
rect 18889 24225 18923 24259
rect 35725 24225 35759 24259
rect 18613 24157 18647 24191
rect 17509 24021 17543 24055
rect 35541 23749 35575 23783
rect 25789 23273 25823 23307
rect 25881 23137 25915 23171
rect 26433 22933 26467 22967
rect 1777 22457 1811 22491
rect 1961 22457 1995 22491
rect 2605 22389 2639 22423
rect 26525 22049 26559 22083
rect 27241 22049 27275 22083
rect 26985 21981 27019 22015
rect 28365 21913 28399 21947
rect 29009 21845 29043 21879
rect 27629 20213 27663 20247
rect 26893 20009 26927 20043
rect 27261 19941 27295 19975
rect 30941 19941 30975 19975
rect 32505 19941 32539 19975
rect 27077 19873 27111 19907
rect 29745 19873 29779 19907
rect 31125 19873 31159 19907
rect 31493 19873 31527 19907
rect 31953 19805 31987 19839
rect 27905 19669 27939 19703
rect 29561 19669 29595 19703
rect 5089 19329 5123 19363
rect 3433 19261 3467 19295
rect 3801 19261 3835 19295
rect 4537 19261 4571 19295
rect 2973 19193 3007 19227
rect 3617 19193 3651 19227
rect 3709 19193 3743 19227
rect 3985 19125 4019 19159
rect 4537 18581 4571 18615
rect 14197 18037 14231 18071
rect 12265 17833 12299 17867
rect 15117 17765 15151 17799
rect 1961 17697 1995 17731
rect 13553 17629 13587 17663
rect 13829 17629 13863 17663
rect 14841 17629 14875 17663
rect 16589 17629 16623 17663
rect 17233 17561 17267 17595
rect 1869 17493 1903 17527
rect 2605 17493 2639 17527
rect 17785 17493 17819 17527
rect 40509 17289 40543 17323
rect 41889 17085 41923 17119
rect 14013 17017 14047 17051
rect 41644 17017 41678 17051
rect 39865 16949 39899 16983
rect 27721 16541 27755 16575
rect 18153 16201 18187 16235
rect 17417 15861 17451 15895
rect 17233 15657 17267 15691
rect 17969 15589 18003 15623
rect 18061 15589 18095 15623
rect 17877 15521 17911 15555
rect 18245 15521 18279 15555
rect 17693 15385 17727 15419
rect 18153 15113 18187 15147
rect 17693 15045 17727 15079
rect 19073 15045 19107 15079
rect 17141 14773 17175 14807
rect 18000 14501 18034 14535
rect 19073 14501 19107 14535
rect 18245 14365 18279 14399
rect 16037 14229 16071 14263
rect 16865 14229 16899 14263
rect 14841 14025 14875 14059
rect 40509 15861 40543 15895
rect 40785 15589 40819 15623
rect 42165 15453 42199 15487
rect 42441 15453 42475 15487
rect 40693 15113 40727 15147
rect 14105 13957 14139 13991
rect 15209 13957 15243 13991
rect 15347 13957 15381 13991
rect 27721 13957 27755 13991
rect 12081 13889 12115 13923
rect 15117 13889 15151 13923
rect 15945 13889 15979 13923
rect 17693 13889 17727 13923
rect 18153 13889 18187 13923
rect 12348 13821 12382 13855
rect 17141 13821 17175 13855
rect 17877 13821 17911 13855
rect 15485 13753 15519 13787
rect 18245 13753 18279 13787
rect 13461 13685 13495 13719
rect 16405 13481 16439 13515
rect 37473 13413 37507 13447
rect 15761 13141 15795 13175
rect 17693 13141 17727 13175
rect 18245 13141 18279 13175
rect 38669 12937 38703 12971
rect 37473 12733 37507 12767
rect 38393 12733 38427 12767
rect 39221 12733 39255 12767
rect 1869 12393 1903 12427
rect 11345 12393 11379 12427
rect 1961 12257 1995 12291
rect 2605 12053 2639 12087
rect 12265 11849 12299 11883
rect 43545 11849 43579 11883
rect 45661 11849 45695 11883
rect 10793 11781 10827 11815
rect 44373 11713 44407 11747
rect 10241 11645 10275 11679
rect 44097 11645 44131 11679
rect 10609 11577 10643 11611
rect 11713 11577 11747 11611
rect 10425 11509 10459 11543
rect 10517 11509 10551 11543
rect 11069 11305 11103 11339
rect 38761 11305 38795 11339
rect 43729 11305 43763 11339
rect 38117 11237 38151 11271
rect 38301 11237 38335 11271
rect 37933 11101 37967 11135
rect 37933 10761 37967 10795
rect 38025 9333 38059 9367
rect 47501 8993 47535 9027
rect 48145 8993 48179 9027
rect 47961 8789 47995 8823
rect 38025 8585 38059 8619
rect 18153 8245 18187 8279
rect 17417 8041 17451 8075
rect 38209 8041 38243 8075
rect 38301 8041 38335 8075
rect 39589 8041 39623 8075
rect 42165 8041 42199 8075
rect 44281 8041 44315 8075
rect 37933 7973 37967 8007
rect 38117 7973 38151 8007
rect 38485 7973 38519 8007
rect 39037 7973 39071 8007
rect 18061 7905 18095 7939
rect 18153 7905 18187 7939
rect 42993 7905 43027 7939
rect 42717 7837 42751 7871
rect 17969 7769 18003 7803
rect 38025 7497 38059 7531
rect 38945 7497 38979 7531
rect 39497 7497 39531 7531
rect 40601 7497 40635 7531
rect 1777 7429 1811 7463
rect 42441 7429 42475 7463
rect 39681 7361 39715 7395
rect 39957 7361 39991 7395
rect 17325 7293 17359 7327
rect 18245 7293 18279 7327
rect 39773 7293 39807 7327
rect 39865 7293 39899 7327
rect 1961 7225 1995 7259
rect 17969 7225 18003 7259
rect 39129 6953 39163 6987
rect 39681 6953 39715 6987
rect 18153 6613 18187 6647
rect 6929 6409 6963 6443
rect 7573 6409 7607 6443
rect 38025 6409 38059 6443
rect 6837 6205 6871 6239
rect 18245 6069 18279 6103
rect 38485 6069 38519 6103
rect 18245 5865 18279 5899
rect 38025 5865 38059 5899
rect 17601 5729 17635 5763
rect 17785 5729 17819 5763
rect 18061 5729 18095 5763
rect 38117 5729 38151 5763
rect 38577 5729 38611 5763
rect 17141 5661 17175 5695
rect 17877 5661 17911 5695
rect 17969 5593 18003 5627
rect 38485 5321 38519 5355
rect 17693 5253 17727 5287
rect 37933 5117 37967 5151
rect 38117 5117 38151 5151
rect 38301 5117 38335 5151
rect 38209 5049 38243 5083
rect 18245 4981 18279 5015
rect 39037 4981 39071 5015
rect 18245 4777 18279 4811
rect 38025 4777 38059 4811
rect 38025 4233 38059 4267
rect 43545 4097 43579 4131
rect 44189 4097 44223 4131
rect 41613 3961 41647 3995
rect 41061 3689 41095 3723
rect 41613 3689 41647 3723
rect 42809 3689 42843 3723
rect 43361 3689 43395 3723
rect 44465 3689 44499 3723
rect 42165 3553 42199 3587
rect 42349 3553 42383 3587
rect 42533 3553 42567 3587
rect 42625 3553 42659 3587
rect 44649 3553 44683 3587
rect 44925 3553 44959 3587
rect 43913 3485 43947 3519
rect 44741 3485 44775 3519
rect 42441 3417 42475 3451
rect 44833 3417 44867 3451
rect 10609 3145 10643 3179
rect 41245 3145 41279 3179
rect 41797 3077 41831 3111
rect 43361 3009 43395 3043
rect 44741 3009 44775 3043
rect 45569 3009 45603 3043
rect 10701 2941 10735 2975
rect 45017 2941 45051 2975
rect 37933 2805 37967 2839
rect 1593 2601 1627 2635
rect 10885 2601 10919 2635
rect 38117 2601 38151 2635
rect 43269 2601 43303 2635
rect 1409 2465 1443 2499
rect 2053 2465 2087 2499
rect 37933 2465 37967 2499
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 9246 47354
rect 9298 47302 9310 47354
rect 9362 47302 9374 47354
rect 9426 47302 9438 47354
rect 9490 47302 19246 47354
rect 19298 47302 19310 47354
rect 19362 47302 19374 47354
rect 19426 47302 19438 47354
rect 19490 47302 29246 47354
rect 29298 47302 29310 47354
rect 29362 47302 29374 47354
rect 29426 47302 29438 47354
rect 29490 47302 39246 47354
rect 39298 47302 39310 47354
rect 39362 47302 39374 47354
rect 39426 47302 39438 47354
rect 39490 47302 48852 47354
rect 1104 47280 48852 47302
rect 1854 47240 1860 47252
rect 1815 47212 1860 47240
rect 1854 47200 1860 47212
rect 1912 47200 1918 47252
rect 1949 47107 2007 47113
rect 1949 47073 1961 47107
rect 1995 47104 2007 47107
rect 2593 47107 2651 47113
rect 2593 47104 2605 47107
rect 1995 47076 2605 47104
rect 1995 47073 2007 47076
rect 1949 47067 2007 47073
rect 2593 47073 2605 47076
rect 2639 47104 2651 47107
rect 17310 47104 17316 47116
rect 2639 47076 17316 47104
rect 2639 47073 2651 47076
rect 2593 47067 2651 47073
rect 17310 47064 17316 47076
rect 17368 47064 17374 47116
rect 1104 46810 48852 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 14246 46810
rect 14298 46758 14310 46810
rect 14362 46758 14374 46810
rect 14426 46758 14438 46810
rect 14490 46758 24246 46810
rect 24298 46758 24310 46810
rect 24362 46758 24374 46810
rect 24426 46758 24438 46810
rect 24490 46758 34246 46810
rect 34298 46758 34310 46810
rect 34362 46758 34374 46810
rect 34426 46758 34438 46810
rect 34490 46758 44246 46810
rect 44298 46758 44310 46810
rect 44362 46758 44374 46810
rect 44426 46758 44438 46810
rect 44490 46758 48852 46810
rect 1104 46736 48852 46758
rect 1104 46266 48852 46288
rect 1104 46214 9246 46266
rect 9298 46214 9310 46266
rect 9362 46214 9374 46266
rect 9426 46214 9438 46266
rect 9490 46214 19246 46266
rect 19298 46214 19310 46266
rect 19362 46214 19374 46266
rect 19426 46214 19438 46266
rect 19490 46214 29246 46266
rect 29298 46214 29310 46266
rect 29362 46214 29374 46266
rect 29426 46214 29438 46266
rect 29490 46214 39246 46266
rect 39298 46214 39310 46266
rect 39362 46214 39374 46266
rect 39426 46214 39438 46266
rect 39490 46214 48852 46266
rect 1104 46192 48852 46214
rect 1104 45722 48852 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 14246 45722
rect 14298 45670 14310 45722
rect 14362 45670 14374 45722
rect 14426 45670 14438 45722
rect 14490 45670 24246 45722
rect 24298 45670 24310 45722
rect 24362 45670 24374 45722
rect 24426 45670 24438 45722
rect 24490 45670 34246 45722
rect 34298 45670 34310 45722
rect 34362 45670 34374 45722
rect 34426 45670 34438 45722
rect 34490 45670 44246 45722
rect 44298 45670 44310 45722
rect 44362 45670 44374 45722
rect 44426 45670 44438 45722
rect 44490 45670 48852 45722
rect 1104 45648 48852 45670
rect 19978 45432 19984 45484
rect 20036 45472 20042 45484
rect 22741 45475 22799 45481
rect 22741 45472 22753 45475
rect 20036 45444 22753 45472
rect 20036 45432 20042 45444
rect 22741 45441 22753 45444
rect 22787 45472 22799 45475
rect 24857 45475 24915 45481
rect 24857 45472 24869 45475
rect 22787 45444 24869 45472
rect 22787 45441 22799 45444
rect 22741 45435 22799 45441
rect 24857 45441 24869 45444
rect 24903 45441 24915 45475
rect 24857 45435 24915 45441
rect 23017 45407 23075 45413
rect 23017 45404 23029 45407
rect 22848 45376 23029 45404
rect 2866 45228 2872 45280
rect 2924 45268 2930 45280
rect 22189 45271 22247 45277
rect 22189 45268 22201 45271
rect 2924 45240 22201 45268
rect 2924 45228 2930 45240
rect 22189 45237 22201 45240
rect 22235 45268 22247 45271
rect 22848 45268 22876 45376
rect 23017 45373 23029 45376
rect 23063 45373 23075 45407
rect 23017 45367 23075 45373
rect 24397 45339 24455 45345
rect 24397 45305 24409 45339
rect 24443 45336 24455 45339
rect 25774 45336 25780 45348
rect 24443 45308 25780 45336
rect 24443 45305 24455 45308
rect 24397 45299 24455 45305
rect 25774 45296 25780 45308
rect 25832 45296 25838 45348
rect 22235 45240 22876 45268
rect 22235 45237 22247 45240
rect 22189 45231 22247 45237
rect 1104 45178 48852 45200
rect 1104 45126 9246 45178
rect 9298 45126 9310 45178
rect 9362 45126 9374 45178
rect 9426 45126 9438 45178
rect 9490 45126 19246 45178
rect 19298 45126 19310 45178
rect 19362 45126 19374 45178
rect 19426 45126 19438 45178
rect 19490 45126 29246 45178
rect 29298 45126 29310 45178
rect 29362 45126 29374 45178
rect 29426 45126 29438 45178
rect 29490 45126 39246 45178
rect 39298 45126 39310 45178
rect 39362 45126 39374 45178
rect 39426 45126 39438 45178
rect 39490 45126 48852 45178
rect 1104 45104 48852 45126
rect 1104 44634 48852 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 14246 44634
rect 14298 44582 14310 44634
rect 14362 44582 14374 44634
rect 14426 44582 14438 44634
rect 14490 44582 24246 44634
rect 24298 44582 24310 44634
rect 24362 44582 24374 44634
rect 24426 44582 24438 44634
rect 24490 44582 34246 44634
rect 34298 44582 34310 44634
rect 34362 44582 34374 44634
rect 34426 44582 34438 44634
rect 34490 44582 44246 44634
rect 44298 44582 44310 44634
rect 44362 44582 44374 44634
rect 44426 44582 44438 44634
rect 44490 44582 48852 44634
rect 1104 44560 48852 44582
rect 1104 44090 48852 44112
rect 1104 44038 9246 44090
rect 9298 44038 9310 44090
rect 9362 44038 9374 44090
rect 9426 44038 9438 44090
rect 9490 44038 19246 44090
rect 19298 44038 19310 44090
rect 19362 44038 19374 44090
rect 19426 44038 19438 44090
rect 19490 44038 29246 44090
rect 29298 44038 29310 44090
rect 29362 44038 29374 44090
rect 29426 44038 29438 44090
rect 29490 44038 39246 44090
rect 39298 44038 39310 44090
rect 39362 44038 39374 44090
rect 39426 44038 39438 44090
rect 39490 44038 48852 44090
rect 1104 44016 48852 44038
rect 1104 43546 48852 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 14246 43546
rect 14298 43494 14310 43546
rect 14362 43494 14374 43546
rect 14426 43494 14438 43546
rect 14490 43494 24246 43546
rect 24298 43494 24310 43546
rect 24362 43494 24374 43546
rect 24426 43494 24438 43546
rect 24490 43494 34246 43546
rect 34298 43494 34310 43546
rect 34362 43494 34374 43546
rect 34426 43494 34438 43546
rect 34490 43494 44246 43546
rect 44298 43494 44310 43546
rect 44362 43494 44374 43546
rect 44426 43494 44438 43546
rect 44490 43494 48852 43546
rect 1104 43472 48852 43494
rect 1104 43002 48852 43024
rect 1104 42950 9246 43002
rect 9298 42950 9310 43002
rect 9362 42950 9374 43002
rect 9426 42950 9438 43002
rect 9490 42950 19246 43002
rect 19298 42950 19310 43002
rect 19362 42950 19374 43002
rect 19426 42950 19438 43002
rect 19490 42950 29246 43002
rect 29298 42950 29310 43002
rect 29362 42950 29374 43002
rect 29426 42950 29438 43002
rect 29490 42950 39246 43002
rect 39298 42950 39310 43002
rect 39362 42950 39374 43002
rect 39426 42950 39438 43002
rect 39490 42950 48852 43002
rect 1104 42928 48852 42950
rect 39666 42761 39672 42764
rect 1949 42755 2007 42761
rect 1949 42721 1961 42755
rect 1995 42752 2007 42755
rect 39623 42755 39672 42761
rect 1995 42724 2636 42752
rect 1995 42721 2007 42724
rect 1949 42715 2007 42721
rect 1854 42548 1860 42560
rect 1815 42520 1860 42548
rect 1854 42508 1860 42520
rect 1912 42508 1918 42560
rect 2608 42557 2636 42724
rect 39623 42721 39635 42755
rect 39669 42721 39672 42755
rect 39623 42715 39672 42721
rect 39666 42712 39672 42715
rect 39724 42752 39730 42764
rect 39724 42724 40724 42752
rect 39724 42712 39730 42724
rect 35342 42644 35348 42696
rect 35400 42684 35406 42696
rect 40696 42693 40724 42724
rect 42794 42712 42800 42764
rect 42852 42752 42858 42764
rect 43605 42755 43663 42761
rect 43605 42752 43617 42755
rect 42852 42724 43617 42752
rect 42852 42712 42858 42724
rect 43605 42721 43617 42724
rect 43651 42721 43663 42755
rect 43605 42715 43663 42721
rect 39025 42687 39083 42693
rect 39025 42684 39037 42687
rect 35400 42656 39037 42684
rect 35400 42644 35406 42656
rect 39025 42653 39037 42656
rect 39071 42653 39083 42687
rect 39025 42647 39083 42653
rect 40681 42687 40739 42693
rect 40681 42653 40693 42687
rect 40727 42684 40739 42687
rect 43346 42684 43352 42696
rect 40727 42656 43024 42684
rect 43307 42656 43352 42684
rect 40727 42653 40739 42656
rect 40681 42647 40739 42653
rect 38930 42576 38936 42628
rect 38988 42616 38994 42628
rect 42996 42616 43024 42656
rect 43346 42644 43352 42656
rect 43404 42644 43410 42696
rect 43254 42616 43260 42628
rect 38988 42588 42932 42616
rect 42996 42588 43260 42616
rect 38988 42576 38994 42588
rect 2593 42551 2651 42557
rect 2593 42517 2605 42551
rect 2639 42548 2651 42551
rect 12250 42548 12256 42560
rect 2639 42520 12256 42548
rect 2639 42517 2651 42520
rect 2593 42511 2651 42517
rect 12250 42508 12256 42520
rect 12308 42508 12314 42560
rect 42794 42548 42800 42560
rect 42755 42520 42800 42548
rect 42794 42508 42800 42520
rect 42852 42508 42858 42560
rect 42904 42548 42932 42588
rect 43254 42576 43260 42588
rect 43312 42576 43318 42628
rect 44729 42551 44787 42557
rect 44729 42548 44741 42551
rect 42904 42520 44741 42548
rect 44729 42517 44741 42520
rect 44775 42517 44787 42551
rect 44729 42511 44787 42517
rect 1104 42458 48852 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 14246 42458
rect 14298 42406 14310 42458
rect 14362 42406 14374 42458
rect 14426 42406 14438 42458
rect 14490 42406 24246 42458
rect 24298 42406 24310 42458
rect 24362 42406 24374 42458
rect 24426 42406 24438 42458
rect 24490 42406 34246 42458
rect 34298 42406 34310 42458
rect 34362 42406 34374 42458
rect 34426 42406 34438 42458
rect 34490 42406 44246 42458
rect 44298 42406 44310 42458
rect 44362 42406 44374 42458
rect 44426 42406 44438 42458
rect 44490 42406 48852 42458
rect 1104 42384 48852 42406
rect 40678 41964 40684 42016
rect 40736 42004 40742 42016
rect 43165 42007 43223 42013
rect 43165 42004 43177 42007
rect 40736 41976 43177 42004
rect 40736 41964 40742 41976
rect 43165 41973 43177 41976
rect 43211 42004 43223 42007
rect 43346 42004 43352 42016
rect 43211 41976 43352 42004
rect 43211 41973 43223 41976
rect 43165 41967 43223 41973
rect 43346 41964 43352 41976
rect 43404 41964 43410 42016
rect 1104 41914 48852 41936
rect 1104 41862 9246 41914
rect 9298 41862 9310 41914
rect 9362 41862 9374 41914
rect 9426 41862 9438 41914
rect 9490 41862 19246 41914
rect 19298 41862 19310 41914
rect 19362 41862 19374 41914
rect 19426 41862 19438 41914
rect 19490 41862 29246 41914
rect 29298 41862 29310 41914
rect 29362 41862 29374 41914
rect 29426 41862 29438 41914
rect 29490 41862 39246 41914
rect 39298 41862 39310 41914
rect 39362 41862 39374 41914
rect 39426 41862 39438 41914
rect 39490 41862 48852 41914
rect 1104 41840 48852 41862
rect 7561 41735 7619 41741
rect 7561 41732 7573 41735
rect 7024 41704 7573 41732
rect 7024 41673 7052 41704
rect 7561 41701 7573 41704
rect 7607 41732 7619 41735
rect 39666 41732 39672 41744
rect 7607 41704 39672 41732
rect 7607 41701 7619 41704
rect 7561 41695 7619 41701
rect 39666 41692 39672 41704
rect 39724 41692 39730 41744
rect 7009 41667 7067 41673
rect 7009 41633 7021 41667
rect 7055 41633 7067 41667
rect 7009 41627 7067 41633
rect 12989 41667 13047 41673
rect 12989 41633 13001 41667
rect 13035 41633 13047 41667
rect 12989 41627 13047 41633
rect 13004 41528 13032 41627
rect 13078 41624 13084 41676
rect 13136 41664 13142 41676
rect 13357 41667 13415 41673
rect 13357 41664 13369 41667
rect 13136 41636 13369 41664
rect 13136 41624 13142 41636
rect 13357 41633 13369 41636
rect 13403 41633 13415 41667
rect 47949 41667 48007 41673
rect 47949 41664 47961 41667
rect 13357 41627 13415 41633
rect 47320 41636 47961 41664
rect 13630 41596 13636 41608
rect 13591 41568 13636 41596
rect 13630 41556 13636 41568
rect 13688 41556 13694 41608
rect 14369 41531 14427 41537
rect 14369 41528 14381 41531
rect 13004 41500 14381 41528
rect 14369 41497 14381 41500
rect 14415 41528 14427 41531
rect 15102 41528 15108 41540
rect 14415 41500 15108 41528
rect 14415 41497 14427 41500
rect 14369 41491 14427 41497
rect 15102 41488 15108 41500
rect 15160 41488 15166 41540
rect 6730 41460 6736 41472
rect 6691 41432 6736 41460
rect 6730 41420 6736 41432
rect 6788 41420 6794 41472
rect 44542 41420 44548 41472
rect 44600 41460 44606 41472
rect 47320 41469 47348 41636
rect 47949 41633 47961 41636
rect 47995 41633 48007 41667
rect 48130 41664 48136 41676
rect 48091 41636 48136 41664
rect 47949 41627 48007 41633
rect 48130 41624 48136 41636
rect 48188 41624 48194 41676
rect 47305 41463 47363 41469
rect 47305 41460 47317 41463
rect 44600 41432 47317 41460
rect 44600 41420 44606 41432
rect 47305 41429 47317 41432
rect 47351 41429 47363 41463
rect 47305 41423 47363 41429
rect 1104 41370 48852 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 14246 41370
rect 14298 41318 14310 41370
rect 14362 41318 14374 41370
rect 14426 41318 14438 41370
rect 14490 41318 24246 41370
rect 24298 41318 24310 41370
rect 24362 41318 24374 41370
rect 24426 41318 24438 41370
rect 24490 41318 34246 41370
rect 34298 41318 34310 41370
rect 34362 41318 34374 41370
rect 34426 41318 34438 41370
rect 34490 41318 44246 41370
rect 44298 41318 44310 41370
rect 44362 41318 44374 41370
rect 44426 41318 44438 41370
rect 44490 41318 48852 41370
rect 1104 41296 48852 41318
rect 13078 40876 13084 40928
rect 13136 40916 13142 40928
rect 13909 40919 13967 40925
rect 13909 40916 13921 40919
rect 13136 40888 13921 40916
rect 13136 40876 13142 40888
rect 13909 40885 13921 40888
rect 13955 40885 13967 40919
rect 13909 40879 13967 40885
rect 1104 40826 48852 40848
rect 1104 40774 9246 40826
rect 9298 40774 9310 40826
rect 9362 40774 9374 40826
rect 9426 40774 9438 40826
rect 9490 40774 19246 40826
rect 19298 40774 19310 40826
rect 19362 40774 19374 40826
rect 19426 40774 19438 40826
rect 19490 40774 29246 40826
rect 29298 40774 29310 40826
rect 29362 40774 29374 40826
rect 29426 40774 29438 40826
rect 29490 40774 39246 40826
rect 39298 40774 39310 40826
rect 39362 40774 39374 40826
rect 39426 40774 39438 40826
rect 39490 40774 48852 40826
rect 1104 40752 48852 40774
rect 1104 40282 48852 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 14246 40282
rect 14298 40230 14310 40282
rect 14362 40230 14374 40282
rect 14426 40230 14438 40282
rect 14490 40230 24246 40282
rect 24298 40230 24310 40282
rect 24362 40230 24374 40282
rect 24426 40230 24438 40282
rect 24490 40230 34246 40282
rect 34298 40230 34310 40282
rect 34362 40230 34374 40282
rect 34426 40230 34438 40282
rect 34490 40230 44246 40282
rect 44298 40230 44310 40282
rect 44362 40230 44374 40282
rect 44426 40230 44438 40282
rect 44490 40230 48852 40282
rect 1104 40208 48852 40230
rect 1104 39738 48852 39760
rect 1104 39686 9246 39738
rect 9298 39686 9310 39738
rect 9362 39686 9374 39738
rect 9426 39686 9438 39738
rect 9490 39686 19246 39738
rect 19298 39686 19310 39738
rect 19362 39686 19374 39738
rect 19426 39686 19438 39738
rect 19490 39686 29246 39738
rect 29298 39686 29310 39738
rect 29362 39686 29374 39738
rect 29426 39686 29438 39738
rect 29490 39686 39246 39738
rect 39298 39686 39310 39738
rect 39362 39686 39374 39738
rect 39426 39686 39438 39738
rect 39490 39686 48852 39738
rect 1104 39664 48852 39686
rect 16669 39627 16727 39633
rect 16669 39624 16681 39627
rect 16546 39596 16681 39624
rect 15102 39516 15108 39568
rect 15160 39556 15166 39568
rect 15473 39559 15531 39565
rect 15473 39556 15485 39559
rect 15160 39528 15485 39556
rect 15160 39516 15166 39528
rect 15473 39525 15485 39528
rect 15519 39525 15531 39559
rect 15473 39519 15531 39525
rect 15488 39420 15516 39519
rect 16025 39491 16083 39497
rect 16025 39457 16037 39491
rect 16071 39488 16083 39491
rect 16546 39488 16574 39596
rect 16669 39593 16681 39596
rect 16715 39624 16727 39627
rect 35342 39624 35348 39636
rect 16715 39596 35348 39624
rect 16715 39593 16727 39596
rect 16669 39587 16727 39593
rect 35342 39584 35348 39596
rect 35400 39584 35406 39636
rect 22664 39528 24256 39556
rect 22664 39497 22692 39528
rect 16071 39460 16574 39488
rect 22649 39491 22707 39497
rect 16071 39457 16083 39460
rect 16025 39451 16083 39457
rect 22649 39457 22661 39491
rect 22695 39457 22707 39491
rect 22649 39451 22707 39457
rect 22925 39491 22983 39497
rect 22925 39457 22937 39491
rect 22971 39457 22983 39491
rect 23106 39488 23112 39500
rect 23067 39460 23112 39488
rect 22925 39451 22983 39457
rect 21910 39420 21916 39432
rect 15488 39392 21916 39420
rect 21910 39380 21916 39392
rect 21968 39420 21974 39432
rect 22833 39423 22891 39429
rect 22833 39420 22845 39423
rect 21968 39392 22845 39420
rect 21968 39380 21974 39392
rect 22833 39389 22845 39392
rect 22879 39389 22891 39423
rect 22940 39420 22968 39451
rect 23106 39448 23112 39460
rect 23164 39448 23170 39500
rect 22940 39392 23704 39420
rect 22833 39383 22891 39389
rect 22738 39352 22744 39364
rect 22699 39324 22744 39352
rect 22738 39312 22744 39324
rect 22796 39312 22802 39364
rect 23676 39296 23704 39392
rect 22465 39287 22523 39293
rect 22465 39253 22477 39287
rect 22511 39284 22523 39287
rect 22554 39284 22560 39296
rect 22511 39256 22560 39284
rect 22511 39253 22523 39256
rect 22465 39247 22523 39253
rect 22554 39244 22560 39256
rect 22612 39244 22618 39296
rect 23658 39284 23664 39296
rect 23619 39256 23664 39284
rect 23658 39244 23664 39256
rect 23716 39244 23722 39296
rect 24228 39293 24256 39528
rect 24213 39287 24271 39293
rect 24213 39253 24225 39287
rect 24259 39284 24271 39287
rect 24578 39284 24584 39296
rect 24259 39256 24584 39284
rect 24259 39253 24271 39256
rect 24213 39247 24271 39253
rect 24578 39244 24584 39256
rect 24636 39244 24642 39296
rect 24762 39244 24768 39296
rect 24820 39284 24826 39296
rect 43990 39284 43996 39296
rect 24820 39256 43996 39284
rect 24820 39244 24826 39256
rect 43990 39244 43996 39256
rect 44048 39284 44054 39296
rect 44542 39284 44548 39296
rect 44048 39256 44548 39284
rect 44048 39244 44054 39256
rect 44542 39244 44548 39256
rect 44600 39244 44606 39296
rect 1104 39194 48852 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 14246 39194
rect 14298 39142 14310 39194
rect 14362 39142 14374 39194
rect 14426 39142 14438 39194
rect 14490 39142 24246 39194
rect 24298 39142 24310 39194
rect 24362 39142 24374 39194
rect 24426 39142 24438 39194
rect 24490 39142 34246 39194
rect 34298 39142 34310 39194
rect 34362 39142 34374 39194
rect 34426 39142 34438 39194
rect 34490 39142 44246 39194
rect 44298 39142 44310 39194
rect 44362 39142 44374 39194
rect 44426 39142 44438 39194
rect 44490 39142 48852 39194
rect 1104 39120 48852 39142
rect 24578 39040 24584 39092
rect 24636 39080 24642 39092
rect 39666 39080 39672 39092
rect 24636 39052 39672 39080
rect 24636 39040 24642 39052
rect 39666 39040 39672 39052
rect 39724 39040 39730 39092
rect 23658 38972 23664 39024
rect 23716 39012 23722 39024
rect 32858 39012 32864 39024
rect 23716 38984 32864 39012
rect 23716 38972 23722 38984
rect 32858 38972 32864 38984
rect 32916 38972 32922 39024
rect 24670 38876 24676 38888
rect 24631 38848 24676 38876
rect 24670 38836 24676 38848
rect 24728 38876 24734 38888
rect 25133 38879 25191 38885
rect 25133 38876 25145 38879
rect 24728 38848 25145 38876
rect 24728 38836 24734 38848
rect 25133 38845 25145 38848
rect 25179 38845 25191 38879
rect 25133 38839 25191 38845
rect 32858 38836 32864 38888
rect 32916 38876 32922 38888
rect 33502 38876 33508 38888
rect 32916 38848 33508 38876
rect 32916 38836 32922 38848
rect 33502 38836 33508 38848
rect 33560 38836 33566 38888
rect 24762 38808 24768 38820
rect 23584 38780 24768 38808
rect 22738 38700 22744 38752
rect 22796 38740 22802 38752
rect 23584 38749 23612 38780
rect 24762 38768 24768 38780
rect 24820 38768 24826 38820
rect 33226 38808 33232 38820
rect 33187 38780 33232 38808
rect 33226 38768 33232 38780
rect 33284 38768 33290 38820
rect 23569 38743 23627 38749
rect 23569 38740 23581 38743
rect 22796 38712 23581 38740
rect 22796 38700 22802 38712
rect 23569 38709 23581 38712
rect 23615 38709 23627 38743
rect 23569 38703 23627 38709
rect 23934 38700 23940 38752
rect 23992 38740 23998 38752
rect 24581 38743 24639 38749
rect 24581 38740 24593 38743
rect 23992 38712 24593 38740
rect 23992 38700 23998 38712
rect 24581 38709 24593 38712
rect 24627 38709 24639 38743
rect 29086 38740 29092 38752
rect 29047 38712 29092 38740
rect 24581 38703 24639 38709
rect 29086 38700 29092 38712
rect 29144 38700 29150 38752
rect 1104 38650 48852 38672
rect 1104 38598 9246 38650
rect 9298 38598 9310 38650
rect 9362 38598 9374 38650
rect 9426 38598 9438 38650
rect 9490 38598 19246 38650
rect 19298 38598 19310 38650
rect 19362 38598 19374 38650
rect 19426 38598 19438 38650
rect 19490 38598 29246 38650
rect 29298 38598 29310 38650
rect 29362 38598 29374 38650
rect 29426 38598 29438 38650
rect 29490 38598 39246 38650
rect 39298 38598 39310 38650
rect 39362 38598 39374 38650
rect 39426 38598 39438 38650
rect 39490 38598 48852 38650
rect 1104 38576 48852 38598
rect 32858 38536 32864 38548
rect 32819 38508 32864 38536
rect 32858 38496 32864 38508
rect 32916 38496 32922 38548
rect 10045 38471 10103 38477
rect 10045 38437 10057 38471
rect 10091 38468 10103 38471
rect 16942 38468 16948 38480
rect 10091 38440 16948 38468
rect 10091 38437 10103 38440
rect 10045 38431 10103 38437
rect 16942 38428 16948 38440
rect 17000 38428 17006 38480
rect 5166 38400 5172 38412
rect 5127 38372 5172 38400
rect 5166 38360 5172 38372
rect 5224 38400 5230 38412
rect 6089 38403 6147 38409
rect 6089 38400 6101 38403
rect 5224 38372 6101 38400
rect 5224 38360 5230 38372
rect 6089 38369 6101 38372
rect 6135 38369 6147 38403
rect 6089 38363 6147 38369
rect 9953 38403 10011 38409
rect 9953 38369 9965 38403
rect 9999 38369 10011 38403
rect 9953 38363 10011 38369
rect 5445 38335 5503 38341
rect 5445 38301 5457 38335
rect 5491 38332 5503 38335
rect 9858 38332 9864 38344
rect 5491 38304 9864 38332
rect 5491 38301 5503 38304
rect 5445 38295 5503 38301
rect 9858 38292 9864 38304
rect 9916 38292 9922 38344
rect 9968 38332 9996 38363
rect 24118 38360 24124 38412
rect 24176 38400 24182 38412
rect 28353 38403 28411 38409
rect 28353 38400 28365 38403
rect 24176 38372 28365 38400
rect 24176 38360 24182 38372
rect 28353 38369 28365 38372
rect 28399 38400 28411 38403
rect 28813 38403 28871 38409
rect 28813 38400 28825 38403
rect 28399 38372 28825 38400
rect 28399 38369 28411 38372
rect 28353 38363 28411 38369
rect 28813 38369 28825 38372
rect 28859 38369 28871 38403
rect 28813 38363 28871 38369
rect 10597 38335 10655 38341
rect 10597 38332 10609 38335
rect 9968 38304 10609 38332
rect 10597 38301 10609 38304
rect 10643 38332 10655 38335
rect 27985 38335 28043 38341
rect 27985 38332 27997 38335
rect 10643 38304 27997 38332
rect 10643 38301 10655 38304
rect 10597 38295 10655 38301
rect 27985 38301 27997 38304
rect 28031 38332 28043 38335
rect 29086 38332 29092 38344
rect 28031 38304 29092 38332
rect 28031 38301 28043 38304
rect 27985 38295 28043 38301
rect 29086 38292 29092 38304
rect 29144 38292 29150 38344
rect 28215 38267 28273 38273
rect 28215 38233 28227 38267
rect 28261 38264 28273 38267
rect 28261 38236 29040 38264
rect 28261 38233 28273 38236
rect 28215 38227 28273 38233
rect 29012 38208 29040 38236
rect 27706 38196 27712 38208
rect 27667 38168 27712 38196
rect 27706 38156 27712 38168
rect 27764 38156 27770 38208
rect 28074 38196 28080 38208
rect 28035 38168 28080 38196
rect 28074 38156 28080 38168
rect 28132 38156 28138 38208
rect 28994 38156 29000 38208
rect 29052 38196 29058 38208
rect 29365 38199 29423 38205
rect 29365 38196 29377 38199
rect 29052 38168 29377 38196
rect 29052 38156 29058 38168
rect 29365 38165 29377 38168
rect 29411 38165 29423 38199
rect 29365 38159 29423 38165
rect 1104 38106 48852 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 14246 38106
rect 14298 38054 14310 38106
rect 14362 38054 14374 38106
rect 14426 38054 14438 38106
rect 14490 38054 24246 38106
rect 24298 38054 24310 38106
rect 24362 38054 24374 38106
rect 24426 38054 24438 38106
rect 24490 38054 34246 38106
rect 34298 38054 34310 38106
rect 34362 38054 34374 38106
rect 34426 38054 34438 38106
rect 34490 38054 44246 38106
rect 44298 38054 44310 38106
rect 44362 38054 44374 38106
rect 44426 38054 44438 38106
rect 44490 38054 48852 38106
rect 1104 38032 48852 38054
rect 29086 37884 29092 37936
rect 29144 37924 29150 37936
rect 42058 37924 42064 37936
rect 29144 37896 42064 37924
rect 29144 37884 29150 37896
rect 42058 37884 42064 37896
rect 42116 37884 42122 37936
rect 28074 37612 28080 37664
rect 28132 37652 28138 37664
rect 28905 37655 28963 37661
rect 28905 37652 28917 37655
rect 28132 37624 28917 37652
rect 28132 37612 28138 37624
rect 28905 37621 28917 37624
rect 28951 37652 28963 37655
rect 39114 37652 39120 37664
rect 28951 37624 39120 37652
rect 28951 37621 28963 37624
rect 28905 37615 28963 37621
rect 39114 37612 39120 37624
rect 39172 37612 39178 37664
rect 1104 37562 48852 37584
rect 1104 37510 9246 37562
rect 9298 37510 9310 37562
rect 9362 37510 9374 37562
rect 9426 37510 9438 37562
rect 9490 37510 19246 37562
rect 19298 37510 19310 37562
rect 19362 37510 19374 37562
rect 19426 37510 19438 37562
rect 19490 37510 29246 37562
rect 29298 37510 29310 37562
rect 29362 37510 29374 37562
rect 29426 37510 29438 37562
rect 29490 37510 39246 37562
rect 39298 37510 39310 37562
rect 39362 37510 39374 37562
rect 39426 37510 39438 37562
rect 39490 37510 48852 37562
rect 1104 37488 48852 37510
rect 1854 37448 1860 37460
rect 1815 37420 1860 37448
rect 1854 37408 1860 37420
rect 1912 37408 1918 37460
rect 1949 37315 2007 37321
rect 1949 37281 1961 37315
rect 1995 37312 2007 37315
rect 2593 37315 2651 37321
rect 2593 37312 2605 37315
rect 1995 37284 2605 37312
rect 1995 37281 2007 37284
rect 1949 37275 2007 37281
rect 2593 37281 2605 37284
rect 2639 37312 2651 37315
rect 38930 37312 38936 37324
rect 2639 37284 38936 37312
rect 2639 37281 2651 37284
rect 2593 37275 2651 37281
rect 38930 37272 38936 37284
rect 38988 37272 38994 37324
rect 1104 37018 48852 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 14246 37018
rect 14298 36966 14310 37018
rect 14362 36966 14374 37018
rect 14426 36966 14438 37018
rect 14490 36966 24246 37018
rect 24298 36966 24310 37018
rect 24362 36966 24374 37018
rect 24426 36966 24438 37018
rect 24490 36966 34246 37018
rect 34298 36966 34310 37018
rect 34362 36966 34374 37018
rect 34426 36966 34438 37018
rect 34490 36966 44246 37018
rect 44298 36966 44310 37018
rect 44362 36966 44374 37018
rect 44426 36966 44438 37018
rect 44490 36966 48852 37018
rect 1104 36944 48852 36966
rect 17589 36907 17647 36913
rect 17589 36904 17601 36907
rect 16546 36876 17601 36904
rect 11698 36796 11704 36848
rect 11756 36836 11762 36848
rect 15013 36839 15071 36845
rect 15013 36836 15025 36839
rect 11756 36808 15025 36836
rect 11756 36796 11762 36808
rect 15013 36805 15025 36808
rect 15059 36805 15071 36839
rect 15013 36799 15071 36805
rect 16393 36771 16451 36777
rect 16393 36737 16405 36771
rect 16439 36768 16451 36771
rect 16546 36768 16574 36876
rect 17589 36873 17601 36876
rect 17635 36904 17647 36907
rect 19978 36904 19984 36916
rect 17635 36876 19984 36904
rect 17635 36873 17647 36876
rect 17589 36867 17647 36873
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 16439 36740 16574 36768
rect 16439 36737 16451 36740
rect 16393 36731 16451 36737
rect 16148 36635 16206 36641
rect 16148 36601 16160 36635
rect 16194 36632 16206 36635
rect 16194 36604 16574 36632
rect 16194 36601 16206 36604
rect 16148 36595 16206 36601
rect 13354 36564 13360 36576
rect 13315 36536 13360 36564
rect 13354 36524 13360 36536
rect 13412 36524 13418 36576
rect 16546 36564 16574 36604
rect 17034 36564 17040 36576
rect 16546 36536 17040 36564
rect 17034 36524 17040 36536
rect 17092 36524 17098 36576
rect 1104 36474 48852 36496
rect 1104 36422 9246 36474
rect 9298 36422 9310 36474
rect 9362 36422 9374 36474
rect 9426 36422 9438 36474
rect 9490 36422 19246 36474
rect 19298 36422 19310 36474
rect 19362 36422 19374 36474
rect 19426 36422 19438 36474
rect 19490 36422 29246 36474
rect 29298 36422 29310 36474
rect 29362 36422 29374 36474
rect 29426 36422 29438 36474
rect 29490 36422 39246 36474
rect 39298 36422 39310 36474
rect 39362 36422 39374 36474
rect 39426 36422 39438 36474
rect 39490 36422 48852 36474
rect 1104 36400 48852 36422
rect 9858 36320 9864 36372
rect 9916 36360 9922 36372
rect 11701 36363 11759 36369
rect 11701 36360 11713 36363
rect 9916 36332 11713 36360
rect 9916 36320 9922 36332
rect 11701 36329 11713 36332
rect 11747 36329 11759 36363
rect 11701 36323 11759 36329
rect 12268 36332 16574 36360
rect 11716 36224 11744 36323
rect 12268 36233 12296 36332
rect 12437 36295 12495 36301
rect 12437 36261 12449 36295
rect 12483 36292 12495 36295
rect 16546 36292 16574 36332
rect 17034 36320 17040 36372
rect 17092 36360 17098 36372
rect 35066 36360 35072 36372
rect 17092 36332 35072 36360
rect 17092 36320 17098 36332
rect 35066 36320 35072 36332
rect 35124 36320 35130 36372
rect 21358 36292 21364 36304
rect 12483 36264 13492 36292
rect 16546 36264 21364 36292
rect 12483 36261 12495 36264
rect 12437 36255 12495 36261
rect 12253 36227 12311 36233
rect 12253 36224 12265 36227
rect 11716 36196 12265 36224
rect 12253 36193 12265 36196
rect 12299 36193 12311 36227
rect 12526 36224 12532 36236
rect 12487 36196 12532 36224
rect 12253 36187 12311 36193
rect 12526 36184 12532 36196
rect 12584 36184 12590 36236
rect 12673 36227 12731 36233
rect 12673 36193 12685 36227
rect 12719 36224 12731 36227
rect 13354 36224 13360 36236
rect 12719 36196 13360 36224
rect 12719 36193 12731 36196
rect 12673 36187 12731 36193
rect 13354 36184 13360 36196
rect 13412 36184 13418 36236
rect 13464 36165 13492 36264
rect 21358 36252 21364 36264
rect 21416 36252 21422 36304
rect 13449 36159 13507 36165
rect 13449 36125 13461 36159
rect 13495 36156 13507 36159
rect 24118 36156 24124 36168
rect 13495 36128 24124 36156
rect 13495 36125 13507 36128
rect 13449 36119 13507 36125
rect 24118 36116 24124 36128
rect 24176 36116 24182 36168
rect 12805 36091 12863 36097
rect 12805 36057 12817 36091
rect 12851 36088 12863 36091
rect 12851 36060 16574 36088
rect 12851 36057 12863 36060
rect 12805 36051 12863 36057
rect 16546 36020 16574 36060
rect 40770 36020 40776 36032
rect 16546 35992 40776 36020
rect 40770 35980 40776 35992
rect 40828 35980 40834 36032
rect 1104 35930 48852 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 14246 35930
rect 14298 35878 14310 35930
rect 14362 35878 14374 35930
rect 14426 35878 14438 35930
rect 14490 35878 24246 35930
rect 24298 35878 24310 35930
rect 24362 35878 24374 35930
rect 24426 35878 24438 35930
rect 24490 35878 34246 35930
rect 34298 35878 34310 35930
rect 34362 35878 34374 35930
rect 34426 35878 34438 35930
rect 34490 35878 44246 35930
rect 44298 35878 44310 35930
rect 44362 35878 44374 35930
rect 44426 35878 44438 35930
rect 44490 35878 48852 35930
rect 1104 35856 48852 35878
rect 47213 35615 47271 35621
rect 47213 35581 47225 35615
rect 47259 35612 47271 35615
rect 47670 35612 47676 35624
rect 47259 35584 47676 35612
rect 47259 35581 47271 35584
rect 47213 35575 47271 35581
rect 47670 35572 47676 35584
rect 47728 35572 47734 35624
rect 47765 35547 47823 35553
rect 47765 35544 47777 35547
rect 45526 35516 47777 35544
rect 12526 35436 12532 35488
rect 12584 35476 12590 35488
rect 13265 35479 13323 35485
rect 13265 35476 13277 35479
rect 12584 35448 13277 35476
rect 12584 35436 12590 35448
rect 13265 35445 13277 35448
rect 13311 35476 13323 35479
rect 21542 35476 21548 35488
rect 13311 35448 21548 35476
rect 13311 35445 13323 35448
rect 13265 35439 13323 35445
rect 21542 35436 21548 35448
rect 21600 35476 21606 35488
rect 28994 35476 29000 35488
rect 21600 35448 29000 35476
rect 21600 35436 21606 35448
rect 28994 35436 29000 35448
rect 29052 35436 29058 35488
rect 39666 35436 39672 35488
rect 39724 35476 39730 35488
rect 45526 35476 45554 35516
rect 47765 35513 47777 35516
rect 47811 35513 47823 35547
rect 47765 35507 47823 35513
rect 39724 35448 45554 35476
rect 39724 35436 39730 35448
rect 1104 35386 48852 35408
rect 1104 35334 9246 35386
rect 9298 35334 9310 35386
rect 9362 35334 9374 35386
rect 9426 35334 9438 35386
rect 9490 35334 19246 35386
rect 19298 35334 19310 35386
rect 19362 35334 19374 35386
rect 19426 35334 19438 35386
rect 19490 35334 29246 35386
rect 29298 35334 29310 35386
rect 29362 35334 29374 35386
rect 29426 35334 29438 35386
rect 29490 35334 39246 35386
rect 39298 35334 39310 35386
rect 39362 35334 39374 35386
rect 39426 35334 39438 35386
rect 39490 35334 48852 35386
rect 1104 35312 48852 35334
rect 1104 34842 48852 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 14246 34842
rect 14298 34790 14310 34842
rect 14362 34790 14374 34842
rect 14426 34790 14438 34842
rect 14490 34790 24246 34842
rect 24298 34790 24310 34842
rect 24362 34790 24374 34842
rect 24426 34790 24438 34842
rect 24490 34790 34246 34842
rect 34298 34790 34310 34842
rect 34362 34790 34374 34842
rect 34426 34790 34438 34842
rect 34490 34790 44246 34842
rect 44298 34790 44310 34842
rect 44362 34790 44374 34842
rect 44426 34790 44438 34842
rect 44490 34790 48852 34842
rect 1104 34768 48852 34790
rect 39022 34484 39028 34536
rect 39080 34524 39086 34536
rect 39666 34524 39672 34536
rect 39080 34496 39672 34524
rect 39080 34484 39086 34496
rect 39666 34484 39672 34496
rect 39724 34484 39730 34536
rect 1104 34298 48852 34320
rect 1104 34246 9246 34298
rect 9298 34246 9310 34298
rect 9362 34246 9374 34298
rect 9426 34246 9438 34298
rect 9490 34246 19246 34298
rect 19298 34246 19310 34298
rect 19362 34246 19374 34298
rect 19426 34246 19438 34298
rect 19490 34246 29246 34298
rect 29298 34246 29310 34298
rect 29362 34246 29374 34298
rect 29426 34246 29438 34298
rect 29490 34246 39246 34298
rect 39298 34246 39310 34298
rect 39362 34246 39374 34298
rect 39426 34246 39438 34298
rect 39490 34246 48852 34298
rect 1104 34224 48852 34246
rect 10410 34048 10416 34060
rect 10371 34020 10416 34048
rect 10410 34008 10416 34020
rect 10468 34048 10474 34060
rect 10873 34051 10931 34057
rect 10873 34048 10885 34051
rect 10468 34020 10885 34048
rect 10468 34008 10474 34020
rect 10873 34017 10885 34020
rect 10919 34017 10931 34051
rect 10873 34011 10931 34017
rect 10229 33983 10287 33989
rect 10229 33949 10241 33983
rect 10275 33980 10287 33983
rect 17402 33980 17408 33992
rect 10275 33952 17408 33980
rect 10275 33949 10287 33952
rect 10229 33943 10287 33949
rect 17402 33940 17408 33952
rect 17460 33940 17466 33992
rect 38194 33844 38200 33856
rect 38155 33816 38200 33844
rect 38194 33804 38200 33816
rect 38252 33804 38258 33856
rect 1104 33754 48852 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 14246 33754
rect 14298 33702 14310 33754
rect 14362 33702 14374 33754
rect 14426 33702 14438 33754
rect 14490 33702 24246 33754
rect 24298 33702 24310 33754
rect 24362 33702 24374 33754
rect 24426 33702 24438 33754
rect 24490 33702 34246 33754
rect 34298 33702 34310 33754
rect 34362 33702 34374 33754
rect 34426 33702 34438 33754
rect 34490 33702 44246 33754
rect 44298 33702 44310 33754
rect 44362 33702 44374 33754
rect 44426 33702 44438 33754
rect 44490 33702 48852 33754
rect 1104 33680 48852 33702
rect 39117 33575 39175 33581
rect 39117 33572 39129 33575
rect 26206 33544 39129 33572
rect 18322 33396 18328 33448
rect 18380 33436 18386 33448
rect 26206 33436 26234 33544
rect 39117 33541 39129 33544
rect 39163 33541 39175 33575
rect 39117 33535 39175 33541
rect 39666 33504 39672 33516
rect 38856 33476 39672 33504
rect 38856 33445 38884 33476
rect 39666 33464 39672 33476
rect 39724 33464 39730 33516
rect 18380 33408 26234 33436
rect 38821 33439 38884 33445
rect 18380 33396 18386 33408
rect 38821 33405 38833 33439
rect 38867 33408 38884 33439
rect 38867 33405 38879 33408
rect 38821 33399 38879 33405
rect 28258 33328 28264 33380
rect 28316 33368 28322 33380
rect 38194 33368 38200 33380
rect 28316 33340 38200 33368
rect 28316 33328 28322 33340
rect 38194 33328 38200 33340
rect 38252 33368 38258 33380
rect 38565 33371 38623 33377
rect 38565 33368 38577 33371
rect 38252 33340 38577 33368
rect 38252 33328 38258 33340
rect 38565 33337 38577 33340
rect 38611 33337 38623 33371
rect 38565 33331 38623 33337
rect 38731 33371 38789 33377
rect 38731 33337 38743 33371
rect 38777 33368 38789 33371
rect 38933 33371 38991 33377
rect 38777 33337 38792 33368
rect 38731 33331 38792 33337
rect 38933 33337 38945 33371
rect 38979 33337 38991 33371
rect 38933 33331 38991 33337
rect 38105 33303 38163 33309
rect 38105 33269 38117 33303
rect 38151 33300 38163 33303
rect 38286 33300 38292 33312
rect 38151 33272 38292 33300
rect 38151 33269 38163 33272
rect 38105 33263 38163 33269
rect 38286 33260 38292 33272
rect 38344 33300 38350 33312
rect 38764 33300 38792 33331
rect 38344 33272 38792 33300
rect 38948 33300 38976 33331
rect 39574 33300 39580 33312
rect 38948 33272 39580 33300
rect 38344 33260 38350 33272
rect 39574 33260 39580 33272
rect 39632 33260 39638 33312
rect 39666 33260 39672 33312
rect 39724 33300 39730 33312
rect 40129 33303 40187 33309
rect 40129 33300 40141 33303
rect 39724 33272 40141 33300
rect 39724 33260 39730 33272
rect 40129 33269 40141 33272
rect 40175 33269 40187 33303
rect 47026 33300 47032 33312
rect 46987 33272 47032 33300
rect 40129 33263 40187 33269
rect 47026 33260 47032 33272
rect 47084 33260 47090 33312
rect 1104 33210 48852 33232
rect 1104 33158 9246 33210
rect 9298 33158 9310 33210
rect 9362 33158 9374 33210
rect 9426 33158 9438 33210
rect 9490 33158 19246 33210
rect 19298 33158 19310 33210
rect 19362 33158 19374 33210
rect 19426 33158 19438 33210
rect 19490 33158 29246 33210
rect 29298 33158 29310 33210
rect 29362 33158 29374 33210
rect 29426 33158 29438 33210
rect 29490 33158 39246 33210
rect 39298 33158 39310 33210
rect 39362 33158 39374 33210
rect 39426 33158 39438 33210
rect 39490 33158 48852 33210
rect 1104 33136 48852 33158
rect 33134 33056 33140 33108
rect 33192 33096 33198 33108
rect 37921 33099 37979 33105
rect 37921 33096 37933 33099
rect 33192 33068 37933 33096
rect 33192 33056 33198 33068
rect 37921 33065 37933 33068
rect 37967 33096 37979 33099
rect 37967 33068 38792 33096
rect 37967 33065 37979 33068
rect 37921 33059 37979 33065
rect 38764 33028 38792 33068
rect 47029 33031 47087 33037
rect 47029 33028 47041 33031
rect 38764 33000 47041 33028
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 30469 32963 30527 32969
rect 30469 32960 30481 32963
rect 29788 32932 30481 32960
rect 29788 32920 29794 32932
rect 30469 32929 30481 32932
rect 30515 32929 30527 32963
rect 30469 32923 30527 32929
rect 38470 32920 38476 32972
rect 38528 32969 38534 32972
rect 38764 32969 38792 33000
rect 47029 32997 47041 33000
rect 47075 33028 47087 33031
rect 47949 33031 48007 33037
rect 47949 33028 47961 33031
rect 47075 33000 47961 33028
rect 47075 32997 47087 33000
rect 47029 32991 47087 32997
rect 47949 32997 47961 33000
rect 47995 32997 48007 33031
rect 47949 32991 48007 32997
rect 38528 32960 38537 32969
rect 38749 32963 38807 32969
rect 38528 32932 38573 32960
rect 38528 32923 38537 32932
rect 38749 32929 38761 32963
rect 38795 32929 38807 32963
rect 47719 32963 47777 32969
rect 47719 32960 47731 32963
rect 38749 32923 38807 32929
rect 47044 32932 47731 32960
rect 38528 32920 38534 32923
rect 47044 32904 47072 32932
rect 47719 32929 47731 32932
rect 47765 32929 47777 32963
rect 47854 32960 47860 32972
rect 47815 32932 47860 32960
rect 47719 32923 47777 32929
rect 47854 32920 47860 32932
rect 47912 32920 47918 32972
rect 48133 32963 48191 32969
rect 48133 32929 48145 32963
rect 48179 32929 48191 32963
rect 48133 32923 48191 32929
rect 38010 32852 38016 32904
rect 38068 32892 38074 32904
rect 38565 32895 38623 32901
rect 38565 32892 38577 32895
rect 38068 32864 38577 32892
rect 38068 32852 38074 32864
rect 38565 32861 38577 32864
rect 38611 32861 38623 32895
rect 38565 32855 38623 32861
rect 38667 32895 38725 32901
rect 38667 32861 38679 32895
rect 38713 32892 38725 32895
rect 39485 32895 39543 32901
rect 39485 32892 39497 32895
rect 38713 32864 39497 32892
rect 38713 32861 38725 32864
rect 38667 32855 38725 32861
rect 39485 32861 39497 32864
rect 39531 32892 39543 32895
rect 39758 32892 39764 32904
rect 39531 32864 39764 32892
rect 39531 32861 39543 32864
rect 39485 32855 39543 32861
rect 39758 32852 39764 32864
rect 39816 32852 39822 32904
rect 47026 32852 47032 32904
rect 47084 32852 47090 32904
rect 38933 32827 38991 32833
rect 38933 32793 38945 32827
rect 38979 32824 38991 32827
rect 42702 32824 42708 32836
rect 38979 32796 42708 32824
rect 38979 32793 38991 32796
rect 38933 32787 38991 32793
rect 42702 32784 42708 32796
rect 42760 32784 42766 32836
rect 48148 32824 48176 32923
rect 46768 32796 48176 32824
rect 46768 32768 46796 32796
rect 30653 32759 30711 32765
rect 30653 32725 30665 32759
rect 30699 32756 30711 32759
rect 32398 32756 32404 32768
rect 30699 32728 32404 32756
rect 30699 32725 30711 32728
rect 30653 32719 30711 32725
rect 32398 32716 32404 32728
rect 32456 32716 32462 32768
rect 38470 32716 38476 32768
rect 38528 32756 38534 32768
rect 40037 32759 40095 32765
rect 40037 32756 40049 32759
rect 38528 32728 40049 32756
rect 38528 32716 38534 32728
rect 40037 32725 40049 32728
rect 40083 32756 40095 32759
rect 40494 32756 40500 32768
rect 40083 32728 40500 32756
rect 40083 32725 40095 32728
rect 40037 32719 40095 32725
rect 40494 32716 40500 32728
rect 40552 32716 40558 32768
rect 46569 32759 46627 32765
rect 46569 32725 46581 32759
rect 46615 32756 46627 32759
rect 46750 32756 46756 32768
rect 46615 32728 46756 32756
rect 46615 32725 46627 32728
rect 46569 32719 46627 32725
rect 46750 32716 46756 32728
rect 46808 32716 46814 32768
rect 47578 32756 47584 32768
rect 47539 32728 47584 32756
rect 47578 32716 47584 32728
rect 47636 32716 47642 32768
rect 1104 32666 48852 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 14246 32666
rect 14298 32614 14310 32666
rect 14362 32614 14374 32666
rect 14426 32614 14438 32666
rect 14490 32614 24246 32666
rect 24298 32614 24310 32666
rect 24362 32614 24374 32666
rect 24426 32614 24438 32666
rect 24490 32614 34246 32666
rect 34298 32614 34310 32666
rect 34362 32614 34374 32666
rect 34426 32614 34438 32666
rect 34490 32614 44246 32666
rect 44298 32614 44310 32666
rect 44362 32614 44374 32666
rect 44426 32614 44438 32666
rect 44490 32614 48852 32666
rect 1104 32592 48852 32614
rect 24670 32512 24676 32564
rect 24728 32552 24734 32564
rect 45554 32552 45560 32564
rect 24728 32524 45560 32552
rect 24728 32512 24734 32524
rect 45554 32512 45560 32524
rect 45612 32552 45618 32564
rect 47213 32555 47271 32561
rect 47213 32552 47225 32555
rect 45612 32524 47225 32552
rect 45612 32512 45618 32524
rect 47213 32521 47225 32524
rect 47259 32552 47271 32555
rect 47854 32552 47860 32564
rect 47259 32524 47860 32552
rect 47259 32521 47271 32524
rect 47213 32515 47271 32521
rect 47854 32512 47860 32524
rect 47912 32512 47918 32564
rect 1762 32416 1768 32428
rect 1723 32388 1768 32416
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 40678 32416 40684 32428
rect 40639 32388 40684 32416
rect 40678 32376 40684 32388
rect 40736 32376 40742 32428
rect 38746 32348 38752 32360
rect 26206 32320 38752 32348
rect 1949 32283 2007 32289
rect 1949 32249 1961 32283
rect 1995 32280 2007 32283
rect 2593 32283 2651 32289
rect 2593 32280 2605 32283
rect 1995 32252 2605 32280
rect 1995 32249 2007 32252
rect 1949 32243 2007 32249
rect 2593 32249 2605 32252
rect 2639 32280 2651 32283
rect 26206 32280 26234 32320
rect 38746 32308 38752 32320
rect 38804 32308 38810 32360
rect 40414 32283 40472 32289
rect 40414 32280 40426 32283
rect 2639 32252 26234 32280
rect 38672 32252 40426 32280
rect 2639 32249 2651 32252
rect 2593 32243 2651 32249
rect 38672 32224 38700 32252
rect 40414 32249 40426 32252
rect 40460 32249 40472 32283
rect 40414 32243 40472 32249
rect 37274 32172 37280 32224
rect 37332 32212 37338 32224
rect 38010 32212 38016 32224
rect 37332 32184 38016 32212
rect 37332 32172 37338 32184
rect 38010 32172 38016 32184
rect 38068 32172 38074 32224
rect 38654 32212 38660 32224
rect 38615 32184 38660 32212
rect 38654 32172 38660 32184
rect 38712 32172 38718 32224
rect 38746 32172 38752 32224
rect 38804 32212 38810 32224
rect 39301 32215 39359 32221
rect 39301 32212 39313 32215
rect 38804 32184 39313 32212
rect 38804 32172 38810 32184
rect 39301 32181 39313 32184
rect 39347 32212 39359 32215
rect 39942 32212 39948 32224
rect 39347 32184 39948 32212
rect 39347 32181 39359 32184
rect 39301 32175 39359 32181
rect 39942 32172 39948 32184
rect 40000 32172 40006 32224
rect 1104 32122 48852 32144
rect 1104 32070 9246 32122
rect 9298 32070 9310 32122
rect 9362 32070 9374 32122
rect 9426 32070 9438 32122
rect 9490 32070 19246 32122
rect 19298 32070 19310 32122
rect 19362 32070 19374 32122
rect 19426 32070 19438 32122
rect 19490 32070 29246 32122
rect 29298 32070 29310 32122
rect 29362 32070 29374 32122
rect 29426 32070 29438 32122
rect 29490 32070 39246 32122
rect 39298 32070 39310 32122
rect 39362 32070 39374 32122
rect 39426 32070 39438 32122
rect 39490 32070 48852 32122
rect 1104 32048 48852 32070
rect 21542 32008 21548 32020
rect 20824 31980 21548 32008
rect 20824 31881 20852 31980
rect 21542 31968 21548 31980
rect 21600 31968 21606 32020
rect 41046 32008 41052 32020
rect 26206 31980 41052 32008
rect 20901 31943 20959 31949
rect 20901 31909 20913 31943
rect 20947 31940 20959 31943
rect 26206 31940 26234 31980
rect 41046 31968 41052 31980
rect 41104 31968 41110 32020
rect 20947 31912 26234 31940
rect 20947 31909 20959 31912
rect 20901 31903 20959 31909
rect 39114 31900 39120 31952
rect 39172 31900 39178 31952
rect 20809 31875 20867 31881
rect 20809 31841 20821 31875
rect 20855 31841 20867 31875
rect 38930 31872 38936 31884
rect 38891 31844 38936 31872
rect 20809 31835 20867 31841
rect 38930 31832 38936 31844
rect 38988 31832 38994 31884
rect 39132 31872 39160 31900
rect 39209 31875 39267 31881
rect 39209 31872 39221 31875
rect 39132 31844 39221 31872
rect 39209 31841 39221 31844
rect 39255 31872 39267 31875
rect 39850 31872 39856 31884
rect 39255 31844 39856 31872
rect 39255 31841 39267 31844
rect 39209 31835 39267 31841
rect 39850 31832 39856 31844
rect 39908 31832 39914 31884
rect 3142 31804 3148 31816
rect 3103 31776 3148 31804
rect 3142 31764 3148 31776
rect 3200 31764 3206 31816
rect 38286 31804 38292 31816
rect 38247 31776 38292 31804
rect 38286 31764 38292 31776
rect 38344 31804 38350 31816
rect 39025 31807 39083 31813
rect 39025 31804 39037 31807
rect 38344 31776 39037 31804
rect 38344 31764 38350 31776
rect 39025 31773 39037 31776
rect 39071 31773 39083 31807
rect 39025 31767 39083 31773
rect 39114 31764 39120 31816
rect 39172 31804 39178 31816
rect 39393 31807 39451 31813
rect 39172 31776 39217 31804
rect 39172 31764 39178 31776
rect 39393 31773 39405 31807
rect 39439 31804 39451 31807
rect 41230 31804 41236 31816
rect 39439 31776 41236 31804
rect 39439 31773 39451 31776
rect 39393 31767 39451 31773
rect 41230 31764 41236 31776
rect 41288 31764 41294 31816
rect 38654 31736 38660 31748
rect 6886 31708 38660 31736
rect 1762 31628 1768 31680
rect 1820 31668 1826 31680
rect 6886 31668 6914 31708
rect 38654 31696 38660 31708
rect 38712 31696 38718 31748
rect 39132 31736 39160 31764
rect 39666 31736 39672 31748
rect 39132 31708 39672 31736
rect 39666 31696 39672 31708
rect 39724 31696 39730 31748
rect 1820 31640 6914 31668
rect 1820 31628 1826 31640
rect 1104 31578 48852 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 14246 31578
rect 14298 31526 14310 31578
rect 14362 31526 14374 31578
rect 14426 31526 14438 31578
rect 14490 31526 24246 31578
rect 24298 31526 24310 31578
rect 24362 31526 24374 31578
rect 24426 31526 24438 31578
rect 24490 31526 34246 31578
rect 34298 31526 34310 31578
rect 34362 31526 34374 31578
rect 34426 31526 34438 31578
rect 34490 31526 44246 31578
rect 44298 31526 44310 31578
rect 44362 31526 44374 31578
rect 44426 31526 44438 31578
rect 44490 31526 48852 31578
rect 1104 31504 48852 31526
rect 1762 31464 1768 31476
rect 1723 31436 1768 31464
rect 1762 31424 1768 31436
rect 1820 31424 1826 31476
rect 38930 31424 38936 31476
rect 38988 31464 38994 31476
rect 39669 31467 39727 31473
rect 39669 31464 39681 31467
rect 38988 31436 39681 31464
rect 38988 31424 38994 31436
rect 39669 31433 39681 31436
rect 39715 31433 39727 31467
rect 39669 31427 39727 31433
rect 3142 31396 3148 31408
rect 1964 31368 3148 31396
rect 1964 31269 1992 31368
rect 3142 31356 3148 31368
rect 3200 31396 3206 31408
rect 3200 31368 6914 31396
rect 3200 31356 3206 31368
rect 2133 31331 2191 31337
rect 2133 31297 2145 31331
rect 2179 31328 2191 31331
rect 3513 31331 3571 31337
rect 3513 31328 3525 31331
rect 2179 31300 3525 31328
rect 2179 31297 2191 31300
rect 2133 31291 2191 31297
rect 3513 31297 3525 31300
rect 3559 31328 3571 31331
rect 6886 31328 6914 31368
rect 38378 31356 38384 31408
rect 38436 31396 38442 31408
rect 39117 31399 39175 31405
rect 39117 31396 39129 31399
rect 38436 31368 39129 31396
rect 38436 31356 38442 31368
rect 39117 31365 39129 31368
rect 39163 31396 39175 31399
rect 40678 31396 40684 31408
rect 39163 31368 40684 31396
rect 39163 31365 39175 31368
rect 39117 31359 39175 31365
rect 40678 31356 40684 31368
rect 40736 31356 40742 31408
rect 25682 31328 25688 31340
rect 3559 31300 4200 31328
rect 6886 31300 25688 31328
rect 3559 31297 3571 31300
rect 3513 31291 3571 31297
rect 1949 31263 2007 31269
rect 1949 31229 1961 31263
rect 1995 31229 2007 31263
rect 1949 31223 2007 31229
rect 2041 31263 2099 31269
rect 2041 31229 2053 31263
rect 2087 31229 2099 31263
rect 2222 31260 2228 31272
rect 2183 31232 2228 31260
rect 2041 31223 2099 31229
rect 2056 31192 2084 31223
rect 2222 31220 2228 31232
rect 2280 31220 2286 31272
rect 2409 31263 2467 31269
rect 2409 31229 2421 31263
rect 2455 31260 2467 31263
rect 4062 31260 4068 31272
rect 2455 31232 4068 31260
rect 2455 31229 2467 31232
rect 2409 31223 2467 31229
rect 4062 31220 4068 31232
rect 4120 31220 4126 31272
rect 4172 31260 4200 31300
rect 25682 31288 25688 31300
rect 25740 31288 25746 31340
rect 15654 31260 15660 31272
rect 4172 31232 15660 31260
rect 15654 31220 15660 31232
rect 15712 31220 15718 31272
rect 2961 31195 3019 31201
rect 2961 31192 2973 31195
rect 2056 31164 2973 31192
rect 2961 31161 2973 31164
rect 3007 31192 3019 31195
rect 38565 31195 38623 31201
rect 3007 31164 6914 31192
rect 3007 31161 3019 31164
rect 2961 31155 3019 31161
rect 4062 31124 4068 31136
rect 4023 31096 4068 31124
rect 4062 31084 4068 31096
rect 4120 31084 4126 31136
rect 6886 31124 6914 31164
rect 38565 31161 38577 31195
rect 38611 31192 38623 31195
rect 39114 31192 39120 31204
rect 38611 31164 39120 31192
rect 38611 31161 38623 31164
rect 38565 31155 38623 31161
rect 39114 31152 39120 31164
rect 39172 31152 39178 31204
rect 21910 31124 21916 31136
rect 6886 31096 21916 31124
rect 21910 31084 21916 31096
rect 21968 31084 21974 31136
rect 1104 31034 48852 31056
rect 1104 30982 9246 31034
rect 9298 30982 9310 31034
rect 9362 30982 9374 31034
rect 9426 30982 9438 31034
rect 9490 30982 19246 31034
rect 19298 30982 19310 31034
rect 19362 30982 19374 31034
rect 19426 30982 19438 31034
rect 19490 30982 29246 31034
rect 29298 30982 29310 31034
rect 29362 30982 29374 31034
rect 29426 30982 29438 31034
rect 29490 30982 39246 31034
rect 39298 30982 39310 31034
rect 39362 30982 39374 31034
rect 39426 30982 39438 31034
rect 39490 30982 48852 31034
rect 1104 30960 48852 30982
rect 4062 30880 4068 30932
rect 4120 30920 4126 30932
rect 37458 30920 37464 30932
rect 4120 30892 37464 30920
rect 4120 30880 4126 30892
rect 37458 30880 37464 30892
rect 37516 30880 37522 30932
rect 15654 30852 15660 30864
rect 15615 30824 15660 30852
rect 15654 30812 15660 30824
rect 15712 30852 15718 30864
rect 31846 30852 31852 30864
rect 15712 30824 31852 30852
rect 15712 30812 15718 30824
rect 31846 30812 31852 30824
rect 31904 30812 31910 30864
rect 15933 30787 15991 30793
rect 15933 30753 15945 30787
rect 15979 30784 15991 30787
rect 16393 30787 16451 30793
rect 16393 30784 16405 30787
rect 15979 30756 16405 30784
rect 15979 30753 15991 30756
rect 15933 30747 15991 30753
rect 16393 30753 16405 30756
rect 16439 30784 16451 30787
rect 34333 30787 34391 30793
rect 16439 30756 16574 30784
rect 16439 30753 16451 30756
rect 16393 30747 16451 30753
rect 2222 30540 2228 30592
rect 2280 30580 2286 30592
rect 2958 30580 2964 30592
rect 2280 30552 2964 30580
rect 2280 30540 2286 30552
rect 2958 30540 2964 30552
rect 3016 30540 3022 30592
rect 16546 30580 16574 30756
rect 34333 30753 34345 30787
rect 34379 30784 34391 30787
rect 47578 30784 47584 30796
rect 34379 30756 47584 30784
rect 34379 30753 34391 30756
rect 34333 30747 34391 30753
rect 47578 30744 47584 30756
rect 47636 30744 47642 30796
rect 32398 30676 32404 30728
rect 32456 30716 32462 30728
rect 32493 30719 32551 30725
rect 32493 30716 32505 30719
rect 32456 30688 32505 30716
rect 32456 30676 32462 30688
rect 32493 30685 32505 30688
rect 32539 30716 32551 30719
rect 34609 30719 34667 30725
rect 34609 30716 34621 30719
rect 32539 30688 34621 30716
rect 32539 30685 32551 30688
rect 32493 30679 32551 30685
rect 34609 30685 34621 30688
rect 34655 30716 34667 30719
rect 38378 30716 38384 30728
rect 34655 30688 38384 30716
rect 34655 30685 34667 30688
rect 34609 30679 34667 30685
rect 38378 30676 38384 30688
rect 38436 30676 38442 30728
rect 22738 30580 22744 30592
rect 16546 30552 22744 30580
rect 22738 30540 22744 30552
rect 22796 30540 22802 30592
rect 33134 30540 33140 30592
rect 33192 30580 33198 30592
rect 33229 30583 33287 30589
rect 33229 30580 33241 30583
rect 33192 30552 33241 30580
rect 33192 30540 33198 30552
rect 33229 30549 33241 30552
rect 33275 30549 33287 30583
rect 33229 30543 33287 30549
rect 1104 30490 48852 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 14246 30490
rect 14298 30438 14310 30490
rect 14362 30438 14374 30490
rect 14426 30438 14438 30490
rect 14490 30438 24246 30490
rect 24298 30438 24310 30490
rect 24362 30438 24374 30490
rect 24426 30438 24438 30490
rect 24490 30438 34246 30490
rect 34298 30438 34310 30490
rect 34362 30438 34374 30490
rect 34426 30438 34438 30490
rect 34490 30438 44246 30490
rect 44298 30438 44310 30490
rect 44362 30438 44374 30490
rect 44426 30438 44438 30490
rect 44490 30438 48852 30490
rect 1104 30416 48852 30438
rect 2958 30336 2964 30388
rect 3016 30376 3022 30388
rect 18230 30376 18236 30388
rect 3016 30348 18236 30376
rect 3016 30336 3022 30348
rect 18230 30336 18236 30348
rect 18288 30336 18294 30388
rect 35066 30308 35072 30320
rect 35027 30280 35072 30308
rect 35066 30268 35072 30280
rect 35124 30268 35130 30320
rect 35342 30308 35348 30320
rect 35303 30280 35348 30308
rect 35342 30268 35348 30280
rect 35400 30308 35406 30320
rect 36173 30311 36231 30317
rect 36173 30308 36185 30311
rect 35400 30280 36185 30308
rect 35400 30268 35406 30280
rect 36173 30277 36185 30280
rect 36219 30308 36231 30311
rect 44082 30308 44088 30320
rect 36219 30280 44088 30308
rect 36219 30277 36231 30280
rect 36173 30271 36231 30277
rect 44082 30268 44088 30280
rect 44140 30268 44146 30320
rect 33502 30240 33508 30252
rect 33415 30212 33508 30240
rect 33502 30200 33508 30212
rect 33560 30240 33566 30252
rect 33560 30212 35756 30240
rect 33560 30200 33566 30212
rect 35618 30181 35624 30184
rect 35229 30175 35287 30181
rect 35229 30172 35241 30175
rect 33980 30144 35241 30172
rect 33980 30113 34008 30144
rect 35229 30141 35241 30144
rect 35275 30141 35287 30175
rect 35229 30135 35287 30141
rect 35437 30175 35495 30181
rect 35437 30141 35449 30175
rect 35483 30141 35495 30175
rect 35437 30135 35495 30141
rect 35574 30175 35624 30181
rect 35574 30141 35586 30175
rect 35620 30141 35624 30175
rect 35574 30135 35624 30141
rect 33965 30107 34023 30113
rect 33965 30104 33977 30107
rect 26206 30076 33977 30104
rect 6914 29996 6920 30048
rect 6972 30036 6978 30048
rect 26206 30036 26234 30076
rect 33965 30073 33977 30076
rect 34011 30073 34023 30107
rect 33965 30067 34023 30073
rect 6972 30008 26234 30036
rect 6972 29996 6978 30008
rect 31846 29996 31852 30048
rect 31904 30036 31910 30048
rect 34517 30039 34575 30045
rect 34517 30036 34529 30039
rect 31904 30008 34529 30036
rect 31904 29996 31910 30008
rect 34517 30005 34529 30008
rect 34563 30036 34575 30039
rect 35452 30036 35480 30135
rect 35618 30132 35624 30135
rect 35676 30132 35682 30184
rect 35728 30181 35756 30212
rect 39574 30200 39580 30252
rect 39632 30240 39638 30252
rect 39758 30240 39764 30252
rect 39632 30212 39764 30240
rect 39632 30200 39638 30212
rect 39758 30200 39764 30212
rect 39816 30200 39822 30252
rect 43254 30200 43260 30252
rect 43312 30240 43318 30252
rect 45373 30243 45431 30249
rect 45373 30240 45385 30243
rect 43312 30212 45385 30240
rect 43312 30200 43318 30212
rect 45373 30209 45385 30212
rect 45419 30209 45431 30243
rect 45373 30203 45431 30209
rect 35713 30175 35771 30181
rect 35713 30141 35725 30175
rect 35759 30141 35771 30175
rect 45002 30172 45008 30184
rect 44963 30144 45008 30172
rect 35713 30135 35771 30141
rect 45002 30132 45008 30144
rect 45060 30132 45066 30184
rect 45465 30175 45523 30181
rect 45465 30141 45477 30175
rect 45511 30141 45523 30175
rect 45465 30135 45523 30141
rect 34563 30008 35480 30036
rect 34563 30005 34575 30008
rect 34517 29999 34575 30005
rect 39850 29996 39856 30048
rect 39908 30036 39914 30048
rect 44453 30039 44511 30045
rect 44453 30036 44465 30039
rect 39908 30008 44465 30036
rect 39908 29996 39914 30008
rect 44453 30005 44465 30008
rect 44499 30036 44511 30039
rect 45480 30036 45508 30135
rect 44499 30008 45508 30036
rect 44499 30005 44511 30008
rect 44453 29999 44511 30005
rect 1104 29946 48852 29968
rect 1104 29894 9246 29946
rect 9298 29894 9310 29946
rect 9362 29894 9374 29946
rect 9426 29894 9438 29946
rect 9490 29894 19246 29946
rect 19298 29894 19310 29946
rect 19362 29894 19374 29946
rect 19426 29894 19438 29946
rect 19490 29894 29246 29946
rect 29298 29894 29310 29946
rect 29362 29894 29374 29946
rect 29426 29894 29438 29946
rect 29490 29894 39246 29946
rect 39298 29894 39310 29946
rect 39362 29894 39374 29946
rect 39426 29894 39438 29946
rect 39490 29894 48852 29946
rect 1104 29872 48852 29894
rect 10686 29792 10692 29844
rect 10744 29832 10750 29844
rect 33502 29832 33508 29844
rect 10744 29804 33508 29832
rect 10744 29792 10750 29804
rect 33502 29792 33508 29804
rect 33560 29792 33566 29844
rect 43990 29832 43996 29844
rect 43951 29804 43996 29832
rect 43990 29792 43996 29804
rect 44048 29792 44054 29844
rect 10410 29656 10416 29708
rect 10468 29696 10474 29708
rect 25961 29699 26019 29705
rect 25961 29696 25973 29699
rect 10468 29668 25973 29696
rect 10468 29656 10474 29668
rect 25961 29665 25973 29668
rect 26007 29696 26019 29699
rect 26007 29668 26740 29696
rect 26007 29665 26019 29668
rect 25961 29659 26019 29665
rect 23106 29588 23112 29640
rect 23164 29628 23170 29640
rect 25593 29631 25651 29637
rect 25593 29628 25605 29631
rect 23164 29600 25605 29628
rect 23164 29588 23170 29600
rect 25593 29597 25605 29600
rect 25639 29597 25651 29631
rect 25774 29628 25780 29640
rect 25735 29600 25780 29628
rect 25593 29591 25651 29597
rect 25774 29588 25780 29600
rect 25832 29588 25838 29640
rect 25869 29631 25927 29637
rect 25869 29597 25881 29631
rect 25915 29597 25927 29631
rect 26050 29628 26056 29640
rect 26011 29600 26056 29628
rect 25869 29591 25927 29597
rect 25133 29563 25191 29569
rect 25133 29529 25145 29563
rect 25179 29560 25191 29563
rect 25792 29560 25820 29588
rect 25179 29532 25820 29560
rect 25884 29560 25912 29591
rect 26050 29588 26056 29600
rect 26108 29588 26114 29640
rect 26712 29569 26740 29668
rect 37550 29628 37556 29640
rect 31726 29600 37556 29628
rect 26697 29563 26755 29569
rect 25884 29532 26234 29560
rect 25179 29529 25191 29532
rect 25133 29523 25191 29529
rect 26206 29492 26234 29532
rect 26697 29529 26709 29563
rect 26743 29560 26755 29563
rect 31726 29560 31754 29600
rect 37550 29588 37556 29600
rect 37608 29628 37614 29640
rect 44637 29631 44695 29637
rect 44637 29628 44649 29631
rect 37608 29600 44649 29628
rect 37608 29588 37614 29600
rect 44637 29597 44649 29600
rect 44683 29628 44695 29631
rect 45002 29628 45008 29640
rect 44683 29600 45008 29628
rect 44683 29597 44695 29600
rect 44637 29591 44695 29597
rect 45002 29588 45008 29600
rect 45060 29588 45066 29640
rect 26743 29532 31754 29560
rect 26743 29529 26755 29532
rect 26697 29523 26755 29529
rect 42702 29520 42708 29572
rect 42760 29560 42766 29572
rect 45186 29560 45192 29572
rect 42760 29532 45192 29560
rect 42760 29520 42766 29532
rect 45186 29520 45192 29532
rect 45244 29520 45250 29572
rect 27249 29495 27307 29501
rect 27249 29492 27261 29495
rect 26206 29464 27261 29492
rect 27249 29461 27261 29464
rect 27295 29492 27307 29495
rect 30834 29492 30840 29504
rect 27295 29464 30840 29492
rect 27295 29461 27307 29464
rect 27249 29455 27307 29461
rect 30834 29452 30840 29464
rect 30892 29452 30898 29504
rect 33778 29452 33784 29504
rect 33836 29492 33842 29504
rect 34701 29495 34759 29501
rect 34701 29492 34713 29495
rect 33836 29464 34713 29492
rect 33836 29452 33842 29464
rect 34701 29461 34713 29464
rect 34747 29492 34759 29495
rect 35618 29492 35624 29504
rect 34747 29464 35624 29492
rect 34747 29461 34759 29464
rect 34701 29455 34759 29461
rect 35618 29452 35624 29464
rect 35676 29452 35682 29504
rect 37274 29452 37280 29504
rect 37332 29492 37338 29504
rect 44542 29492 44548 29504
rect 37332 29464 44548 29492
rect 37332 29452 37338 29464
rect 44542 29452 44548 29464
rect 44600 29452 44606 29504
rect 1104 29402 48852 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 14246 29402
rect 14298 29350 14310 29402
rect 14362 29350 14374 29402
rect 14426 29350 14438 29402
rect 14490 29350 24246 29402
rect 24298 29350 24310 29402
rect 24362 29350 24374 29402
rect 24426 29350 24438 29402
rect 24490 29350 34246 29402
rect 34298 29350 34310 29402
rect 34362 29350 34374 29402
rect 34426 29350 34438 29402
rect 34490 29350 44246 29402
rect 44298 29350 44310 29402
rect 44362 29350 44374 29402
rect 44426 29350 44438 29402
rect 44490 29350 48852 29402
rect 1104 29328 48852 29350
rect 44082 29288 44088 29300
rect 44043 29260 44088 29288
rect 44082 29248 44088 29260
rect 44140 29248 44146 29300
rect 43990 29180 43996 29232
rect 44048 29220 44054 29232
rect 44913 29223 44971 29229
rect 44913 29220 44925 29223
rect 44048 29192 44925 29220
rect 44048 29180 44054 29192
rect 44913 29189 44925 29192
rect 44959 29189 44971 29223
rect 44913 29183 44971 29189
rect 44082 29112 44088 29164
rect 44140 29152 44146 29164
rect 44821 29155 44879 29161
rect 44821 29152 44833 29155
rect 44140 29124 44833 29152
rect 44140 29112 44146 29124
rect 44821 29121 44833 29124
rect 44867 29121 44879 29155
rect 44821 29115 44879 29121
rect 35618 29044 35624 29096
rect 35676 29084 35682 29096
rect 44174 29084 44180 29096
rect 35676 29056 44180 29084
rect 35676 29044 35682 29056
rect 44174 29044 44180 29056
rect 44232 29044 44238 29096
rect 44542 29044 44548 29096
rect 44600 29084 44606 29096
rect 44729 29087 44787 29093
rect 44729 29084 44741 29087
rect 44600 29056 44741 29084
rect 44600 29044 44606 29056
rect 44729 29053 44741 29056
rect 44775 29053 44787 29087
rect 44729 29047 44787 29053
rect 45005 29087 45063 29093
rect 45005 29053 45017 29087
rect 45051 29053 45063 29087
rect 45186 29084 45192 29096
rect 45147 29056 45192 29084
rect 45005 29047 45063 29053
rect 25038 28976 25044 29028
rect 25096 29016 25102 29028
rect 25225 29019 25283 29025
rect 25225 29016 25237 29019
rect 25096 28988 25237 29016
rect 25096 28976 25102 28988
rect 25225 28985 25237 28988
rect 25271 29016 25283 29019
rect 26050 29016 26056 29028
rect 25271 28988 26056 29016
rect 25271 28985 25283 28988
rect 25225 28979 25283 28985
rect 26050 28976 26056 28988
rect 26108 28976 26114 29028
rect 30834 28976 30840 29028
rect 30892 29016 30898 29028
rect 39574 29016 39580 29028
rect 30892 28988 39580 29016
rect 30892 28976 30898 28988
rect 39574 28976 39580 28988
rect 39632 28976 39638 29028
rect 44192 29016 44220 29044
rect 45020 29016 45048 29047
rect 45186 29044 45192 29056
rect 45244 29044 45250 29096
rect 43916 28988 44128 29016
rect 44192 28988 45048 29016
rect 41690 28908 41696 28960
rect 41748 28948 41754 28960
rect 43916 28948 43944 28988
rect 41748 28920 43944 28948
rect 44100 28948 44128 28988
rect 44545 28951 44603 28957
rect 44545 28948 44557 28951
rect 44100 28920 44557 28948
rect 41748 28908 41754 28920
rect 44545 28917 44557 28920
rect 44591 28917 44603 28951
rect 44545 28911 44603 28917
rect 1104 28858 48852 28880
rect 1104 28806 9246 28858
rect 9298 28806 9310 28858
rect 9362 28806 9374 28858
rect 9426 28806 9438 28858
rect 9490 28806 19246 28858
rect 19298 28806 19310 28858
rect 19362 28806 19374 28858
rect 19426 28806 19438 28858
rect 19490 28806 29246 28858
rect 29298 28806 29310 28858
rect 29362 28806 29374 28858
rect 29426 28806 29438 28858
rect 29490 28806 39246 28858
rect 39298 28806 39310 28858
rect 39362 28806 39374 28858
rect 39426 28806 39438 28858
rect 39490 28806 48852 28858
rect 1104 28784 48852 28806
rect 21358 28704 21364 28756
rect 21416 28744 21422 28756
rect 22002 28744 22008 28756
rect 21416 28716 22008 28744
rect 21416 28704 21422 28716
rect 22002 28704 22008 28716
rect 22060 28744 22066 28756
rect 22189 28747 22247 28753
rect 22189 28744 22201 28747
rect 22060 28716 22201 28744
rect 22060 28704 22066 28716
rect 22189 28713 22201 28716
rect 22235 28713 22247 28747
rect 22189 28707 22247 28713
rect 31021 28747 31079 28753
rect 31021 28713 31033 28747
rect 31067 28744 31079 28747
rect 31846 28744 31852 28756
rect 31067 28716 31852 28744
rect 31067 28713 31079 28716
rect 31021 28707 31079 28713
rect 31846 28704 31852 28716
rect 31904 28704 31910 28756
rect 36265 28747 36323 28753
rect 36265 28713 36277 28747
rect 36311 28744 36323 28747
rect 38378 28744 38384 28756
rect 36311 28716 38384 28744
rect 36311 28713 36323 28716
rect 36265 28707 36323 28713
rect 38378 28704 38384 28716
rect 38436 28704 38442 28756
rect 44174 28744 44180 28756
rect 44135 28716 44180 28744
rect 44174 28704 44180 28716
rect 44232 28704 44238 28756
rect 23014 28568 23020 28620
rect 23072 28608 23078 28620
rect 47026 28608 47032 28620
rect 23072 28580 47032 28608
rect 23072 28568 23078 28580
rect 47026 28568 47032 28580
rect 47084 28568 47090 28620
rect 32674 28500 32680 28552
rect 32732 28540 32738 28552
rect 37366 28540 37372 28552
rect 32732 28512 37372 28540
rect 32732 28500 32738 28512
rect 37366 28500 37372 28512
rect 37424 28500 37430 28552
rect 38102 28540 38108 28552
rect 38063 28512 38108 28540
rect 38102 28500 38108 28512
rect 38160 28500 38166 28552
rect 38378 28540 38384 28552
rect 38339 28512 38384 28540
rect 38378 28500 38384 28512
rect 38436 28500 38442 28552
rect 28994 28432 29000 28484
rect 29052 28472 29058 28484
rect 29052 28444 37044 28472
rect 29052 28432 29058 28444
rect 18230 28364 18236 28416
rect 18288 28404 18294 28416
rect 24854 28404 24860 28416
rect 18288 28376 24860 28404
rect 18288 28364 18294 28376
rect 24854 28364 24860 28376
rect 24912 28364 24918 28416
rect 37016 28413 37044 28444
rect 37001 28407 37059 28413
rect 37001 28373 37013 28407
rect 37047 28404 37059 28407
rect 38010 28404 38016 28416
rect 37047 28376 38016 28404
rect 37047 28373 37059 28376
rect 37001 28367 37059 28373
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 38102 28364 38108 28416
rect 38160 28404 38166 28416
rect 38562 28404 38568 28416
rect 38160 28376 38568 28404
rect 38160 28364 38166 28376
rect 38562 28364 38568 28376
rect 38620 28404 38626 28416
rect 38841 28407 38899 28413
rect 38841 28404 38853 28407
rect 38620 28376 38853 28404
rect 38620 28364 38626 28376
rect 38841 28373 38853 28376
rect 38887 28373 38899 28407
rect 38841 28367 38899 28373
rect 1104 28314 48852 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 14246 28314
rect 14298 28262 14310 28314
rect 14362 28262 14374 28314
rect 14426 28262 14438 28314
rect 14490 28262 24246 28314
rect 24298 28262 24310 28314
rect 24362 28262 24374 28314
rect 24426 28262 24438 28314
rect 24490 28262 34246 28314
rect 34298 28262 34310 28314
rect 34362 28262 34374 28314
rect 34426 28262 34438 28314
rect 34490 28262 44246 28314
rect 44298 28262 44310 28314
rect 44362 28262 44374 28314
rect 44426 28262 44438 28314
rect 44490 28262 48852 28314
rect 1104 28240 48852 28262
rect 24118 28200 24124 28212
rect 22848 28172 24124 28200
rect 22002 27956 22008 28008
rect 22060 27996 22066 28008
rect 22848 28005 22876 28172
rect 24118 28160 24124 28172
rect 24176 28200 24182 28212
rect 24213 28203 24271 28209
rect 24213 28200 24225 28203
rect 24176 28172 24225 28200
rect 24176 28160 24182 28172
rect 24213 28169 24225 28172
rect 24259 28200 24271 28203
rect 24670 28200 24676 28212
rect 24259 28172 24676 28200
rect 24259 28169 24271 28172
rect 24213 28163 24271 28169
rect 24670 28160 24676 28172
rect 24728 28160 24734 28212
rect 24762 28160 24768 28212
rect 24820 28200 24826 28212
rect 32674 28200 32680 28212
rect 24820 28172 32680 28200
rect 24820 28160 24826 28172
rect 32674 28160 32680 28172
rect 32732 28160 32738 28212
rect 32769 28203 32827 28209
rect 32769 28169 32781 28203
rect 32815 28200 32827 28203
rect 33226 28200 33232 28212
rect 32815 28172 33232 28200
rect 32815 28169 32827 28172
rect 32769 28163 32827 28169
rect 33226 28160 33232 28172
rect 33284 28160 33290 28212
rect 23109 28135 23167 28141
rect 23109 28101 23121 28135
rect 23155 28132 23167 28135
rect 43438 28132 43444 28144
rect 23155 28104 43444 28132
rect 23155 28101 23167 28104
rect 23109 28095 23167 28101
rect 43438 28092 43444 28104
rect 43496 28092 43502 28144
rect 23753 28067 23811 28073
rect 23753 28064 23765 28067
rect 23124 28036 23765 28064
rect 23014 28005 23020 28008
rect 22557 27999 22615 28005
rect 22557 27996 22569 27999
rect 22060 27968 22569 27996
rect 22060 27956 22066 27968
rect 22557 27965 22569 27968
rect 22603 27965 22615 27999
rect 22557 27959 22615 27965
rect 22833 27999 22891 28005
rect 22833 27965 22845 27999
rect 22879 27965 22891 27999
rect 22833 27959 22891 27965
rect 22977 27999 23020 28005
rect 22977 27965 22989 27999
rect 22977 27959 23020 27965
rect 22572 27860 22600 27959
rect 23014 27956 23020 27959
rect 23072 27956 23078 28008
rect 22646 27888 22652 27940
rect 22704 27928 22710 27940
rect 22741 27931 22799 27937
rect 22741 27928 22753 27931
rect 22704 27900 22753 27928
rect 22704 27888 22710 27900
rect 22741 27897 22753 27900
rect 22787 27928 22799 27931
rect 23124 27928 23152 28036
rect 23753 28033 23765 28036
rect 23799 28064 23811 28067
rect 24578 28064 24584 28076
rect 23799 28036 24584 28064
rect 23799 28033 23811 28036
rect 23753 28027 23811 28033
rect 24578 28024 24584 28036
rect 24636 28024 24642 28076
rect 24854 28024 24860 28076
rect 24912 28064 24918 28076
rect 31570 28064 31576 28076
rect 24912 28036 31576 28064
rect 24912 28024 24918 28036
rect 31570 28024 31576 28036
rect 31628 28024 31634 28076
rect 31846 28064 31852 28076
rect 31807 28036 31852 28064
rect 31846 28024 31852 28036
rect 31904 28024 31910 28076
rect 33226 28064 33232 28076
rect 31956 28036 33232 28064
rect 31665 27999 31723 28005
rect 31665 27996 31677 27999
rect 22787 27900 23152 27928
rect 30944 27968 31677 27996
rect 22787 27897 22799 27900
rect 22741 27891 22799 27897
rect 30944 27872 30972 27968
rect 31665 27965 31677 27968
rect 31711 27965 31723 27999
rect 31665 27959 31723 27965
rect 31754 27956 31760 28008
rect 31812 27996 31818 28008
rect 31956 28005 31984 28036
rect 33226 28024 33232 28036
rect 33284 28024 33290 28076
rect 31941 27999 31999 28005
rect 31812 27968 31857 27996
rect 31812 27956 31818 27968
rect 31941 27965 31953 27999
rect 31987 27965 31999 27999
rect 31941 27959 31999 27965
rect 32125 27999 32183 28005
rect 32125 27965 32137 27999
rect 32171 27996 32183 27999
rect 32171 27968 33364 27996
rect 32171 27965 32183 27968
rect 32125 27959 32183 27965
rect 24762 27860 24768 27872
rect 22572 27832 24768 27860
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 30926 27860 30932 27872
rect 30887 27832 30932 27860
rect 30926 27820 30932 27832
rect 30984 27820 30990 27872
rect 31478 27860 31484 27872
rect 31439 27832 31484 27860
rect 31478 27820 31484 27832
rect 31536 27820 31542 27872
rect 31570 27820 31576 27872
rect 31628 27860 31634 27872
rect 31956 27860 31984 27959
rect 33336 27869 33364 27968
rect 31628 27832 31984 27860
rect 33321 27863 33379 27869
rect 31628 27820 31634 27832
rect 33321 27829 33333 27863
rect 33367 27860 33379 27863
rect 38930 27860 38936 27872
rect 33367 27832 38936 27860
rect 33367 27829 33379 27832
rect 33321 27823 33379 27829
rect 38930 27820 38936 27832
rect 38988 27820 38994 27872
rect 1104 27770 48852 27792
rect 1104 27718 9246 27770
rect 9298 27718 9310 27770
rect 9362 27718 9374 27770
rect 9426 27718 9438 27770
rect 9490 27718 19246 27770
rect 19298 27718 19310 27770
rect 19362 27718 19374 27770
rect 19426 27718 19438 27770
rect 19490 27718 29246 27770
rect 29298 27718 29310 27770
rect 29362 27718 29374 27770
rect 29426 27718 29438 27770
rect 29490 27718 39246 27770
rect 39298 27718 39310 27770
rect 39362 27718 39374 27770
rect 39426 27718 39438 27770
rect 39490 27718 48852 27770
rect 1104 27696 48852 27718
rect 10594 27616 10600 27668
rect 10652 27656 10658 27668
rect 30926 27656 30932 27668
rect 10652 27628 30932 27656
rect 10652 27616 10658 27628
rect 30926 27616 30932 27628
rect 30984 27616 30990 27668
rect 31846 27616 31852 27668
rect 31904 27656 31910 27668
rect 32766 27656 32772 27668
rect 31904 27628 32772 27656
rect 31904 27616 31910 27628
rect 32766 27616 32772 27628
rect 32824 27616 32830 27668
rect 1762 27588 1768 27600
rect 1723 27560 1768 27588
rect 1762 27548 1768 27560
rect 1820 27548 1826 27600
rect 4614 27548 4620 27600
rect 4672 27588 4678 27600
rect 5166 27588 5172 27600
rect 4672 27560 5172 27588
rect 4672 27548 4678 27560
rect 5166 27548 5172 27560
rect 5224 27548 5230 27600
rect 17218 27548 17224 27600
rect 17276 27588 17282 27600
rect 22465 27591 22523 27597
rect 22465 27588 22477 27591
rect 17276 27560 22477 27588
rect 17276 27548 17282 27560
rect 22465 27557 22477 27560
rect 22511 27588 22523 27591
rect 23014 27588 23020 27600
rect 22511 27560 23020 27588
rect 22511 27557 22523 27560
rect 22465 27551 22523 27557
rect 23014 27548 23020 27560
rect 23072 27548 23078 27600
rect 1949 27523 2007 27529
rect 1949 27489 1961 27523
rect 1995 27520 2007 27523
rect 2593 27523 2651 27529
rect 2593 27520 2605 27523
rect 1995 27492 2605 27520
rect 1995 27489 2007 27492
rect 1949 27483 2007 27489
rect 2593 27489 2605 27492
rect 2639 27520 2651 27523
rect 28258 27520 28264 27532
rect 2639 27492 28264 27520
rect 2639 27489 2651 27492
rect 2593 27483 2651 27489
rect 28258 27480 28264 27492
rect 28316 27480 28322 27532
rect 21910 27412 21916 27464
rect 21968 27452 21974 27464
rect 31113 27455 31171 27461
rect 31113 27452 31125 27455
rect 21968 27424 31125 27452
rect 21968 27412 21974 27424
rect 31113 27421 31125 27424
rect 31159 27452 31171 27455
rect 31754 27452 31760 27464
rect 31159 27424 31760 27452
rect 31159 27421 31171 27424
rect 31113 27415 31171 27421
rect 31754 27412 31760 27424
rect 31812 27452 31818 27464
rect 33042 27452 33048 27464
rect 31812 27424 33048 27452
rect 31812 27412 31818 27424
rect 33042 27412 33048 27424
rect 33100 27412 33106 27464
rect 1104 27226 48852 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 14246 27226
rect 14298 27174 14310 27226
rect 14362 27174 14374 27226
rect 14426 27174 14438 27226
rect 14490 27174 24246 27226
rect 24298 27174 24310 27226
rect 24362 27174 24374 27226
rect 24426 27174 24438 27226
rect 24490 27174 34246 27226
rect 34298 27174 34310 27226
rect 34362 27174 34374 27226
rect 34426 27174 34438 27226
rect 34490 27174 44246 27226
rect 44298 27174 44310 27226
rect 44362 27174 44374 27226
rect 44426 27174 44438 27226
rect 44490 27174 48852 27226
rect 1104 27152 48852 27174
rect 15930 27072 15936 27124
rect 15988 27112 15994 27124
rect 33134 27112 33140 27124
rect 15988 27084 33140 27112
rect 15988 27072 15994 27084
rect 33134 27072 33140 27084
rect 33192 27072 33198 27124
rect 34425 27115 34483 27121
rect 34425 27081 34437 27115
rect 34471 27112 34483 27115
rect 37274 27112 37280 27124
rect 34471 27084 37280 27112
rect 34471 27081 34483 27084
rect 34425 27075 34483 27081
rect 37274 27072 37280 27084
rect 37332 27072 37338 27124
rect 33042 27004 33048 27056
rect 33100 27044 33106 27056
rect 41598 27044 41604 27056
rect 33100 27016 41604 27044
rect 33100 27004 33106 27016
rect 41598 27004 41604 27016
rect 41656 27004 41662 27056
rect 17954 26936 17960 26988
rect 18012 26976 18018 26988
rect 25774 26976 25780 26988
rect 18012 26948 25780 26976
rect 18012 26936 18018 26948
rect 25774 26936 25780 26948
rect 25832 26976 25838 26988
rect 25832 26948 31754 26976
rect 25832 26936 25838 26948
rect 2958 26868 2964 26920
rect 3016 26908 3022 26920
rect 4065 26911 4123 26917
rect 4065 26908 4077 26911
rect 3016 26880 4077 26908
rect 3016 26868 3022 26880
rect 4065 26877 4077 26880
rect 4111 26908 4123 26911
rect 6730 26908 6736 26920
rect 4111 26880 6736 26908
rect 4111 26877 4123 26880
rect 4065 26871 4123 26877
rect 6730 26868 6736 26880
rect 6788 26908 6794 26920
rect 17218 26908 17224 26920
rect 6788 26880 17224 26908
rect 6788 26868 6794 26880
rect 17218 26868 17224 26880
rect 17276 26868 17282 26920
rect 19978 26868 19984 26920
rect 20036 26908 20042 26920
rect 30006 26908 30012 26920
rect 20036 26880 30012 26908
rect 20036 26868 20042 26880
rect 30006 26868 30012 26880
rect 30064 26868 30070 26920
rect 31726 26908 31754 26948
rect 34333 26911 34391 26917
rect 34333 26908 34345 26911
rect 31726 26880 34345 26908
rect 34333 26877 34345 26880
rect 34379 26908 34391 26911
rect 34379 26880 35112 26908
rect 34379 26877 34391 26880
rect 34333 26871 34391 26877
rect 30285 26843 30343 26849
rect 30285 26809 30297 26843
rect 30331 26809 30343 26843
rect 31510 26812 32720 26840
rect 30285 26803 30343 26809
rect 13630 26732 13636 26784
rect 13688 26772 13694 26784
rect 29457 26775 29515 26781
rect 29457 26772 29469 26775
rect 13688 26744 29469 26772
rect 13688 26732 13694 26744
rect 29457 26741 29469 26744
rect 29503 26772 29515 26775
rect 30300 26772 30328 26803
rect 32692 26784 32720 26812
rect 29503 26744 30328 26772
rect 29503 26741 29515 26744
rect 29457 26735 29515 26741
rect 31754 26732 31760 26784
rect 31812 26772 31818 26784
rect 32674 26772 32680 26784
rect 31812 26744 31857 26772
rect 32635 26744 32680 26772
rect 31812 26732 31818 26744
rect 32674 26732 32680 26744
rect 32732 26732 32738 26784
rect 35084 26781 35112 26880
rect 35069 26775 35127 26781
rect 35069 26741 35081 26775
rect 35115 26772 35127 26775
rect 37734 26772 37740 26784
rect 35115 26744 37740 26772
rect 35115 26741 35127 26744
rect 35069 26735 35127 26741
rect 37734 26732 37740 26744
rect 37792 26732 37798 26784
rect 1104 26682 48852 26704
rect 1104 26630 9246 26682
rect 9298 26630 9310 26682
rect 9362 26630 9374 26682
rect 9426 26630 9438 26682
rect 9490 26630 19246 26682
rect 19298 26630 19310 26682
rect 19362 26630 19374 26682
rect 19426 26630 19438 26682
rect 19490 26630 29246 26682
rect 29298 26630 29310 26682
rect 29362 26630 29374 26682
rect 29426 26630 29438 26682
rect 29490 26630 39246 26682
rect 39298 26630 39310 26682
rect 39362 26630 39374 26682
rect 39426 26630 39438 26682
rect 39490 26630 48852 26682
rect 1104 26608 48852 26630
rect 30006 26528 30012 26580
rect 30064 26568 30070 26580
rect 32217 26571 32275 26577
rect 32217 26568 32229 26571
rect 30064 26540 32229 26568
rect 30064 26528 30070 26540
rect 32217 26537 32229 26540
rect 32263 26568 32275 26571
rect 32398 26568 32404 26580
rect 32263 26540 32404 26568
rect 32263 26537 32275 26540
rect 32217 26531 32275 26537
rect 32398 26528 32404 26540
rect 32456 26528 32462 26580
rect 2958 26441 2964 26444
rect 2956 26432 2964 26441
rect 2919 26404 2964 26432
rect 2956 26395 2964 26404
rect 2958 26392 2964 26395
rect 3016 26392 3022 26444
rect 3053 26435 3111 26441
rect 3053 26401 3065 26435
rect 3099 26401 3111 26435
rect 3053 26395 3111 26401
rect 3145 26435 3203 26441
rect 3145 26401 3157 26435
rect 3191 26401 3203 26435
rect 3145 26395 3203 26401
rect 3329 26435 3387 26441
rect 3329 26401 3341 26435
rect 3375 26432 3387 26435
rect 4614 26432 4620 26444
rect 3375 26404 4620 26432
rect 3375 26401 3387 26404
rect 3329 26395 3387 26401
rect 2777 26299 2835 26305
rect 2777 26265 2789 26299
rect 2823 26296 2835 26299
rect 2866 26296 2872 26308
rect 2823 26268 2872 26296
rect 2823 26265 2835 26268
rect 2777 26259 2835 26265
rect 2866 26256 2872 26268
rect 2924 26256 2930 26308
rect 3068 26296 3096 26395
rect 3160 26364 3188 26395
rect 4614 26392 4620 26404
rect 4672 26392 4678 26444
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3160 26336 3985 26364
rect 3973 26333 3985 26336
rect 4019 26364 4031 26367
rect 17954 26364 17960 26376
rect 4019 26336 17960 26364
rect 4019 26333 4031 26336
rect 3973 26327 4031 26333
rect 17954 26324 17960 26336
rect 18012 26324 18018 26376
rect 4525 26299 4583 26305
rect 4525 26296 4537 26299
rect 3068 26268 4537 26296
rect 4525 26265 4537 26268
rect 4571 26296 4583 26299
rect 15930 26296 15936 26308
rect 4571 26268 15936 26296
rect 4571 26265 4583 26268
rect 4525 26259 4583 26265
rect 15930 26256 15936 26268
rect 15988 26256 15994 26308
rect 1104 26138 48852 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 14246 26138
rect 14298 26086 14310 26138
rect 14362 26086 14374 26138
rect 14426 26086 14438 26138
rect 14490 26086 24246 26138
rect 24298 26086 24310 26138
rect 24362 26086 24374 26138
rect 24426 26086 24438 26138
rect 24490 26086 34246 26138
rect 34298 26086 34310 26138
rect 34362 26086 34374 26138
rect 34426 26086 34438 26138
rect 34490 26086 44246 26138
rect 44298 26086 44310 26138
rect 44362 26086 44374 26138
rect 44426 26086 44438 26138
rect 44490 26086 48852 26138
rect 1104 26064 48852 26086
rect 3881 25687 3939 25693
rect 3881 25653 3893 25687
rect 3927 25684 3939 25687
rect 4614 25684 4620 25696
rect 3927 25656 4620 25684
rect 3927 25653 3939 25656
rect 3881 25647 3939 25653
rect 4614 25644 4620 25656
rect 4672 25684 4678 25696
rect 18138 25684 18144 25696
rect 4672 25656 18144 25684
rect 4672 25644 4678 25656
rect 18138 25644 18144 25656
rect 18196 25644 18202 25696
rect 42058 25644 42064 25696
rect 42116 25684 42122 25696
rect 45922 25684 45928 25696
rect 42116 25656 45928 25684
rect 42116 25644 42122 25656
rect 45922 25644 45928 25656
rect 45980 25644 45986 25696
rect 1104 25594 48852 25616
rect 1104 25542 9246 25594
rect 9298 25542 9310 25594
rect 9362 25542 9374 25594
rect 9426 25542 9438 25594
rect 9490 25542 19246 25594
rect 19298 25542 19310 25594
rect 19362 25542 19374 25594
rect 19426 25542 19438 25594
rect 19490 25542 29246 25594
rect 29298 25542 29310 25594
rect 29362 25542 29374 25594
rect 29426 25542 29438 25594
rect 29490 25542 39246 25594
rect 39298 25542 39310 25594
rect 39362 25542 39374 25594
rect 39426 25542 39438 25594
rect 39490 25542 48852 25594
rect 1104 25520 48852 25542
rect 45646 25480 45652 25492
rect 45526 25452 45652 25480
rect 37366 25372 37372 25424
rect 37424 25412 37430 25424
rect 38010 25412 38016 25424
rect 37424 25384 38016 25412
rect 37424 25372 37430 25384
rect 38010 25372 38016 25384
rect 38068 25412 38074 25424
rect 45526 25412 45554 25452
rect 45646 25440 45652 25452
rect 45704 25480 45710 25492
rect 46750 25480 46756 25492
rect 45704 25452 46756 25480
rect 45704 25440 45710 25452
rect 46750 25440 46756 25452
rect 46808 25440 46814 25492
rect 38068 25384 45554 25412
rect 38068 25372 38074 25384
rect 45922 25372 45928 25424
rect 45980 25412 45986 25424
rect 46477 25415 46535 25421
rect 46477 25412 46489 25415
rect 45980 25384 46489 25412
rect 45980 25372 45986 25384
rect 46477 25381 46489 25384
rect 46523 25381 46535 25415
rect 46477 25375 46535 25381
rect 45186 25304 45192 25356
rect 45244 25344 45250 25356
rect 46385 25347 46443 25353
rect 46385 25344 46397 25347
rect 45244 25316 46397 25344
rect 45244 25304 45250 25316
rect 46385 25313 46397 25316
rect 46431 25313 46443 25347
rect 46566 25344 46572 25356
rect 46527 25316 46572 25344
rect 46385 25307 46443 25313
rect 46566 25304 46572 25316
rect 46624 25304 46630 25356
rect 46750 25344 46756 25356
rect 46711 25316 46756 25344
rect 46750 25304 46756 25316
rect 46808 25304 46814 25356
rect 47489 25347 47547 25353
rect 47489 25313 47501 25347
rect 47535 25344 47547 25347
rect 48130 25344 48136 25356
rect 47535 25316 48136 25344
rect 47535 25313 47547 25316
rect 47489 25307 47547 25313
rect 48130 25304 48136 25316
rect 48188 25304 48194 25356
rect 45186 25140 45192 25152
rect 45147 25112 45192 25140
rect 45186 25100 45192 25112
rect 45244 25100 45250 25152
rect 46198 25140 46204 25152
rect 46159 25112 46204 25140
rect 46198 25100 46204 25112
rect 46256 25100 46262 25152
rect 47946 25140 47952 25152
rect 47907 25112 47952 25140
rect 47946 25100 47952 25112
rect 48004 25100 48010 25152
rect 1104 25050 48852 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 14246 25050
rect 14298 24998 14310 25050
rect 14362 24998 14374 25050
rect 14426 24998 14438 25050
rect 14490 24998 24246 25050
rect 24298 24998 24310 25050
rect 24362 24998 24374 25050
rect 24426 24998 24438 25050
rect 24490 24998 34246 25050
rect 34298 24998 34310 25050
rect 34362 24998 34374 25050
rect 34426 24998 34438 25050
rect 34490 24998 44246 25050
rect 44298 24998 44310 25050
rect 44362 24998 44374 25050
rect 44426 24998 44438 25050
rect 44490 24998 48852 25050
rect 1104 24976 48852 24998
rect 46109 24939 46167 24945
rect 46109 24936 46121 24939
rect 45526 24908 46121 24936
rect 39758 24828 39764 24880
rect 39816 24828 39822 24880
rect 42058 24828 42064 24880
rect 42116 24868 42122 24880
rect 42610 24868 42616 24880
rect 42116 24840 42616 24868
rect 42116 24828 42122 24840
rect 42610 24828 42616 24840
rect 42668 24828 42674 24880
rect 38930 24760 38936 24812
rect 38988 24800 38994 24812
rect 39776 24800 39804 24828
rect 45526 24800 45554 24908
rect 46109 24905 46121 24908
rect 46155 24936 46167 24939
rect 46566 24936 46572 24948
rect 46155 24908 46572 24936
rect 46155 24905 46167 24908
rect 46109 24899 46167 24905
rect 46566 24896 46572 24908
rect 46624 24896 46630 24948
rect 38988 24772 45554 24800
rect 38988 24760 38994 24772
rect 39666 24692 39672 24744
rect 39724 24732 39730 24744
rect 39761 24735 39819 24741
rect 39761 24732 39773 24735
rect 39724 24704 39773 24732
rect 39724 24692 39730 24704
rect 39761 24701 39773 24704
rect 39807 24732 39819 24735
rect 39850 24732 39856 24744
rect 39807 24704 39856 24732
rect 39807 24701 39819 24704
rect 39761 24695 39819 24701
rect 39850 24692 39856 24704
rect 39908 24732 39914 24744
rect 40589 24735 40647 24741
rect 40589 24732 40601 24735
rect 39908 24704 40601 24732
rect 39908 24692 39914 24704
rect 40589 24701 40601 24704
rect 40635 24701 40647 24735
rect 40589 24695 40647 24701
rect 45557 24735 45615 24741
rect 45557 24701 45569 24735
rect 45603 24732 45615 24735
rect 45646 24732 45652 24744
rect 45603 24704 45652 24732
rect 45603 24701 45615 24704
rect 45557 24695 45615 24701
rect 45646 24692 45652 24704
rect 45704 24692 45710 24744
rect 28537 24667 28595 24673
rect 28537 24633 28549 24667
rect 28583 24633 28595 24667
rect 28537 24627 28595 24633
rect 13722 24556 13728 24608
rect 13780 24596 13786 24608
rect 27985 24599 28043 24605
rect 27985 24596 27997 24599
rect 13780 24568 27997 24596
rect 13780 24556 13786 24568
rect 27985 24565 27997 24568
rect 28031 24596 28043 24599
rect 28552 24596 28580 24627
rect 39482 24624 39488 24676
rect 39540 24664 39546 24676
rect 40221 24667 40279 24673
rect 40221 24664 40233 24667
rect 39540 24636 40233 24664
rect 39540 24624 39546 24636
rect 40221 24633 40233 24636
rect 40267 24633 40279 24667
rect 40221 24627 40279 24633
rect 28031 24568 28580 24596
rect 28031 24565 28043 24568
rect 27985 24559 28043 24565
rect 29730 24556 29736 24608
rect 29788 24596 29794 24608
rect 29825 24599 29883 24605
rect 29825 24596 29837 24599
rect 29788 24568 29837 24596
rect 29788 24556 29794 24568
rect 29825 24565 29837 24568
rect 29871 24565 29883 24599
rect 29825 24559 29883 24565
rect 1104 24506 48852 24528
rect 1104 24454 9246 24506
rect 9298 24454 9310 24506
rect 9362 24454 9374 24506
rect 9426 24454 9438 24506
rect 9490 24454 19246 24506
rect 19298 24454 19310 24506
rect 19362 24454 19374 24506
rect 19426 24454 19438 24506
rect 19490 24454 29246 24506
rect 29298 24454 29310 24506
rect 29362 24454 29374 24506
rect 29426 24454 29438 24506
rect 29490 24454 39246 24506
rect 39298 24454 39310 24506
rect 39362 24454 39374 24506
rect 39426 24454 39438 24506
rect 39490 24454 48852 24506
rect 1104 24432 48852 24454
rect 19705 24395 19763 24401
rect 19705 24361 19717 24395
rect 19751 24392 19763 24395
rect 19978 24392 19984 24404
rect 19751 24364 19984 24392
rect 19751 24361 19763 24364
rect 19705 24355 19763 24361
rect 18877 24259 18935 24265
rect 18877 24225 18889 24259
rect 18923 24256 18935 24259
rect 19720 24256 19748 24355
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 36081 24327 36139 24333
rect 36081 24293 36093 24327
rect 36127 24324 36139 24327
rect 37550 24324 37556 24336
rect 36127 24296 37556 24324
rect 36127 24293 36139 24296
rect 36081 24287 36139 24293
rect 37550 24284 37556 24296
rect 37608 24284 37614 24336
rect 35710 24256 35716 24268
rect 18923 24228 19748 24256
rect 35671 24228 35716 24256
rect 18923 24225 18935 24228
rect 18877 24219 18935 24225
rect 35710 24216 35716 24228
rect 35768 24216 35774 24268
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 23474 24188 23480 24200
rect 18647 24160 23480 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 23474 24148 23480 24160
rect 23532 24148 23538 24200
rect 17310 24012 17316 24064
rect 17368 24052 17374 24064
rect 17494 24052 17500 24064
rect 17368 24024 17500 24052
rect 17368 24012 17374 24024
rect 17494 24012 17500 24024
rect 17552 24012 17558 24064
rect 1104 23962 48852 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 14246 23962
rect 14298 23910 14310 23962
rect 14362 23910 14374 23962
rect 14426 23910 14438 23962
rect 14490 23910 24246 23962
rect 24298 23910 24310 23962
rect 24362 23910 24374 23962
rect 24426 23910 24438 23962
rect 24490 23910 34246 23962
rect 34298 23910 34310 23962
rect 34362 23910 34374 23962
rect 34426 23910 34438 23962
rect 34490 23910 44246 23962
rect 44298 23910 44310 23962
rect 44362 23910 44374 23962
rect 44426 23910 44438 23962
rect 44490 23910 48852 23962
rect 1104 23888 48852 23910
rect 17494 23808 17500 23860
rect 17552 23848 17558 23860
rect 43530 23848 43536 23860
rect 17552 23820 43536 23848
rect 17552 23808 17558 23820
rect 43530 23808 43536 23820
rect 43588 23808 43594 23860
rect 31754 23740 31760 23792
rect 31812 23780 31818 23792
rect 35529 23783 35587 23789
rect 35529 23780 35541 23783
rect 31812 23752 35541 23780
rect 31812 23740 31818 23752
rect 35529 23749 35541 23752
rect 35575 23780 35587 23783
rect 35710 23780 35716 23792
rect 35575 23752 35716 23780
rect 35575 23749 35587 23752
rect 35529 23743 35587 23749
rect 35710 23740 35716 23752
rect 35768 23740 35774 23792
rect 1104 23418 48852 23440
rect 1104 23366 9246 23418
rect 9298 23366 9310 23418
rect 9362 23366 9374 23418
rect 9426 23366 9438 23418
rect 9490 23366 19246 23418
rect 19298 23366 19310 23418
rect 19362 23366 19374 23418
rect 19426 23366 19438 23418
rect 19490 23366 29246 23418
rect 29298 23366 29310 23418
rect 29362 23366 29374 23418
rect 29426 23366 29438 23418
rect 29490 23366 39246 23418
rect 39298 23366 39310 23418
rect 39362 23366 39374 23418
rect 39426 23366 39438 23418
rect 39490 23366 48852 23418
rect 1104 23344 48852 23366
rect 25682 23264 25688 23316
rect 25740 23304 25746 23316
rect 25777 23307 25835 23313
rect 25777 23304 25789 23307
rect 25740 23276 25789 23304
rect 25740 23264 25746 23276
rect 25777 23273 25789 23276
rect 25823 23273 25835 23307
rect 25777 23267 25835 23273
rect 24670 23128 24676 23180
rect 24728 23168 24734 23180
rect 25869 23171 25927 23177
rect 25869 23168 25881 23171
rect 24728 23140 25881 23168
rect 24728 23128 24734 23140
rect 25869 23137 25881 23140
rect 25915 23168 25927 23171
rect 25915 23140 26234 23168
rect 25915 23137 25927 23140
rect 25869 23131 25927 23137
rect 26206 22964 26234 23140
rect 26421 22967 26479 22973
rect 26421 22964 26433 22967
rect 26206 22936 26433 22964
rect 26421 22933 26433 22936
rect 26467 22964 26479 22967
rect 39574 22964 39580 22976
rect 26467 22936 39580 22964
rect 26467 22933 26479 22936
rect 26421 22927 26479 22933
rect 39574 22924 39580 22936
rect 39632 22924 39638 22976
rect 1104 22874 48852 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 14246 22874
rect 14298 22822 14310 22874
rect 14362 22822 14374 22874
rect 14426 22822 14438 22874
rect 14490 22822 24246 22874
rect 24298 22822 24310 22874
rect 24362 22822 24374 22874
rect 24426 22822 24438 22874
rect 24490 22822 34246 22874
rect 34298 22822 34310 22874
rect 34362 22822 34374 22874
rect 34426 22822 34438 22874
rect 34490 22822 44246 22874
rect 44298 22822 44310 22874
rect 44362 22822 44374 22874
rect 44426 22822 44438 22874
rect 44490 22822 48852 22874
rect 1104 22800 48852 22822
rect 1762 22488 1768 22500
rect 1723 22460 1768 22488
rect 1762 22448 1768 22460
rect 1820 22448 1826 22500
rect 1949 22491 2007 22497
rect 1949 22457 1961 22491
rect 1995 22457 2007 22491
rect 1949 22451 2007 22457
rect 1964 22420 1992 22451
rect 2593 22423 2651 22429
rect 2593 22420 2605 22423
rect 1964 22392 2605 22420
rect 2593 22389 2605 22392
rect 2639 22420 2651 22423
rect 11698 22420 11704 22432
rect 2639 22392 11704 22420
rect 2639 22389 2651 22392
rect 2593 22383 2651 22389
rect 11698 22380 11704 22392
rect 11756 22380 11762 22432
rect 1104 22330 48852 22352
rect 1104 22278 9246 22330
rect 9298 22278 9310 22330
rect 9362 22278 9374 22330
rect 9426 22278 9438 22330
rect 9490 22278 19246 22330
rect 19298 22278 19310 22330
rect 19362 22278 19374 22330
rect 19426 22278 19438 22330
rect 19490 22278 29246 22330
rect 29298 22278 29310 22330
rect 29362 22278 29374 22330
rect 29426 22278 29438 22330
rect 29490 22278 39246 22330
rect 39298 22278 39310 22330
rect 39362 22278 39374 22330
rect 39426 22278 39438 22330
rect 39490 22278 48852 22330
rect 1104 22256 48852 22278
rect 11698 22108 11704 22160
rect 11756 22148 11762 22160
rect 12158 22148 12164 22160
rect 11756 22120 12164 22148
rect 11756 22108 11762 22120
rect 12158 22108 12164 22120
rect 12216 22108 12222 22160
rect 26513 22083 26571 22089
rect 26513 22080 26525 22083
rect 26206 22052 26525 22080
rect 18414 21836 18420 21888
rect 18472 21876 18478 21888
rect 26206 21876 26234 22052
rect 26513 22049 26525 22052
rect 26559 22080 26571 22083
rect 27229 22083 27287 22089
rect 27229 22080 27241 22083
rect 26559 22052 27241 22080
rect 26559 22049 26571 22052
rect 26513 22043 26571 22049
rect 27229 22049 27241 22052
rect 27275 22049 27287 22083
rect 27229 22043 27287 22049
rect 26973 22015 27031 22021
rect 26973 21981 26985 22015
rect 27019 21981 27031 22015
rect 26973 21975 27031 21981
rect 18472 21848 26234 21876
rect 26988 21876 27016 21975
rect 28258 21904 28264 21956
rect 28316 21944 28322 21956
rect 28353 21947 28411 21953
rect 28353 21944 28365 21947
rect 28316 21916 28365 21944
rect 28316 21904 28322 21916
rect 28353 21913 28365 21916
rect 28399 21913 28411 21947
rect 28353 21907 28411 21913
rect 28997 21879 29055 21885
rect 28997 21876 29009 21879
rect 26988 21848 29009 21876
rect 18472 21836 18478 21848
rect 28997 21845 29009 21848
rect 29043 21876 29055 21879
rect 29546 21876 29552 21888
rect 29043 21848 29552 21876
rect 29043 21845 29055 21848
rect 28997 21839 29055 21845
rect 29546 21836 29552 21848
rect 29604 21836 29610 21888
rect 1104 21786 48852 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 14246 21786
rect 14298 21734 14310 21786
rect 14362 21734 14374 21786
rect 14426 21734 14438 21786
rect 14490 21734 24246 21786
rect 24298 21734 24310 21786
rect 24362 21734 24374 21786
rect 24426 21734 24438 21786
rect 24490 21734 34246 21786
rect 34298 21734 34310 21786
rect 34362 21734 34374 21786
rect 34426 21734 34438 21786
rect 34490 21734 44246 21786
rect 44298 21734 44310 21786
rect 44362 21734 44374 21786
rect 44426 21734 44438 21786
rect 44490 21734 48852 21786
rect 1104 21712 48852 21734
rect 1104 21242 48852 21264
rect 1104 21190 9246 21242
rect 9298 21190 9310 21242
rect 9362 21190 9374 21242
rect 9426 21190 9438 21242
rect 9490 21190 19246 21242
rect 19298 21190 19310 21242
rect 19362 21190 19374 21242
rect 19426 21190 19438 21242
rect 19490 21190 29246 21242
rect 29298 21190 29310 21242
rect 29362 21190 29374 21242
rect 29426 21190 29438 21242
rect 29490 21190 39246 21242
rect 39298 21190 39310 21242
rect 39362 21190 39374 21242
rect 39426 21190 39438 21242
rect 39490 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 14246 20698
rect 14298 20646 14310 20698
rect 14362 20646 14374 20698
rect 14426 20646 14438 20698
rect 14490 20646 24246 20698
rect 24298 20646 24310 20698
rect 24362 20646 24374 20698
rect 24426 20646 24438 20698
rect 24490 20646 34246 20698
rect 34298 20646 34310 20698
rect 34362 20646 34374 20698
rect 34426 20646 34438 20698
rect 34490 20646 44246 20698
rect 44298 20646 44310 20698
rect 44362 20646 44374 20698
rect 44426 20646 44438 20698
rect 44490 20646 48852 20698
rect 1104 20624 48852 20646
rect 27246 20204 27252 20256
rect 27304 20244 27310 20256
rect 27617 20247 27675 20253
rect 27617 20244 27629 20247
rect 27304 20216 27629 20244
rect 27304 20204 27310 20216
rect 27617 20213 27629 20216
rect 27663 20244 27675 20247
rect 44542 20244 44548 20256
rect 27663 20216 44548 20244
rect 27663 20213 27675 20216
rect 27617 20207 27675 20213
rect 44542 20204 44548 20216
rect 44600 20204 44606 20256
rect 1104 20154 48852 20176
rect 1104 20102 9246 20154
rect 9298 20102 9310 20154
rect 9362 20102 9374 20154
rect 9426 20102 9438 20154
rect 9490 20102 19246 20154
rect 19298 20102 19310 20154
rect 19362 20102 19374 20154
rect 19426 20102 19438 20154
rect 19490 20102 29246 20154
rect 29298 20102 29310 20154
rect 29362 20102 29374 20154
rect 29426 20102 29438 20154
rect 29490 20102 39246 20154
rect 39298 20102 39310 20154
rect 39362 20102 39374 20154
rect 39426 20102 39438 20154
rect 39490 20102 48852 20154
rect 1104 20080 48852 20102
rect 23474 20000 23480 20052
rect 23532 20040 23538 20052
rect 26881 20043 26939 20049
rect 26881 20040 26893 20043
rect 23532 20012 26893 20040
rect 23532 20000 23538 20012
rect 26881 20009 26893 20012
rect 26927 20009 26939 20043
rect 26881 20003 26939 20009
rect 27246 19972 27252 19984
rect 27207 19944 27252 19972
rect 27246 19932 27252 19944
rect 27304 19932 27310 19984
rect 30834 19932 30840 19984
rect 30892 19972 30898 19984
rect 30929 19975 30987 19981
rect 30929 19972 30941 19975
rect 30892 19944 30941 19972
rect 30892 19932 30898 19944
rect 30929 19941 30941 19944
rect 30975 19972 30987 19975
rect 31570 19972 31576 19984
rect 30975 19944 31576 19972
rect 30975 19941 30987 19944
rect 30929 19935 30987 19941
rect 31570 19932 31576 19944
rect 31628 19972 31634 19984
rect 32493 19975 32551 19981
rect 32493 19972 32505 19975
rect 31628 19944 32505 19972
rect 31628 19932 31634 19944
rect 32493 19941 32505 19944
rect 32539 19941 32551 19975
rect 32493 19935 32551 19941
rect 27065 19907 27123 19913
rect 27065 19873 27077 19907
rect 27111 19904 27123 19907
rect 27522 19904 27528 19916
rect 27111 19876 27528 19904
rect 27111 19873 27123 19876
rect 27065 19867 27123 19873
rect 27522 19864 27528 19876
rect 27580 19864 27586 19916
rect 29730 19904 29736 19916
rect 29691 19876 29736 19904
rect 29730 19864 29736 19876
rect 29788 19864 29794 19916
rect 31113 19907 31171 19913
rect 31113 19873 31125 19907
rect 31159 19873 31171 19907
rect 31113 19867 31171 19873
rect 31481 19907 31539 19913
rect 31481 19873 31493 19907
rect 31527 19904 31539 19907
rect 33778 19904 33784 19916
rect 31527 19876 33784 19904
rect 31527 19873 31539 19876
rect 31481 19867 31539 19873
rect 18138 19796 18144 19848
rect 18196 19836 18202 19848
rect 31128 19836 31156 19867
rect 33778 19864 33784 19876
rect 33836 19864 33842 19916
rect 31754 19836 31760 19848
rect 18196 19808 31760 19836
rect 18196 19796 18202 19808
rect 31754 19796 31760 19808
rect 31812 19836 31818 19848
rect 31941 19839 31999 19845
rect 31941 19836 31953 19839
rect 31812 19808 31953 19836
rect 31812 19796 31818 19808
rect 31941 19805 31953 19808
rect 31987 19805 31999 19839
rect 31941 19799 31999 19805
rect 27522 19660 27528 19712
rect 27580 19700 27586 19712
rect 27893 19703 27951 19709
rect 27893 19700 27905 19703
rect 27580 19672 27905 19700
rect 27580 19660 27586 19672
rect 27893 19669 27905 19672
rect 27939 19669 27951 19703
rect 29546 19700 29552 19712
rect 29507 19672 29552 19700
rect 27893 19663 27951 19669
rect 29546 19660 29552 19672
rect 29604 19660 29610 19712
rect 1104 19610 48852 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 14246 19610
rect 14298 19558 14310 19610
rect 14362 19558 14374 19610
rect 14426 19558 14438 19610
rect 14490 19558 24246 19610
rect 24298 19558 24310 19610
rect 24362 19558 24374 19610
rect 24426 19558 24438 19610
rect 24490 19558 34246 19610
rect 34298 19558 34310 19610
rect 34362 19558 34374 19610
rect 34426 19558 34438 19610
rect 34490 19558 44246 19610
rect 44298 19558 44310 19610
rect 44362 19558 44374 19610
rect 44426 19558 44438 19610
rect 44490 19558 48852 19610
rect 1104 19536 48852 19558
rect 5077 19363 5135 19369
rect 5077 19360 5089 19363
rect 3804 19332 5089 19360
rect 3418 19292 3424 19304
rect 3379 19264 3424 19292
rect 3418 19252 3424 19264
rect 3476 19252 3482 19304
rect 3804 19301 3832 19332
rect 5077 19329 5089 19332
rect 5123 19360 5135 19363
rect 5123 19332 5672 19360
rect 5123 19329 5135 19332
rect 5077 19323 5135 19329
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19261 3847 19295
rect 4525 19295 4583 19301
rect 4525 19292 4537 19295
rect 3789 19255 3847 19261
rect 3896 19264 4537 19292
rect 2961 19227 3019 19233
rect 2961 19193 2973 19227
rect 3007 19224 3019 19227
rect 3602 19224 3608 19236
rect 3007 19196 3608 19224
rect 3007 19193 3019 19196
rect 2961 19187 3019 19193
rect 3602 19184 3608 19196
rect 3660 19184 3666 19236
rect 3697 19227 3755 19233
rect 3697 19193 3709 19227
rect 3743 19224 3755 19227
rect 3896 19224 3924 19264
rect 4525 19261 4537 19264
rect 4571 19292 4583 19295
rect 5644 19292 5672 19332
rect 13078 19292 13084 19304
rect 4571 19264 5580 19292
rect 5644 19264 13084 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 5552 19224 5580 19264
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 13354 19224 13360 19236
rect 3743 19196 3924 19224
rect 3988 19196 5488 19224
rect 5552 19196 13360 19224
rect 3743 19193 3755 19196
rect 3697 19187 3755 19193
rect 3988 19165 4016 19196
rect 3973 19159 4031 19165
rect 3973 19125 3985 19159
rect 4019 19125 4031 19159
rect 5460 19156 5488 19196
rect 13354 19184 13360 19196
rect 13412 19224 13418 19236
rect 17862 19224 17868 19236
rect 13412 19196 17868 19224
rect 13412 19184 13418 19196
rect 17862 19184 17868 19196
rect 17920 19184 17926 19236
rect 15102 19156 15108 19168
rect 5460 19128 15108 19156
rect 3973 19119 4031 19125
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 1104 19066 18952 19088
rect 1104 19014 9246 19066
rect 9298 19014 9310 19066
rect 9362 19014 9374 19066
rect 9426 19014 9438 19066
rect 9490 19014 18952 19066
rect 1104 18992 18952 19014
rect 37628 19066 48852 19088
rect 37628 19014 39246 19066
rect 39298 19014 39310 19066
rect 39362 19014 39374 19066
rect 39426 19014 39438 19066
rect 39490 19014 48852 19066
rect 37628 18992 48852 19014
rect 3418 18572 3424 18624
rect 3476 18612 3482 18624
rect 4525 18615 4583 18621
rect 4525 18612 4537 18615
rect 3476 18584 4537 18612
rect 3476 18572 3482 18584
rect 4525 18581 4537 18584
rect 4571 18612 4583 18615
rect 27522 18612 27528 18624
rect 4571 18584 27528 18612
rect 4571 18581 4583 18584
rect 4525 18575 4583 18581
rect 27522 18572 27528 18584
rect 27580 18612 27586 18624
rect 37642 18612 37648 18624
rect 27580 18584 37648 18612
rect 27580 18572 27586 18584
rect 37642 18572 37648 18584
rect 37700 18572 37706 18624
rect 1104 18522 18952 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 14246 18522
rect 14298 18470 14310 18522
rect 14362 18470 14374 18522
rect 14426 18470 14438 18522
rect 14490 18470 18952 18522
rect 1104 18448 18952 18470
rect 37628 18522 48852 18544
rect 37628 18470 44246 18522
rect 44298 18470 44310 18522
rect 44362 18470 44374 18522
rect 44426 18470 44438 18522
rect 44490 18470 48852 18522
rect 37628 18448 48852 18470
rect 14182 18068 14188 18080
rect 14143 18040 14188 18068
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 1104 17978 18952 18000
rect 1104 17926 9246 17978
rect 9298 17926 9310 17978
rect 9362 17926 9374 17978
rect 9426 17926 9438 17978
rect 9490 17926 18952 17978
rect 1104 17904 18952 17926
rect 37628 17978 48852 18000
rect 37628 17926 39246 17978
rect 39298 17926 39310 17978
rect 39362 17926 39374 17978
rect 39426 17926 39438 17978
rect 39490 17926 48852 17978
rect 37628 17904 48852 17926
rect 12250 17864 12256 17876
rect 12211 17836 12256 17864
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 15102 17796 15108 17808
rect 15063 17768 15108 17796
rect 15102 17756 15108 17768
rect 15160 17756 15166 17808
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 1995 17700 2636 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 2608 17536 2636 17700
rect 13538 17660 13544 17672
rect 13499 17632 13544 17660
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 13817 17663 13875 17669
rect 13817 17629 13829 17663
rect 13863 17660 13875 17663
rect 14182 17660 14188 17672
rect 13863 17632 14188 17660
rect 13863 17629 13875 17632
rect 13817 17623 13875 17629
rect 14182 17620 14188 17632
rect 14240 17660 14246 17672
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 14240 17632 14841 17660
rect 14240 17620 14246 17632
rect 14829 17629 14841 17632
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 1854 17524 1860 17536
rect 1815 17496 1860 17524
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 2590 17524 2596 17536
rect 2551 17496 2596 17524
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 14844 17524 14872 17623
rect 16224 17592 16252 17714
rect 16577 17663 16635 17669
rect 16577 17629 16589 17663
rect 16623 17660 16635 17663
rect 39666 17660 39672 17672
rect 16623 17632 39672 17660
rect 16623 17629 16635 17632
rect 16577 17623 16635 17629
rect 39666 17620 39672 17632
rect 39724 17620 39730 17672
rect 17221 17595 17279 17601
rect 17221 17592 17233 17595
rect 16224 17564 17233 17592
rect 17221 17561 17233 17564
rect 17267 17592 17279 17595
rect 32306 17592 32312 17604
rect 17267 17564 32312 17592
rect 17267 17561 17279 17564
rect 17221 17555 17279 17561
rect 32306 17552 32312 17564
rect 32364 17592 32370 17604
rect 32674 17592 32680 17604
rect 32364 17564 32680 17592
rect 32364 17552 32370 17564
rect 32674 17552 32680 17564
rect 32732 17552 32738 17604
rect 17773 17527 17831 17533
rect 17773 17524 17785 17527
rect 14844 17496 17785 17524
rect 17773 17493 17785 17496
rect 17819 17524 17831 17527
rect 18046 17524 18052 17536
rect 17819 17496 18052 17524
rect 17819 17493 17831 17496
rect 17773 17487 17831 17493
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 1104 17434 18952 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 14246 17434
rect 14298 17382 14310 17434
rect 14362 17382 14374 17434
rect 14426 17382 14438 17434
rect 14490 17382 18952 17434
rect 1104 17360 18952 17382
rect 37628 17434 48852 17456
rect 37628 17382 44246 17434
rect 44298 17382 44310 17434
rect 44362 17382 44374 17434
rect 44426 17382 44438 17434
rect 44490 17382 48852 17434
rect 37628 17360 48852 17382
rect 2590 17280 2596 17332
rect 2648 17320 2654 17332
rect 40494 17320 40500 17332
rect 2648 17292 40500 17320
rect 2648 17280 2654 17292
rect 40494 17280 40500 17292
rect 40552 17280 40558 17332
rect 18046 17212 18052 17264
rect 18104 17252 18110 17264
rect 29546 17252 29552 17264
rect 18104 17224 29552 17252
rect 18104 17212 18110 17224
rect 29546 17212 29552 17224
rect 29604 17212 29610 17264
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 39666 17184 39672 17196
rect 12308 17156 39672 17184
rect 12308 17144 12314 17156
rect 39666 17144 39672 17156
rect 39724 17144 39730 17196
rect 41877 17119 41935 17125
rect 41877 17116 41889 17119
rect 39868 17088 41889 17116
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 14001 17051 14059 17057
rect 14001 17048 14013 17051
rect 13596 17020 14013 17048
rect 13596 17008 13602 17020
rect 14001 17017 14013 17020
rect 14047 17048 14059 17051
rect 31478 17048 31484 17060
rect 14047 17020 31484 17048
rect 14047 17017 14059 17020
rect 14001 17011 14059 17017
rect 31478 17008 31484 17020
rect 31536 17008 31542 17060
rect 29546 16940 29552 16992
rect 29604 16980 29610 16992
rect 39868 16989 39896 17088
rect 41877 17085 41889 17088
rect 41923 17116 41935 17119
rect 42702 17116 42708 17128
rect 41923 17088 42708 17116
rect 41923 17085 41935 17088
rect 41877 17079 41935 17085
rect 42702 17076 42708 17088
rect 42760 17076 42766 17128
rect 41690 17057 41696 17060
rect 41632 17051 41696 17057
rect 41632 17017 41644 17051
rect 41678 17017 41696 17051
rect 41632 17011 41696 17017
rect 41690 17008 41696 17011
rect 41748 17008 41754 17060
rect 39853 16983 39911 16989
rect 39853 16980 39865 16983
rect 29604 16952 39865 16980
rect 29604 16940 29610 16952
rect 39853 16949 39865 16952
rect 39899 16949 39911 16983
rect 39853 16943 39911 16949
rect 1104 16890 18952 16912
rect 1104 16838 9246 16890
rect 9298 16838 9310 16890
rect 9362 16838 9374 16890
rect 9426 16838 9438 16890
rect 9490 16838 18952 16890
rect 1104 16816 18952 16838
rect 37628 16890 48852 16912
rect 37628 16838 39246 16890
rect 39298 16838 39310 16890
rect 39362 16838 39374 16890
rect 39426 16838 39438 16890
rect 39490 16838 48852 16890
rect 37628 16816 48852 16838
rect 32306 16600 32312 16652
rect 32364 16640 32370 16652
rect 37826 16640 37832 16652
rect 32364 16612 37832 16640
rect 32364 16600 32370 16612
rect 37826 16600 37832 16612
rect 37884 16600 37890 16652
rect 27706 16572 27712 16584
rect 27667 16544 27712 16572
rect 27706 16532 27712 16544
rect 27764 16532 27770 16584
rect 1104 16346 18952 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 14246 16346
rect 14298 16294 14310 16346
rect 14362 16294 14374 16346
rect 14426 16294 14438 16346
rect 14490 16294 18952 16346
rect 1104 16272 18952 16294
rect 37628 16346 48852 16368
rect 37628 16294 44246 16346
rect 44298 16294 44310 16346
rect 44362 16294 44374 16346
rect 44426 16294 44438 16346
rect 44490 16294 48852 16346
rect 37628 16272 48852 16294
rect 18138 16232 18144 16244
rect 18099 16204 18144 16232
rect 18138 16192 18144 16204
rect 18196 16192 18202 16244
rect 43346 15988 43352 16040
rect 43404 16028 43410 16040
rect 43990 16028 43996 16040
rect 43404 16000 43996 16028
rect 43404 15988 43410 16000
rect 43990 15988 43996 16000
rect 44048 15988 44054 16040
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17276 15864 17417 15892
rect 17276 15852 17282 15864
rect 17405 15861 17417 15864
rect 17451 15892 17463 15895
rect 17862 15892 17868 15904
rect 17451 15864 17868 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 40497 15895 40555 15901
rect 40497 15861 40509 15895
rect 40543 15892 40555 15895
rect 42426 15892 42432 15904
rect 40543 15864 42432 15892
rect 40543 15861 40555 15864
rect 40497 15855 40555 15861
rect 42426 15852 42432 15864
rect 42484 15892 42490 15904
rect 42702 15892 42708 15904
rect 42484 15864 42708 15892
rect 42484 15852 42490 15864
rect 42702 15852 42708 15864
rect 42760 15852 42766 15904
rect 1104 15802 18952 15824
rect 1104 15750 9246 15802
rect 9298 15750 9310 15802
rect 9362 15750 9374 15802
rect 9426 15750 9438 15802
rect 9490 15750 18952 15802
rect 1104 15728 18952 15750
rect 37628 15802 48852 15824
rect 37628 15750 39246 15802
rect 39298 15750 39310 15802
rect 39362 15750 39374 15802
rect 39426 15750 39438 15802
rect 39490 15750 48852 15802
rect 37628 15728 48852 15750
rect 17218 15688 17224 15700
rect 17131 15660 17224 15688
rect 17218 15648 17224 15660
rect 17276 15688 17282 15700
rect 17276 15660 18092 15688
rect 17276 15648 17282 15660
rect 17954 15620 17960 15632
rect 17915 15592 17960 15620
rect 17954 15580 17960 15592
rect 18012 15580 18018 15632
rect 18064 15629 18092 15660
rect 32582 15648 32588 15700
rect 32640 15688 32646 15700
rect 43346 15688 43352 15700
rect 32640 15660 43352 15688
rect 32640 15648 32646 15660
rect 43346 15648 43352 15660
rect 43404 15648 43410 15700
rect 18049 15623 18107 15629
rect 18049 15589 18061 15623
rect 18095 15620 18107 15623
rect 18095 15592 26234 15620
rect 18095 15589 18107 15592
rect 18049 15583 18107 15589
rect 17862 15552 17868 15564
rect 17823 15524 17868 15552
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 18138 15512 18144 15564
rect 18196 15552 18202 15564
rect 18233 15555 18291 15561
rect 18233 15552 18245 15555
rect 18196 15524 18245 15552
rect 18196 15512 18202 15524
rect 18233 15521 18245 15524
rect 18279 15521 18291 15555
rect 26206 15552 26234 15592
rect 39574 15580 39580 15632
rect 39632 15620 39638 15632
rect 40773 15623 40831 15629
rect 40773 15620 40785 15623
rect 39632 15592 40785 15620
rect 39632 15580 39638 15592
rect 40773 15589 40785 15592
rect 40819 15589 40831 15623
rect 40773 15583 40831 15589
rect 47670 15552 47676 15564
rect 26206 15524 47676 15552
rect 18233 15515 18291 15521
rect 47670 15512 47676 15524
rect 47728 15512 47734 15564
rect 40770 15444 40776 15496
rect 40828 15484 40834 15496
rect 42153 15487 42211 15493
rect 42153 15484 42165 15487
rect 40828 15456 42165 15484
rect 40828 15444 40834 15456
rect 42153 15453 42165 15456
rect 42199 15453 42211 15487
rect 42426 15484 42432 15496
rect 42387 15456 42432 15484
rect 42153 15447 42211 15453
rect 42426 15444 42432 15456
rect 42484 15444 42490 15496
rect 15378 15376 15384 15428
rect 15436 15416 15442 15428
rect 17681 15419 17739 15425
rect 17681 15416 17693 15419
rect 15436 15388 17693 15416
rect 15436 15376 15442 15388
rect 17681 15385 17693 15388
rect 17727 15385 17739 15419
rect 17681 15379 17739 15385
rect 1104 15258 18952 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 14246 15258
rect 14298 15206 14310 15258
rect 14362 15206 14374 15258
rect 14426 15206 14438 15258
rect 14490 15206 18952 15258
rect 1104 15184 18952 15206
rect 37628 15258 48852 15280
rect 37628 15206 44246 15258
rect 44298 15206 44310 15258
rect 44362 15206 44374 15258
rect 44426 15206 44438 15258
rect 44490 15206 48852 15258
rect 37628 15184 48852 15206
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18141 15147 18199 15153
rect 18141 15144 18153 15147
rect 18012 15116 18153 15144
rect 18012 15104 18018 15116
rect 18141 15113 18153 15116
rect 18187 15113 18199 15147
rect 18141 15107 18199 15113
rect 40681 15147 40739 15153
rect 40681 15113 40693 15147
rect 40727 15144 40739 15147
rect 40770 15144 40776 15156
rect 40727 15116 40776 15144
rect 40727 15113 40739 15116
rect 40681 15107 40739 15113
rect 40770 15104 40776 15116
rect 40828 15104 40834 15156
rect 17681 15079 17739 15085
rect 17681 15045 17693 15079
rect 17727 15076 17739 15079
rect 19061 15079 19119 15085
rect 19061 15076 19073 15079
rect 17727 15048 19073 15076
rect 17727 15045 17739 15048
rect 17681 15039 17739 15045
rect 19061 15045 19073 15048
rect 19107 15076 19119 15079
rect 22554 15076 22560 15088
rect 19107 15048 22560 15076
rect 19107 15045 19119 15048
rect 19061 15039 19119 15045
rect 22554 15036 22560 15048
rect 22612 15036 22618 15088
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 14148 14844 17172 14872
rect 14148 14832 14154 14844
rect 17144 14813 17172 14844
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 18138 14804 18144 14816
rect 17175 14776 18144 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 1104 14714 18952 14736
rect 1104 14662 9246 14714
rect 9298 14662 9310 14714
rect 9362 14662 9374 14714
rect 9426 14662 9438 14714
rect 9490 14662 18952 14714
rect 1104 14640 18952 14662
rect 37628 14714 48852 14736
rect 37628 14662 39246 14714
rect 39298 14662 39310 14714
rect 39362 14662 39374 14714
rect 39426 14662 39438 14714
rect 39490 14662 48852 14714
rect 37628 14640 48852 14662
rect 15102 14560 15108 14612
rect 15160 14600 15166 14612
rect 22646 14600 22652 14612
rect 15160 14572 22652 14600
rect 15160 14560 15166 14572
rect 22646 14560 22652 14572
rect 22704 14560 22710 14612
rect 44634 14600 44640 14612
rect 26206 14572 44640 14600
rect 17988 14535 18046 14541
rect 17988 14501 18000 14535
rect 18034 14532 18046 14535
rect 19061 14535 19119 14541
rect 19061 14532 19073 14535
rect 18034 14504 19073 14532
rect 18034 14501 18046 14504
rect 17988 14495 18046 14501
rect 19061 14501 19073 14504
rect 19107 14501 19119 14535
rect 19061 14495 19119 14501
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 17678 14464 17684 14476
rect 17092 14436 17684 14464
rect 17092 14424 17098 14436
rect 17678 14424 17684 14436
rect 17736 14464 17742 14476
rect 26206 14464 26234 14572
rect 44634 14560 44640 14572
rect 44692 14560 44698 14612
rect 17736 14436 26234 14464
rect 17736 14424 17742 14436
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18506 14396 18512 14408
rect 18279 14368 18512 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 15378 14260 15384 14272
rect 13412 14232 15384 14260
rect 13412 14220 13418 14232
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 16022 14260 16028 14272
rect 15983 14232 16028 14260
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 16850 14260 16856 14272
rect 16763 14232 16856 14260
rect 16850 14220 16856 14232
rect 16908 14260 16914 14272
rect 24946 14260 24952 14272
rect 16908 14232 24952 14260
rect 16908 14220 16914 14232
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 1104 14170 18952 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 14246 14170
rect 14298 14118 14310 14170
rect 14362 14118 14374 14170
rect 14426 14118 14438 14170
rect 14490 14118 18952 14170
rect 1104 14096 18952 14118
rect 37628 14170 48852 14192
rect 37628 14118 44246 14170
rect 44298 14118 44310 14170
rect 44362 14118 44374 14170
rect 44426 14118 44438 14170
rect 44490 14118 48852 14170
rect 37628 14096 48852 14118
rect 12084 14028 13032 14056
rect 12084 13929 12112 14028
rect 13004 13988 13032 14028
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 14829 14059 14887 14065
rect 14829 14056 14841 14059
rect 13136 14028 14841 14056
rect 13136 14016 13142 14028
rect 14829 14025 14841 14028
rect 14875 14025 14887 14059
rect 14829 14019 14887 14025
rect 18138 14016 18144 14068
rect 18196 14056 18202 14068
rect 18506 14056 18512 14068
rect 18196 14028 18512 14056
rect 18196 14016 18202 14028
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 14090 13988 14096 14000
rect 13004 13960 14096 13988
rect 14090 13948 14096 13960
rect 14148 13948 14154 14000
rect 15197 13991 15255 13997
rect 15197 13957 15209 13991
rect 15243 13957 15255 13991
rect 15197 13951 15255 13957
rect 15335 13991 15393 13997
rect 15335 13957 15347 13991
rect 15381 13988 15393 13991
rect 16022 13988 16028 14000
rect 15381 13960 16028 13988
rect 15381 13957 15393 13960
rect 15335 13951 15393 13957
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13889 12127 13923
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 12069 13883 12127 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15212 13920 15240 13951
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 27709 13991 27767 13997
rect 27709 13988 27721 13991
rect 16448 13960 27721 13988
rect 16448 13948 16454 13960
rect 27709 13957 27721 13960
rect 27755 13957 27767 13991
rect 27709 13951 27767 13957
rect 15930 13920 15936 13932
rect 15212 13892 15936 13920
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 17218 13920 17224 13932
rect 16546 13892 17224 13920
rect 12336 13855 12394 13861
rect 12336 13821 12348 13855
rect 12382 13852 12394 13855
rect 13354 13852 13360 13864
rect 12382 13824 13360 13852
rect 12382 13821 12394 13824
rect 12336 13815 12394 13821
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 16546 13852 16574 13892
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 17678 13920 17684 13932
rect 17639 13892 17684 13920
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 18141 13923 18199 13929
rect 18141 13889 18153 13923
rect 18187 13920 18199 13923
rect 42150 13920 42156 13932
rect 18187 13892 42156 13920
rect 18187 13889 18199 13892
rect 18141 13883 18199 13889
rect 42150 13880 42156 13892
rect 42208 13880 42214 13932
rect 13464 13824 16574 13852
rect 17129 13855 17187 13861
rect 13464 13725 13492 13824
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17696 13852 17724 13880
rect 17175 13824 17724 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 17865 13855 17923 13861
rect 17865 13852 17877 13855
rect 17828 13824 17877 13852
rect 17828 13812 17834 13824
rect 17865 13821 17877 13824
rect 17911 13821 17923 13855
rect 17865 13815 17923 13821
rect 15473 13787 15531 13793
rect 15473 13753 15485 13787
rect 15519 13784 15531 13787
rect 16390 13784 16396 13796
rect 15519 13756 16396 13784
rect 15519 13753 15531 13756
rect 15473 13747 15531 13753
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 18230 13784 18236 13796
rect 18191 13756 18236 13784
rect 18230 13744 18236 13756
rect 18288 13744 18294 13796
rect 13449 13719 13507 13725
rect 13449 13685 13461 13719
rect 13495 13685 13507 13719
rect 13449 13679 13507 13685
rect 1104 13626 18952 13648
rect 1104 13574 9246 13626
rect 9298 13574 9310 13626
rect 9362 13574 9374 13626
rect 9426 13574 9438 13626
rect 9490 13574 18952 13626
rect 1104 13552 18952 13574
rect 37628 13626 48852 13648
rect 37628 13574 39246 13626
rect 39298 13574 39310 13626
rect 39362 13574 39374 13626
rect 39426 13574 39438 13626
rect 39490 13574 48852 13626
rect 37628 13552 48852 13574
rect 16390 13512 16396 13524
rect 16351 13484 16396 13512
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 31662 13404 31668 13456
rect 31720 13444 31726 13456
rect 37461 13447 37519 13453
rect 37461 13444 37473 13447
rect 31720 13416 37473 13444
rect 31720 13404 31726 13416
rect 37461 13413 37473 13416
rect 37507 13413 37519 13447
rect 37461 13407 37519 13413
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 31680 13308 31708 13404
rect 11388 13280 31708 13308
rect 11388 13268 11394 13280
rect 17402 13200 17408 13252
rect 17460 13240 17466 13252
rect 38286 13240 38292 13252
rect 17460 13212 38292 13240
rect 17460 13200 17466 13212
rect 38286 13200 38292 13212
rect 38344 13200 38350 13252
rect 15102 13132 15108 13184
rect 15160 13172 15166 13184
rect 15749 13175 15807 13181
rect 15749 13172 15761 13175
rect 15160 13144 15761 13172
rect 15160 13132 15166 13144
rect 15749 13141 15761 13144
rect 15795 13141 15807 13175
rect 15749 13135 15807 13141
rect 17681 13175 17739 13181
rect 17681 13141 17693 13175
rect 17727 13172 17739 13175
rect 17770 13172 17776 13184
rect 17727 13144 17776 13172
rect 17727 13141 17739 13144
rect 17681 13135 17739 13141
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 18230 13172 18236 13184
rect 18191 13144 18236 13172
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 1104 13082 18952 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 14246 13082
rect 14298 13030 14310 13082
rect 14362 13030 14374 13082
rect 14426 13030 14438 13082
rect 14490 13030 18952 13082
rect 1104 13008 18952 13030
rect 37628 13082 48852 13104
rect 37628 13030 44246 13082
rect 44298 13030 44310 13082
rect 44362 13030 44374 13082
rect 44426 13030 44438 13082
rect 44490 13030 48852 13082
rect 37628 13008 48852 13030
rect 38657 12971 38715 12977
rect 38657 12937 38669 12971
rect 38703 12968 38715 12971
rect 39114 12968 39120 12980
rect 38703 12940 39120 12968
rect 38703 12937 38715 12940
rect 38657 12931 38715 12937
rect 39114 12928 39120 12940
rect 39172 12928 39178 12980
rect 37461 12767 37519 12773
rect 37461 12733 37473 12767
rect 37507 12764 37519 12767
rect 38381 12767 38439 12773
rect 38381 12764 38393 12767
rect 37507 12736 38393 12764
rect 37507 12733 37519 12736
rect 37461 12727 37519 12733
rect 38381 12733 38393 12736
rect 38427 12764 38439 12767
rect 39209 12767 39267 12773
rect 39209 12764 39221 12767
rect 38427 12736 39221 12764
rect 38427 12733 38439 12736
rect 38381 12727 38439 12733
rect 39209 12733 39221 12736
rect 39255 12733 39267 12767
rect 39209 12727 39267 12733
rect 1104 12538 18952 12560
rect 1104 12486 9246 12538
rect 9298 12486 9310 12538
rect 9362 12486 9374 12538
rect 9426 12486 9438 12538
rect 9490 12486 18952 12538
rect 1104 12464 18952 12486
rect 37628 12538 48852 12560
rect 37628 12486 39246 12538
rect 39298 12486 39310 12538
rect 39362 12486 39374 12538
rect 39426 12486 39438 12538
rect 39490 12486 48852 12538
rect 37628 12464 48852 12486
rect 1854 12424 1860 12436
rect 1815 12396 1860 12424
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 11330 12424 11336 12436
rect 11291 12396 11336 12424
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 1995 12260 2636 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2608 12093 2636 12260
rect 6886 12124 16574 12152
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12084 2651 12087
rect 6886 12084 6914 12124
rect 2639 12056 6914 12084
rect 16546 12084 16574 12124
rect 16850 12084 16856 12096
rect 16546 12056 16856 12084
rect 2639 12053 2651 12056
rect 2593 12047 2651 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 1104 11994 18952 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 14246 11994
rect 14298 11942 14310 11994
rect 14362 11942 14374 11994
rect 14426 11942 14438 11994
rect 14490 11942 18952 11994
rect 1104 11920 18952 11942
rect 37628 11994 48852 12016
rect 37628 11942 44246 11994
rect 44298 11942 44310 11994
rect 44362 11942 44374 11994
rect 44426 11942 44438 11994
rect 44490 11942 48852 11994
rect 37628 11920 48852 11942
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12253 11883 12311 11889
rect 12253 11880 12265 11883
rect 12216 11852 12265 11880
rect 12216 11840 12222 11852
rect 12253 11849 12265 11852
rect 12299 11849 12311 11883
rect 12253 11843 12311 11849
rect 43438 11840 43444 11892
rect 43496 11880 43502 11892
rect 43533 11883 43591 11889
rect 43533 11880 43545 11883
rect 43496 11852 43545 11880
rect 43496 11840 43502 11852
rect 43533 11849 43545 11852
rect 43579 11849 43591 11883
rect 43533 11843 43591 11849
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 10781 11815 10839 11821
rect 10781 11812 10793 11815
rect 10744 11784 10793 11812
rect 10744 11772 10750 11784
rect 10781 11781 10793 11784
rect 10827 11781 10839 11815
rect 10781 11775 10839 11781
rect 43548 11744 43576 11843
rect 45554 11840 45560 11892
rect 45612 11880 45618 11892
rect 45649 11883 45707 11889
rect 45649 11880 45661 11883
rect 45612 11852 45661 11880
rect 45612 11840 45618 11852
rect 45649 11849 45661 11852
rect 45695 11849 45707 11883
rect 45649 11843 45707 11849
rect 44361 11747 44419 11753
rect 44361 11744 44373 11747
rect 43548 11716 44373 11744
rect 44361 11713 44373 11716
rect 44407 11713 44419 11747
rect 44361 11707 44419 11713
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 12158 11676 12164 11688
rect 10275 11648 12164 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 42426 11636 42432 11688
rect 42484 11676 42490 11688
rect 43714 11676 43720 11688
rect 42484 11648 43720 11676
rect 42484 11636 42490 11648
rect 43714 11636 43720 11648
rect 43772 11676 43778 11688
rect 44085 11679 44143 11685
rect 44085 11676 44097 11679
rect 43772 11648 44097 11676
rect 43772 11636 43778 11648
rect 44085 11645 44097 11648
rect 44131 11645 44143 11679
rect 44085 11639 44143 11645
rect 10597 11611 10655 11617
rect 10597 11577 10609 11611
rect 10643 11608 10655 11611
rect 11701 11611 11759 11617
rect 11701 11608 11713 11611
rect 10643 11580 11713 11608
rect 10643 11577 10655 11580
rect 10597 11571 10655 11577
rect 11701 11577 11713 11580
rect 11747 11608 11759 11611
rect 15102 11608 15108 11620
rect 11747 11580 15108 11608
rect 11747 11577 11759 11580
rect 11701 11571 11759 11577
rect 15102 11568 15108 11580
rect 15160 11568 15166 11620
rect 10410 11540 10416 11552
rect 10371 11512 10416 11540
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 11330 11540 11336 11552
rect 10551 11512 11336 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 1104 11450 18952 11472
rect 1104 11398 9246 11450
rect 9298 11398 9310 11450
rect 9362 11398 9374 11450
rect 9426 11398 9438 11450
rect 9490 11398 18952 11450
rect 1104 11376 18952 11398
rect 37628 11450 48852 11472
rect 37628 11398 39246 11450
rect 39298 11398 39310 11450
rect 39362 11398 39374 11450
rect 39426 11398 39438 11450
rect 39490 11398 48852 11450
rect 37628 11376 48852 11398
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10468 11308 11069 11336
rect 10468 11296 10474 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 38746 11336 38752 11348
rect 11057 11299 11115 11305
rect 38304 11308 38752 11336
rect 37734 11228 37740 11280
rect 37792 11268 37798 11280
rect 38304 11277 38332 11308
rect 38746 11296 38752 11308
rect 38804 11296 38810 11348
rect 43714 11336 43720 11348
rect 43675 11308 43720 11336
rect 43714 11296 43720 11308
rect 43772 11296 43778 11348
rect 38105 11271 38163 11277
rect 38105 11268 38117 11271
rect 37792 11240 38117 11268
rect 37792 11228 37798 11240
rect 38105 11237 38117 11240
rect 38151 11237 38163 11271
rect 38105 11231 38163 11237
rect 38289 11271 38347 11277
rect 38289 11237 38301 11271
rect 38335 11237 38347 11271
rect 38289 11231 38347 11237
rect 37918 11132 37924 11144
rect 37879 11104 37924 11132
rect 37918 11092 37924 11104
rect 37976 11092 37982 11144
rect 1104 10906 18952 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 14246 10906
rect 14298 10854 14310 10906
rect 14362 10854 14374 10906
rect 14426 10854 14438 10906
rect 14490 10854 18952 10906
rect 1104 10832 18952 10854
rect 37628 10906 48852 10928
rect 37628 10854 44246 10906
rect 44298 10854 44310 10906
rect 44362 10854 44374 10906
rect 44426 10854 44438 10906
rect 44490 10854 48852 10906
rect 37628 10832 48852 10854
rect 37734 10752 37740 10804
rect 37792 10792 37798 10804
rect 37921 10795 37979 10801
rect 37921 10792 37933 10795
rect 37792 10764 37933 10792
rect 37792 10752 37798 10764
rect 37921 10761 37933 10764
rect 37967 10761 37979 10795
rect 37921 10755 37979 10761
rect 1104 10362 18952 10384
rect 1104 10310 9246 10362
rect 9298 10310 9310 10362
rect 9362 10310 9374 10362
rect 9426 10310 9438 10362
rect 9490 10310 18952 10362
rect 1104 10288 18952 10310
rect 37628 10362 48852 10384
rect 37628 10310 39246 10362
rect 39298 10310 39310 10362
rect 39362 10310 39374 10362
rect 39426 10310 39438 10362
rect 39490 10310 48852 10362
rect 37628 10288 48852 10310
rect 1104 9818 18952 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 14246 9818
rect 14298 9766 14310 9818
rect 14362 9766 14374 9818
rect 14426 9766 14438 9818
rect 14490 9766 18952 9818
rect 1104 9744 18952 9766
rect 37628 9818 48852 9840
rect 37628 9766 44246 9818
rect 44298 9766 44310 9818
rect 44362 9766 44374 9818
rect 44426 9766 44438 9818
rect 44490 9766 48852 9818
rect 37628 9744 48852 9766
rect 32858 9324 32864 9376
rect 32916 9364 32922 9376
rect 38013 9367 38071 9373
rect 38013 9364 38025 9367
rect 32916 9336 38025 9364
rect 32916 9324 32922 9336
rect 38013 9333 38025 9336
rect 38059 9364 38071 9367
rect 47946 9364 47952 9376
rect 38059 9336 47952 9364
rect 38059 9333 38071 9336
rect 38013 9327 38071 9333
rect 47946 9324 47952 9336
rect 48004 9324 48010 9376
rect 1104 9274 18952 9296
rect 1104 9222 9246 9274
rect 9298 9222 9310 9274
rect 9362 9222 9374 9274
rect 9426 9222 9438 9274
rect 9490 9222 18952 9274
rect 1104 9200 18952 9222
rect 24028 9277 25127 9303
rect 24028 9164 24045 9277
rect 25084 9215 25127 9277
rect 24028 9163 25033 9164
rect 25085 9163 25127 9215
rect 37628 9274 48852 9296
rect 37628 9222 39246 9274
rect 39298 9222 39310 9274
rect 39362 9222 39374 9274
rect 39426 9222 39438 9274
rect 39490 9222 48852 9274
rect 37628 9200 48852 9222
rect 24028 9148 25127 9163
rect 24028 9096 24046 9148
rect 24098 9096 24101 9148
rect 24254 9096 24257 9148
rect 24408 9096 24411 9148
rect 24564 9096 24567 9148
rect 24720 9096 24723 9148
rect 24876 9096 24879 9148
rect 25030 9147 25127 9148
rect 25030 9096 25032 9147
rect 24028 9095 25032 9096
rect 25084 9095 25127 9147
rect 24028 8982 25127 9095
rect 37274 9052 37280 9104
rect 37332 9092 37338 9104
rect 45186 9092 45192 9104
rect 37332 9064 45192 9092
rect 37332 9052 37338 9064
rect 45186 9052 45192 9064
rect 45244 9052 45250 9104
rect 47489 9027 47547 9033
rect 47489 8993 47501 9027
rect 47535 9024 47547 9027
rect 48130 9024 48136 9036
rect 47535 8996 48136 9024
rect 47535 8993 47547 8996
rect 47489 8987 47547 8993
rect 48130 8984 48136 8996
rect 48188 8984 48194 9036
rect 22000 8956 25127 8982
rect 22000 8843 22032 8956
rect 22139 8955 25127 8956
rect 22251 8954 22317 8955
rect 22000 8842 22144 8843
rect 22424 8842 25127 8955
rect 22000 8841 22260 8842
rect 22312 8841 25127 8842
rect 22000 8827 25127 8841
rect 1104 8730 18952 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 14246 8730
rect 14298 8678 14310 8730
rect 14362 8678 14374 8730
rect 14426 8678 14438 8730
rect 14490 8678 18952 8730
rect 1104 8656 18952 8678
rect 22000 8664 22033 8827
rect 22140 8826 25127 8827
rect 22252 8825 22318 8826
rect 22000 8663 22145 8664
rect 22425 8663 25127 8826
rect 47946 8820 47952 8832
rect 47907 8792 47952 8820
rect 47946 8780 47952 8792
rect 48004 8780 48010 8832
rect 22000 8662 22261 8663
rect 22313 8662 25127 8663
rect 22000 8648 25127 8662
rect 37628 8730 48852 8752
rect 37628 8678 44246 8730
rect 44298 8678 44310 8730
rect 44362 8678 44374 8730
rect 44426 8678 44438 8730
rect 44490 8678 48852 8730
rect 37628 8656 48852 8678
rect 22000 8596 22034 8648
rect 22141 8647 22262 8648
rect 22314 8647 25127 8648
rect 22000 8481 22035 8596
rect 22426 8593 25127 8647
rect 22000 8480 22147 8481
rect 22254 8480 22320 8481
rect 22427 8480 25127 8593
rect 38013 8619 38071 8625
rect 38013 8585 38025 8619
rect 38059 8616 38071 8619
rect 38286 8616 38292 8628
rect 38059 8588 38292 8616
rect 38059 8585 38071 8588
rect 38013 8579 38071 8585
rect 38286 8576 38292 8588
rect 38344 8576 38350 8628
rect 38470 8576 38476 8628
rect 38528 8616 38534 8628
rect 47946 8616 47952 8628
rect 38528 8588 47952 8616
rect 38528 8576 38534 8588
rect 47946 8576 47952 8588
rect 48004 8576 48010 8628
rect 22000 8421 25127 8480
rect 17770 8304 17776 8356
rect 17828 8304 17834 8356
rect 17788 8276 17816 8304
rect 17954 8276 17960 8288
rect 17788 8248 17960 8276
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 18046 8236 18052 8288
rect 18104 8276 18110 8288
rect 18141 8279 18199 8285
rect 18141 8276 18153 8279
rect 18104 8248 18153 8276
rect 18104 8236 18110 8248
rect 18141 8245 18153 8248
rect 18187 8245 18199 8279
rect 18141 8239 18199 8245
rect 1104 8186 18952 8208
rect 1104 8134 9246 8186
rect 9298 8134 9310 8186
rect 9362 8134 9374 8186
rect 9426 8134 9438 8186
rect 9490 8134 18952 8186
rect 1104 8112 18952 8134
rect 37628 8186 48852 8208
rect 37628 8134 39246 8186
rect 39298 8134 39310 8186
rect 39362 8134 39374 8186
rect 39426 8134 39438 8186
rect 39490 8134 48852 8186
rect 37628 8112 48852 8134
rect 17402 8072 17408 8084
rect 17363 8044 17408 8072
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 34606 8032 34612 8084
rect 34664 8072 34670 8084
rect 38197 8075 38255 8081
rect 38197 8072 38209 8075
rect 34664 8044 38209 8072
rect 34664 8032 34670 8044
rect 38197 8041 38209 8044
rect 38243 8041 38255 8075
rect 38197 8035 38255 8041
rect 17420 8004 17448 8032
rect 17420 7976 18184 8004
rect 18046 7936 18052 7948
rect 18007 7908 18052 7936
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18156 7945 18184 7976
rect 37458 7964 37464 8016
rect 37516 8004 37522 8016
rect 37921 8007 37979 8013
rect 37921 8004 37933 8007
rect 37516 7976 37933 8004
rect 37516 7964 37522 7976
rect 37921 7973 37933 7976
rect 37967 7973 37979 8007
rect 38102 8004 38108 8016
rect 38063 7976 38108 8004
rect 37921 7967 37979 7973
rect 38102 7964 38108 7976
rect 38160 7964 38166 8016
rect 18141 7939 18199 7945
rect 18141 7905 18153 7939
rect 18187 7905 18199 7939
rect 38212 7936 38240 8035
rect 38286 8032 38292 8084
rect 38344 8072 38350 8084
rect 39577 8075 39635 8081
rect 39577 8072 39589 8075
rect 38344 8044 38389 8072
rect 38488 8044 39589 8072
rect 38344 8032 38350 8044
rect 38488 8013 38516 8044
rect 39577 8041 39589 8044
rect 39623 8072 39635 8075
rect 39942 8072 39948 8084
rect 39623 8044 39948 8072
rect 39623 8041 39635 8044
rect 39577 8035 39635 8041
rect 39942 8032 39948 8044
rect 40000 8032 40006 8084
rect 42150 8072 42156 8084
rect 42111 8044 42156 8072
rect 42150 8032 42156 8044
rect 42208 8032 42214 8084
rect 42610 8032 42616 8084
rect 42668 8072 42674 8084
rect 44269 8075 44327 8081
rect 44269 8072 44281 8075
rect 42668 8044 44281 8072
rect 42668 8032 42674 8044
rect 44269 8041 44281 8044
rect 44315 8041 44327 8075
rect 44269 8035 44327 8041
rect 38473 8007 38531 8013
rect 38473 7973 38485 8007
rect 38519 7973 38531 8007
rect 38473 7967 38531 7973
rect 39025 8007 39083 8013
rect 39025 7973 39037 8007
rect 39071 8004 39083 8007
rect 39114 8004 39120 8016
rect 39071 7976 39120 8004
rect 39071 7973 39083 7976
rect 39025 7967 39083 7973
rect 39040 7936 39068 7967
rect 39114 7964 39120 7976
rect 39172 7964 39178 8016
rect 38212 7908 39068 7936
rect 42168 7936 42196 8032
rect 42981 7939 43039 7945
rect 42981 7936 42993 7939
rect 42168 7908 42993 7936
rect 18141 7899 18199 7905
rect 42981 7905 42993 7908
rect 43027 7905 43039 7939
rect 42981 7899 43039 7905
rect 42426 7828 42432 7880
rect 42484 7868 42490 7880
rect 42705 7871 42763 7877
rect 42705 7868 42717 7871
rect 42484 7840 42717 7868
rect 42484 7828 42490 7840
rect 42705 7837 42717 7840
rect 42751 7837 42763 7871
rect 42705 7831 42763 7837
rect 11698 7760 11704 7812
rect 11756 7800 11762 7812
rect 17957 7803 18015 7809
rect 17957 7800 17969 7803
rect 11756 7772 17969 7800
rect 11756 7760 11762 7772
rect 17957 7769 17969 7772
rect 18003 7769 18015 7803
rect 17957 7763 18015 7769
rect 1104 7642 18952 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 14246 7642
rect 14298 7590 14310 7642
rect 14362 7590 14374 7642
rect 14426 7590 14438 7642
rect 14490 7590 18952 7642
rect 1104 7568 18952 7590
rect 37628 7642 48852 7664
rect 37628 7590 44246 7642
rect 44298 7590 44310 7642
rect 44362 7590 44374 7642
rect 44426 7590 44438 7642
rect 44490 7590 48852 7642
rect 37628 7568 48852 7590
rect 38013 7531 38071 7537
rect 38013 7497 38025 7531
rect 38059 7528 38071 7531
rect 38102 7528 38108 7540
rect 38059 7500 38108 7528
rect 38059 7497 38071 7500
rect 38013 7491 38071 7497
rect 38102 7488 38108 7500
rect 38160 7488 38166 7540
rect 38286 7488 38292 7540
rect 38344 7528 38350 7540
rect 38933 7531 38991 7537
rect 38933 7528 38945 7531
rect 38344 7500 38945 7528
rect 38344 7488 38350 7500
rect 38933 7497 38945 7500
rect 38979 7497 38991 7531
rect 38933 7491 38991 7497
rect 1762 7460 1768 7472
rect 1723 7432 1768 7460
rect 1762 7420 1768 7432
rect 1820 7420 1826 7472
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 17862 7324 17868 7336
rect 17359 7296 17868 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17862 7284 17868 7296
rect 17920 7324 17926 7336
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 17920 7296 18245 7324
rect 17920 7284 17926 7296
rect 18233 7293 18245 7296
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 11698 7256 11704 7268
rect 1995 7228 11704 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 11698 7216 11704 7228
rect 11756 7216 11762 7268
rect 17954 7256 17960 7268
rect 17867 7228 17960 7256
rect 17954 7216 17960 7228
rect 18012 7256 18018 7268
rect 21726 7256 21732 7268
rect 18012 7228 21732 7256
rect 18012 7216 18018 7228
rect 21726 7216 21732 7228
rect 21784 7216 21790 7268
rect 38948 7256 38976 7491
rect 39022 7488 39028 7540
rect 39080 7528 39086 7540
rect 39485 7531 39543 7537
rect 39485 7528 39497 7531
rect 39080 7500 39497 7528
rect 39080 7488 39086 7500
rect 39485 7497 39497 7500
rect 39531 7497 39543 7531
rect 40589 7531 40647 7537
rect 40589 7528 40601 7531
rect 39485 7491 39543 7497
rect 39592 7500 40601 7528
rect 39592 7392 39620 7500
rect 40589 7497 40601 7500
rect 40635 7528 40647 7531
rect 42610 7528 42616 7540
rect 40635 7500 42616 7528
rect 40635 7497 40647 7500
rect 40589 7491 40647 7497
rect 42610 7488 42616 7500
rect 42668 7488 42674 7540
rect 39758 7420 39764 7472
rect 39816 7460 39822 7472
rect 42426 7460 42432 7472
rect 39816 7432 39988 7460
rect 42387 7432 42432 7460
rect 39816 7420 39822 7432
rect 39960 7401 39988 7432
rect 42426 7420 42432 7432
rect 42484 7460 42490 7472
rect 43254 7460 43260 7472
rect 42484 7432 43260 7460
rect 42484 7420 42490 7432
rect 43254 7420 43260 7432
rect 43312 7420 43318 7472
rect 39669 7395 39727 7401
rect 39669 7392 39681 7395
rect 39592 7364 39681 7392
rect 39669 7361 39681 7364
rect 39715 7361 39727 7395
rect 39669 7355 39727 7361
rect 39945 7395 40003 7401
rect 39945 7361 39957 7395
rect 39991 7361 40003 7395
rect 39945 7355 40003 7361
rect 39758 7324 39764 7336
rect 39719 7296 39764 7324
rect 39758 7284 39764 7296
rect 39816 7284 39822 7336
rect 39853 7327 39911 7333
rect 39853 7293 39865 7327
rect 39899 7293 39911 7327
rect 39853 7287 39911 7293
rect 39868 7256 39896 7287
rect 38948 7228 39896 7256
rect 39114 7148 39120 7200
rect 39172 7188 39178 7200
rect 39758 7188 39764 7200
rect 39172 7160 39764 7188
rect 39172 7148 39178 7160
rect 39758 7148 39764 7160
rect 39816 7148 39822 7200
rect 1104 7098 18952 7120
rect 1104 7046 9246 7098
rect 9298 7046 9310 7098
rect 9362 7046 9374 7098
rect 9426 7046 9438 7098
rect 9490 7046 18952 7098
rect 1104 7024 18952 7046
rect 37628 7098 48852 7120
rect 37628 7046 39246 7098
rect 39298 7046 39310 7098
rect 39362 7046 39374 7098
rect 39426 7046 39438 7098
rect 39490 7046 48852 7098
rect 37628 7024 48852 7046
rect 39114 6984 39120 6996
rect 39075 6956 39120 6984
rect 39114 6944 39120 6956
rect 39172 6944 39178 6996
rect 39666 6984 39672 6996
rect 39627 6956 39672 6984
rect 39666 6944 39672 6956
rect 39724 6944 39730 6996
rect 18138 6644 18144 6656
rect 18099 6616 18144 6644
rect 18138 6604 18144 6616
rect 18196 6644 18202 6656
rect 18322 6644 18328 6656
rect 18196 6616 18328 6644
rect 18196 6604 18202 6616
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 1104 6554 18952 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 14246 6554
rect 14298 6502 14310 6554
rect 14362 6502 14374 6554
rect 14426 6502 14438 6554
rect 14490 6502 18952 6554
rect 1104 6480 18952 6502
rect 37628 6554 48852 6576
rect 37628 6502 44246 6554
rect 44298 6502 44310 6554
rect 44362 6502 44374 6554
rect 44426 6502 44438 6554
rect 44490 6502 48852 6554
rect 37628 6480 48852 6502
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7561 6443 7619 6449
rect 6972 6412 7017 6440
rect 6972 6400 6978 6412
rect 7561 6409 7573 6443
rect 7607 6440 7619 6443
rect 15930 6440 15936 6452
rect 7607 6412 15936 6440
rect 7607 6409 7619 6412
rect 7561 6403 7619 6409
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 7576 6236 7604 6403
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 38010 6440 38016 6452
rect 37971 6412 38016 6440
rect 38010 6400 38016 6412
rect 38068 6400 38074 6452
rect 6871 6208 7604 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 17954 6060 17960 6112
rect 18012 6100 18018 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 18012 6072 18245 6100
rect 18012 6060 18018 6072
rect 18233 6069 18245 6072
rect 18279 6100 18291 6103
rect 18322 6100 18328 6112
rect 18279 6072 18328 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 18322 6060 18328 6072
rect 18380 6060 18386 6112
rect 32858 6060 32864 6112
rect 32916 6100 32922 6112
rect 38470 6100 38476 6112
rect 32916 6072 38476 6100
rect 32916 6060 32922 6072
rect 38470 6060 38476 6072
rect 38528 6060 38534 6112
rect 1104 6010 18952 6032
rect 1104 5958 9246 6010
rect 9298 5958 9310 6010
rect 9362 5958 9374 6010
rect 9426 5958 9438 6010
rect 9490 5958 18952 6010
rect 1104 5936 18952 5958
rect 37628 6010 48852 6032
rect 37628 5958 39246 6010
rect 39298 5958 39310 6010
rect 39362 5958 39374 6010
rect 39426 5958 39438 6010
rect 39490 5958 48852 6010
rect 37628 5936 48852 5958
rect 18233 5899 18291 5905
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18414 5896 18420 5908
rect 18279 5868 18420 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 38013 5899 38071 5905
rect 38013 5896 38025 5899
rect 37700 5868 38025 5896
rect 37700 5856 37706 5868
rect 38013 5865 38025 5868
rect 38059 5865 38071 5899
rect 38013 5859 38071 5865
rect 18138 5828 18144 5840
rect 17604 5800 18144 5828
rect 17604 5769 17632 5800
rect 18138 5788 18144 5800
rect 18196 5788 18202 5840
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17773 5763 17831 5769
rect 17773 5729 17785 5763
rect 17819 5760 17831 5763
rect 17954 5760 17960 5772
rect 17819 5732 17960 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 18049 5763 18107 5769
rect 18049 5729 18061 5763
rect 18095 5760 18107 5763
rect 18230 5760 18236 5772
rect 18095 5732 18236 5760
rect 18095 5729 18107 5732
rect 18049 5723 18107 5729
rect 18230 5720 18236 5732
rect 18288 5760 18294 5772
rect 23934 5760 23940 5772
rect 18288 5732 23940 5760
rect 18288 5720 18294 5732
rect 23934 5720 23940 5732
rect 23992 5720 23998 5772
rect 33870 5720 33876 5772
rect 33928 5760 33934 5772
rect 38105 5763 38163 5769
rect 38105 5760 38117 5763
rect 33928 5732 38117 5760
rect 33928 5720 33934 5732
rect 38105 5729 38117 5732
rect 38151 5760 38163 5763
rect 38565 5763 38623 5769
rect 38565 5760 38577 5763
rect 38151 5732 38577 5760
rect 38151 5729 38163 5732
rect 38105 5723 38163 5729
rect 38565 5729 38577 5732
rect 38611 5729 38623 5763
rect 38565 5723 38623 5729
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5692 17187 5695
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17175 5664 17877 5692
rect 17175 5661 17187 5664
rect 17129 5655 17187 5661
rect 17865 5661 17877 5664
rect 17911 5692 17923 5695
rect 24946 5692 24952 5704
rect 17911 5664 24952 5692
rect 17911 5661 17923 5664
rect 17865 5655 17923 5661
rect 24946 5652 24952 5664
rect 25004 5652 25010 5704
rect 17954 5584 17960 5636
rect 18012 5624 18018 5636
rect 18012 5596 18057 5624
rect 18012 5584 18018 5596
rect 1104 5466 18952 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 14246 5466
rect 14298 5414 14310 5466
rect 14362 5414 14374 5466
rect 14426 5414 14438 5466
rect 14490 5414 18952 5466
rect 1104 5392 18952 5414
rect 37628 5466 48852 5488
rect 37628 5414 44246 5466
rect 44298 5414 44310 5466
rect 44362 5414 44374 5466
rect 44426 5414 44438 5466
rect 44490 5414 48852 5466
rect 37628 5392 48852 5414
rect 38473 5355 38531 5361
rect 38473 5321 38485 5355
rect 38519 5352 38531 5355
rect 38562 5352 38568 5364
rect 38519 5324 38568 5352
rect 38519 5321 38531 5324
rect 38473 5315 38531 5321
rect 38562 5312 38568 5324
rect 38620 5312 38626 5364
rect 17681 5287 17739 5293
rect 17681 5253 17693 5287
rect 17727 5284 17739 5287
rect 18046 5284 18052 5296
rect 17727 5256 18052 5284
rect 17727 5253 17739 5256
rect 17681 5247 17739 5253
rect 18046 5244 18052 5256
rect 18104 5284 18110 5296
rect 23750 5284 23756 5296
rect 18104 5256 23756 5284
rect 18104 5244 18110 5256
rect 23750 5244 23756 5256
rect 23808 5244 23814 5296
rect 37274 5176 37280 5228
rect 37332 5216 37338 5228
rect 37332 5188 38332 5216
rect 37332 5176 37338 5188
rect 38304 5160 38332 5188
rect 37921 5151 37979 5157
rect 37921 5117 37933 5151
rect 37967 5148 37979 5151
rect 38010 5148 38016 5160
rect 37967 5120 38016 5148
rect 37967 5117 37979 5120
rect 37921 5111 37979 5117
rect 38010 5108 38016 5120
rect 38068 5108 38074 5160
rect 38102 5108 38108 5160
rect 38160 5148 38166 5160
rect 38286 5148 38292 5160
rect 38160 5120 38205 5148
rect 38247 5120 38292 5148
rect 38160 5108 38166 5120
rect 38286 5108 38292 5120
rect 38344 5108 38350 5160
rect 38197 5083 38255 5089
rect 38197 5049 38209 5083
rect 38243 5080 38255 5083
rect 38838 5080 38844 5092
rect 38243 5052 38844 5080
rect 38243 5049 38255 5052
rect 38197 5043 38255 5049
rect 38838 5040 38844 5052
rect 38896 5080 38902 5092
rect 38896 5052 39068 5080
rect 38896 5040 38902 5052
rect 39040 5024 39068 5052
rect 17954 4972 17960 5024
rect 18012 5012 18018 5024
rect 18233 5015 18291 5021
rect 18233 5012 18245 5015
rect 18012 4984 18245 5012
rect 18012 4972 18018 4984
rect 18233 4981 18245 4984
rect 18279 5012 18291 5015
rect 35250 5012 35256 5024
rect 18279 4984 35256 5012
rect 18279 4981 18291 4984
rect 18233 4975 18291 4981
rect 35250 4972 35256 4984
rect 35308 4972 35314 5024
rect 39022 5012 39028 5024
rect 38983 4984 39028 5012
rect 39022 4972 39028 4984
rect 39080 4972 39086 5024
rect 1104 4922 18952 4944
rect 1104 4870 9246 4922
rect 9298 4870 9310 4922
rect 9362 4870 9374 4922
rect 9426 4870 9438 4922
rect 9490 4870 18952 4922
rect 1104 4848 18952 4870
rect 37628 4922 48852 4944
rect 37628 4870 39246 4922
rect 39298 4870 39310 4922
rect 39362 4870 39374 4922
rect 39426 4870 39438 4922
rect 39490 4870 48852 4922
rect 37628 4848 48852 4870
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 38013 4811 38071 4817
rect 38013 4777 38025 4811
rect 38059 4808 38071 4811
rect 38102 4808 38108 4820
rect 38059 4780 38108 4808
rect 38059 4777 38071 4780
rect 38013 4771 38071 4777
rect 38102 4768 38108 4780
rect 38160 4768 38166 4820
rect 1104 4378 18952 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 14246 4378
rect 14298 4326 14310 4378
rect 14362 4326 14374 4378
rect 14426 4326 14438 4378
rect 14490 4326 18952 4378
rect 1104 4304 18952 4326
rect 37628 4378 48852 4400
rect 37628 4326 44246 4378
rect 44298 4326 44310 4378
rect 44362 4326 44374 4378
rect 44426 4326 44438 4378
rect 44490 4326 48852 4378
rect 37628 4304 48852 4326
rect 38013 4267 38071 4273
rect 38013 4233 38025 4267
rect 38059 4264 38071 4267
rect 38286 4264 38292 4276
rect 38059 4236 38292 4264
rect 38059 4233 38071 4236
rect 38013 4227 38071 4233
rect 38286 4224 38292 4236
rect 38344 4224 38350 4276
rect 43530 4128 43536 4140
rect 43491 4100 43536 4128
rect 43530 4088 43536 4100
rect 43588 4088 43594 4140
rect 44177 4131 44235 4137
rect 44177 4097 44189 4131
rect 44223 4128 44235 4131
rect 44634 4128 44640 4140
rect 44223 4100 44640 4128
rect 44223 4097 44235 4100
rect 44177 4091 44235 4097
rect 44634 4088 44640 4100
rect 44692 4088 44698 4140
rect 41601 3995 41659 4001
rect 41601 3992 41613 3995
rect 22066 3964 41613 3992
rect 1104 3834 18952 3856
rect 1104 3782 9246 3834
rect 9298 3782 9310 3834
rect 9362 3782 9374 3834
rect 9426 3782 9438 3834
rect 9490 3782 18952 3834
rect 1104 3760 18952 3782
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 22066 3584 22094 3964
rect 41601 3961 41613 3964
rect 41647 3992 41659 3995
rect 42334 3992 42340 4004
rect 41647 3964 42340 3992
rect 41647 3961 41659 3964
rect 41601 3955 41659 3961
rect 42334 3952 42340 3964
rect 42392 3952 42398 4004
rect 37628 3834 48852 3856
rect 37628 3782 39246 3834
rect 39298 3782 39310 3834
rect 39362 3782 39374 3834
rect 39426 3782 39438 3834
rect 39490 3782 48852 3834
rect 37628 3760 48852 3782
rect 41046 3720 41052 3732
rect 41007 3692 41052 3720
rect 41046 3680 41052 3692
rect 41104 3680 41110 3732
rect 41598 3720 41604 3732
rect 41559 3692 41604 3720
rect 41598 3680 41604 3692
rect 41656 3720 41662 3732
rect 42518 3720 42524 3732
rect 41656 3692 42524 3720
rect 41656 3680 41662 3692
rect 42518 3680 42524 3692
rect 42576 3680 42582 3732
rect 42794 3720 42800 3732
rect 42755 3692 42800 3720
rect 42794 3680 42800 3692
rect 42852 3680 42858 3732
rect 43346 3720 43352 3732
rect 43307 3692 43352 3720
rect 43346 3680 43352 3692
rect 43404 3680 43410 3732
rect 44453 3723 44511 3729
rect 44453 3689 44465 3723
rect 44499 3720 44511 3723
rect 44542 3720 44548 3732
rect 44499 3692 44548 3720
rect 44499 3689 44511 3692
rect 44453 3683 44511 3689
rect 44542 3680 44548 3692
rect 44600 3680 44606 3732
rect 41064 3652 41092 3680
rect 41064 3624 42656 3652
rect 18380 3556 22094 3584
rect 18380 3544 18386 3556
rect 41230 3544 41236 3596
rect 41288 3584 41294 3596
rect 42153 3587 42211 3593
rect 42153 3584 42165 3587
rect 41288 3556 42165 3584
rect 41288 3544 41294 3556
rect 42153 3553 42165 3556
rect 42199 3553 42211 3587
rect 42334 3584 42340 3596
rect 42295 3556 42340 3584
rect 42153 3547 42211 3553
rect 42334 3544 42340 3556
rect 42392 3544 42398 3596
rect 42518 3584 42524 3596
rect 42479 3556 42524 3584
rect 42518 3544 42524 3556
rect 42576 3544 42582 3596
rect 42628 3593 42656 3624
rect 43530 3612 43536 3664
rect 43588 3652 43594 3664
rect 43588 3624 44956 3652
rect 43588 3612 43594 3624
rect 42613 3587 42671 3593
rect 42613 3553 42625 3587
rect 42659 3553 42671 3587
rect 44634 3584 44640 3596
rect 44595 3556 44640 3584
rect 42613 3547 42671 3553
rect 44634 3544 44640 3556
rect 44692 3544 44698 3596
rect 44928 3593 44956 3624
rect 44913 3587 44971 3593
rect 44913 3553 44925 3587
rect 44959 3553 44971 3587
rect 44913 3547 44971 3553
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 13722 3516 13728 3528
rect 12492 3488 13728 3516
rect 12492 3476 12498 3488
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 35250 3476 35256 3528
rect 35308 3516 35314 3528
rect 43901 3519 43959 3525
rect 43901 3516 43913 3519
rect 35308 3488 43913 3516
rect 35308 3476 35314 3488
rect 43901 3485 43913 3488
rect 43947 3516 43959 3519
rect 44729 3519 44787 3525
rect 44729 3516 44741 3519
rect 43947 3488 44741 3516
rect 43947 3485 43959 3488
rect 43901 3479 43959 3485
rect 44729 3485 44741 3488
rect 44775 3485 44787 3519
rect 44729 3479 44787 3485
rect 42426 3448 42432 3460
rect 42387 3420 42432 3448
rect 42426 3408 42432 3420
rect 42484 3408 42490 3460
rect 43346 3408 43352 3460
rect 43404 3448 43410 3460
rect 44821 3451 44879 3457
rect 44821 3448 44833 3451
rect 43404 3420 44833 3448
rect 43404 3408 43410 3420
rect 44821 3417 44833 3420
rect 44867 3417 44879 3451
rect 44821 3411 44879 3417
rect 1104 3290 18952 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 14246 3290
rect 14298 3238 14310 3290
rect 14362 3238 14374 3290
rect 14426 3238 14438 3290
rect 14490 3238 18952 3290
rect 1104 3216 18952 3238
rect 37628 3290 48852 3312
rect 37628 3238 44246 3290
rect 44298 3238 44310 3290
rect 44362 3238 44374 3290
rect 44426 3238 44438 3290
rect 44490 3238 48852 3290
rect 37628 3216 48852 3238
rect 10594 3176 10600 3188
rect 10555 3148 10600 3176
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 41230 3176 41236 3188
rect 41191 3148 41236 3176
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 32950 3068 32956 3120
rect 33008 3108 33014 3120
rect 41785 3111 41843 3117
rect 41785 3108 41797 3111
rect 33008 3080 41797 3108
rect 33008 3068 33014 3080
rect 41785 3077 41797 3080
rect 41831 3108 41843 3111
rect 42426 3108 42432 3120
rect 41831 3080 42432 3108
rect 41831 3077 41843 3080
rect 41785 3071 41843 3077
rect 42426 3068 42432 3080
rect 42484 3068 42490 3120
rect 39022 3040 39028 3052
rect 22066 3012 39028 3040
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 10870 2972 10876 2984
rect 10735 2944 10876 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 10870 2932 10876 2944
rect 10928 2972 10934 2984
rect 22066 2972 22094 3012
rect 39022 3000 39028 3012
rect 39080 3040 39086 3052
rect 43349 3043 43407 3049
rect 43349 3040 43361 3043
rect 39080 3012 43361 3040
rect 39080 3000 39086 3012
rect 43349 3009 43361 3012
rect 43395 3009 43407 3043
rect 43349 3003 43407 3009
rect 44729 3043 44787 3049
rect 44729 3009 44741 3043
rect 44775 3040 44787 3043
rect 45557 3043 45615 3049
rect 45557 3040 45569 3043
rect 44775 3012 45569 3040
rect 44775 3009 44787 3012
rect 44729 3003 44787 3009
rect 45557 3009 45569 3012
rect 45603 3040 45615 3043
rect 46198 3040 46204 3052
rect 45603 3012 46204 3040
rect 45603 3009 45615 3012
rect 45557 3003 45615 3009
rect 46198 3000 46204 3012
rect 46256 3000 46262 3052
rect 10928 2944 22094 2972
rect 10928 2932 10934 2944
rect 43254 2932 43260 2984
rect 43312 2972 43318 2984
rect 45005 2975 45063 2981
rect 45005 2972 45017 2975
rect 43312 2944 45017 2972
rect 43312 2932 43318 2944
rect 45005 2941 45017 2944
rect 45051 2941 45063 2975
rect 45005 2935 45063 2941
rect 37918 2836 37924 2848
rect 37879 2808 37924 2836
rect 37918 2796 37924 2808
rect 37976 2796 37982 2848
rect 1104 2746 18952 2768
rect 1104 2694 9246 2746
rect 9298 2694 9310 2746
rect 9362 2694 9374 2746
rect 9426 2694 9438 2746
rect 9490 2694 18952 2746
rect 1104 2672 18952 2694
rect 37628 2746 48852 2768
rect 37628 2694 39246 2746
rect 39298 2694 39310 2746
rect 39362 2694 39374 2746
rect 39426 2694 39438 2746
rect 39490 2694 48852 2746
rect 37628 2672 48852 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 3602 2632 3608 2644
rect 1627 2604 3608 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 3602 2592 3608 2604
rect 3660 2592 3666 2644
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 37826 2592 37832 2644
rect 37884 2632 37890 2644
rect 38105 2635 38163 2641
rect 38105 2632 38117 2635
rect 37884 2604 38117 2632
rect 37884 2592 37890 2604
rect 38105 2601 38117 2604
rect 38151 2601 38163 2635
rect 43254 2632 43260 2644
rect 43215 2604 43260 2632
rect 38105 2595 38163 2601
rect 43254 2592 43260 2604
rect 43312 2592 43318 2644
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2496 1458 2508
rect 2041 2499 2099 2505
rect 2041 2496 2053 2499
rect 1452 2468 2053 2496
rect 1452 2456 1458 2468
rect 2041 2465 2053 2468
rect 2087 2465 2099 2499
rect 2041 2459 2099 2465
rect 37366 2456 37372 2508
rect 37424 2496 37430 2508
rect 37918 2496 37924 2508
rect 37424 2468 37924 2496
rect 37424 2456 37430 2468
rect 37918 2456 37924 2468
rect 37976 2456 37982 2508
rect 1104 2202 18952 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 14246 2202
rect 14298 2150 14310 2202
rect 14362 2150 14374 2202
rect 14426 2150 14438 2202
rect 14490 2150 18952 2202
rect 1104 2128 18952 2150
rect 37628 2202 48852 2224
rect 37628 2150 44246 2202
rect 44298 2150 44310 2202
rect 44362 2150 44374 2202
rect 44426 2150 44438 2202
rect 44490 2150 48852 2202
rect 37628 2128 48852 2150
<< via1 >>
rect 9246 47302 9298 47354
rect 9310 47302 9362 47354
rect 9374 47302 9426 47354
rect 9438 47302 9490 47354
rect 19246 47302 19298 47354
rect 19310 47302 19362 47354
rect 19374 47302 19426 47354
rect 19438 47302 19490 47354
rect 29246 47302 29298 47354
rect 29310 47302 29362 47354
rect 29374 47302 29426 47354
rect 29438 47302 29490 47354
rect 39246 47302 39298 47354
rect 39310 47302 39362 47354
rect 39374 47302 39426 47354
rect 39438 47302 39490 47354
rect 1860 47243 1912 47252
rect 1860 47209 1869 47243
rect 1869 47209 1903 47243
rect 1903 47209 1912 47243
rect 1860 47200 1912 47209
rect 17316 47064 17368 47116
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 14246 46758 14298 46810
rect 14310 46758 14362 46810
rect 14374 46758 14426 46810
rect 14438 46758 14490 46810
rect 24246 46758 24298 46810
rect 24310 46758 24362 46810
rect 24374 46758 24426 46810
rect 24438 46758 24490 46810
rect 34246 46758 34298 46810
rect 34310 46758 34362 46810
rect 34374 46758 34426 46810
rect 34438 46758 34490 46810
rect 44246 46758 44298 46810
rect 44310 46758 44362 46810
rect 44374 46758 44426 46810
rect 44438 46758 44490 46810
rect 9246 46214 9298 46266
rect 9310 46214 9362 46266
rect 9374 46214 9426 46266
rect 9438 46214 9490 46266
rect 19246 46214 19298 46266
rect 19310 46214 19362 46266
rect 19374 46214 19426 46266
rect 19438 46214 19490 46266
rect 29246 46214 29298 46266
rect 29310 46214 29362 46266
rect 29374 46214 29426 46266
rect 29438 46214 29490 46266
rect 39246 46214 39298 46266
rect 39310 46214 39362 46266
rect 39374 46214 39426 46266
rect 39438 46214 39490 46266
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 14246 45670 14298 45722
rect 14310 45670 14362 45722
rect 14374 45670 14426 45722
rect 14438 45670 14490 45722
rect 24246 45670 24298 45722
rect 24310 45670 24362 45722
rect 24374 45670 24426 45722
rect 24438 45670 24490 45722
rect 34246 45670 34298 45722
rect 34310 45670 34362 45722
rect 34374 45670 34426 45722
rect 34438 45670 34490 45722
rect 44246 45670 44298 45722
rect 44310 45670 44362 45722
rect 44374 45670 44426 45722
rect 44438 45670 44490 45722
rect 19984 45432 20036 45484
rect 2872 45228 2924 45280
rect 25780 45296 25832 45348
rect 9246 45126 9298 45178
rect 9310 45126 9362 45178
rect 9374 45126 9426 45178
rect 9438 45126 9490 45178
rect 19246 45126 19298 45178
rect 19310 45126 19362 45178
rect 19374 45126 19426 45178
rect 19438 45126 19490 45178
rect 29246 45126 29298 45178
rect 29310 45126 29362 45178
rect 29374 45126 29426 45178
rect 29438 45126 29490 45178
rect 39246 45126 39298 45178
rect 39310 45126 39362 45178
rect 39374 45126 39426 45178
rect 39438 45126 39490 45178
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 14246 44582 14298 44634
rect 14310 44582 14362 44634
rect 14374 44582 14426 44634
rect 14438 44582 14490 44634
rect 24246 44582 24298 44634
rect 24310 44582 24362 44634
rect 24374 44582 24426 44634
rect 24438 44582 24490 44634
rect 34246 44582 34298 44634
rect 34310 44582 34362 44634
rect 34374 44582 34426 44634
rect 34438 44582 34490 44634
rect 44246 44582 44298 44634
rect 44310 44582 44362 44634
rect 44374 44582 44426 44634
rect 44438 44582 44490 44634
rect 9246 44038 9298 44090
rect 9310 44038 9362 44090
rect 9374 44038 9426 44090
rect 9438 44038 9490 44090
rect 19246 44038 19298 44090
rect 19310 44038 19362 44090
rect 19374 44038 19426 44090
rect 19438 44038 19490 44090
rect 29246 44038 29298 44090
rect 29310 44038 29362 44090
rect 29374 44038 29426 44090
rect 29438 44038 29490 44090
rect 39246 44038 39298 44090
rect 39310 44038 39362 44090
rect 39374 44038 39426 44090
rect 39438 44038 39490 44090
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 14246 43494 14298 43546
rect 14310 43494 14362 43546
rect 14374 43494 14426 43546
rect 14438 43494 14490 43546
rect 24246 43494 24298 43546
rect 24310 43494 24362 43546
rect 24374 43494 24426 43546
rect 24438 43494 24490 43546
rect 34246 43494 34298 43546
rect 34310 43494 34362 43546
rect 34374 43494 34426 43546
rect 34438 43494 34490 43546
rect 44246 43494 44298 43546
rect 44310 43494 44362 43546
rect 44374 43494 44426 43546
rect 44438 43494 44490 43546
rect 9246 42950 9298 43002
rect 9310 42950 9362 43002
rect 9374 42950 9426 43002
rect 9438 42950 9490 43002
rect 19246 42950 19298 43002
rect 19310 42950 19362 43002
rect 19374 42950 19426 43002
rect 19438 42950 19490 43002
rect 29246 42950 29298 43002
rect 29310 42950 29362 43002
rect 29374 42950 29426 43002
rect 29438 42950 29490 43002
rect 39246 42950 39298 43002
rect 39310 42950 39362 43002
rect 39374 42950 39426 43002
rect 39438 42950 39490 43002
rect 1860 42551 1912 42560
rect 1860 42517 1869 42551
rect 1869 42517 1903 42551
rect 1903 42517 1912 42551
rect 1860 42508 1912 42517
rect 39672 42712 39724 42764
rect 35348 42644 35400 42696
rect 42800 42712 42852 42764
rect 43352 42687 43404 42696
rect 38936 42576 38988 42628
rect 43352 42653 43361 42687
rect 43361 42653 43395 42687
rect 43395 42653 43404 42687
rect 43352 42644 43404 42653
rect 12256 42508 12308 42560
rect 42800 42551 42852 42560
rect 42800 42517 42809 42551
rect 42809 42517 42843 42551
rect 42843 42517 42852 42551
rect 42800 42508 42852 42517
rect 43260 42576 43312 42628
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 14246 42406 14298 42458
rect 14310 42406 14362 42458
rect 14374 42406 14426 42458
rect 14438 42406 14490 42458
rect 24246 42406 24298 42458
rect 24310 42406 24362 42458
rect 24374 42406 24426 42458
rect 24438 42406 24490 42458
rect 34246 42406 34298 42458
rect 34310 42406 34362 42458
rect 34374 42406 34426 42458
rect 34438 42406 34490 42458
rect 44246 42406 44298 42458
rect 44310 42406 44362 42458
rect 44374 42406 44426 42458
rect 44438 42406 44490 42458
rect 40684 41964 40736 42016
rect 43352 41964 43404 42016
rect 9246 41862 9298 41914
rect 9310 41862 9362 41914
rect 9374 41862 9426 41914
rect 9438 41862 9490 41914
rect 19246 41862 19298 41914
rect 19310 41862 19362 41914
rect 19374 41862 19426 41914
rect 19438 41862 19490 41914
rect 29246 41862 29298 41914
rect 29310 41862 29362 41914
rect 29374 41862 29426 41914
rect 29438 41862 29490 41914
rect 39246 41862 39298 41914
rect 39310 41862 39362 41914
rect 39374 41862 39426 41914
rect 39438 41862 39490 41914
rect 39672 41692 39724 41744
rect 13084 41624 13136 41676
rect 13636 41599 13688 41608
rect 13636 41565 13645 41599
rect 13645 41565 13679 41599
rect 13679 41565 13688 41599
rect 13636 41556 13688 41565
rect 15108 41488 15160 41540
rect 6736 41463 6788 41472
rect 6736 41429 6745 41463
rect 6745 41429 6779 41463
rect 6779 41429 6788 41463
rect 6736 41420 6788 41429
rect 44548 41420 44600 41472
rect 48136 41667 48188 41676
rect 48136 41633 48145 41667
rect 48145 41633 48179 41667
rect 48179 41633 48188 41667
rect 48136 41624 48188 41633
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 14246 41318 14298 41370
rect 14310 41318 14362 41370
rect 14374 41318 14426 41370
rect 14438 41318 14490 41370
rect 24246 41318 24298 41370
rect 24310 41318 24362 41370
rect 24374 41318 24426 41370
rect 24438 41318 24490 41370
rect 34246 41318 34298 41370
rect 34310 41318 34362 41370
rect 34374 41318 34426 41370
rect 34438 41318 34490 41370
rect 44246 41318 44298 41370
rect 44310 41318 44362 41370
rect 44374 41318 44426 41370
rect 44438 41318 44490 41370
rect 13084 40876 13136 40928
rect 9246 40774 9298 40826
rect 9310 40774 9362 40826
rect 9374 40774 9426 40826
rect 9438 40774 9490 40826
rect 19246 40774 19298 40826
rect 19310 40774 19362 40826
rect 19374 40774 19426 40826
rect 19438 40774 19490 40826
rect 29246 40774 29298 40826
rect 29310 40774 29362 40826
rect 29374 40774 29426 40826
rect 29438 40774 29490 40826
rect 39246 40774 39298 40826
rect 39310 40774 39362 40826
rect 39374 40774 39426 40826
rect 39438 40774 39490 40826
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 14246 40230 14298 40282
rect 14310 40230 14362 40282
rect 14374 40230 14426 40282
rect 14438 40230 14490 40282
rect 24246 40230 24298 40282
rect 24310 40230 24362 40282
rect 24374 40230 24426 40282
rect 24438 40230 24490 40282
rect 34246 40230 34298 40282
rect 34310 40230 34362 40282
rect 34374 40230 34426 40282
rect 34438 40230 34490 40282
rect 44246 40230 44298 40282
rect 44310 40230 44362 40282
rect 44374 40230 44426 40282
rect 44438 40230 44490 40282
rect 9246 39686 9298 39738
rect 9310 39686 9362 39738
rect 9374 39686 9426 39738
rect 9438 39686 9490 39738
rect 19246 39686 19298 39738
rect 19310 39686 19362 39738
rect 19374 39686 19426 39738
rect 19438 39686 19490 39738
rect 29246 39686 29298 39738
rect 29310 39686 29362 39738
rect 29374 39686 29426 39738
rect 29438 39686 29490 39738
rect 39246 39686 39298 39738
rect 39310 39686 39362 39738
rect 39374 39686 39426 39738
rect 39438 39686 39490 39738
rect 15108 39516 15160 39568
rect 35348 39584 35400 39636
rect 23112 39491 23164 39500
rect 21916 39423 21968 39432
rect 21916 39389 21925 39423
rect 21925 39389 21959 39423
rect 21959 39389 21968 39423
rect 21916 39380 21968 39389
rect 23112 39457 23121 39491
rect 23121 39457 23155 39491
rect 23155 39457 23164 39491
rect 23112 39448 23164 39457
rect 22744 39355 22796 39364
rect 22744 39321 22753 39355
rect 22753 39321 22787 39355
rect 22787 39321 22796 39355
rect 22744 39312 22796 39321
rect 22560 39244 22612 39296
rect 23664 39287 23716 39296
rect 23664 39253 23673 39287
rect 23673 39253 23707 39287
rect 23707 39253 23716 39287
rect 23664 39244 23716 39253
rect 24584 39244 24636 39296
rect 24768 39244 24820 39296
rect 43996 39244 44048 39296
rect 44548 39244 44600 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 14246 39142 14298 39194
rect 14310 39142 14362 39194
rect 14374 39142 14426 39194
rect 14438 39142 14490 39194
rect 24246 39142 24298 39194
rect 24310 39142 24362 39194
rect 24374 39142 24426 39194
rect 24438 39142 24490 39194
rect 34246 39142 34298 39194
rect 34310 39142 34362 39194
rect 34374 39142 34426 39194
rect 34438 39142 34490 39194
rect 44246 39142 44298 39194
rect 44310 39142 44362 39194
rect 44374 39142 44426 39194
rect 44438 39142 44490 39194
rect 24584 39040 24636 39092
rect 39672 39040 39724 39092
rect 23664 38972 23716 39024
rect 32864 38972 32916 39024
rect 24676 38879 24728 38888
rect 24676 38845 24685 38879
rect 24685 38845 24719 38879
rect 24719 38845 24728 38879
rect 24676 38836 24728 38845
rect 32864 38836 32916 38888
rect 33508 38879 33560 38888
rect 33508 38845 33517 38879
rect 33517 38845 33551 38879
rect 33551 38845 33560 38879
rect 33508 38836 33560 38845
rect 22744 38700 22796 38752
rect 24768 38768 24820 38820
rect 33232 38811 33284 38820
rect 33232 38777 33241 38811
rect 33241 38777 33275 38811
rect 33275 38777 33284 38811
rect 33232 38768 33284 38777
rect 23940 38700 23992 38752
rect 29092 38743 29144 38752
rect 29092 38709 29101 38743
rect 29101 38709 29135 38743
rect 29135 38709 29144 38743
rect 29092 38700 29144 38709
rect 9246 38598 9298 38650
rect 9310 38598 9362 38650
rect 9374 38598 9426 38650
rect 9438 38598 9490 38650
rect 19246 38598 19298 38650
rect 19310 38598 19362 38650
rect 19374 38598 19426 38650
rect 19438 38598 19490 38650
rect 29246 38598 29298 38650
rect 29310 38598 29362 38650
rect 29374 38598 29426 38650
rect 29438 38598 29490 38650
rect 39246 38598 39298 38650
rect 39310 38598 39362 38650
rect 39374 38598 39426 38650
rect 39438 38598 39490 38650
rect 32864 38539 32916 38548
rect 32864 38505 32873 38539
rect 32873 38505 32907 38539
rect 32907 38505 32916 38539
rect 32864 38496 32916 38505
rect 16948 38428 17000 38480
rect 5172 38403 5224 38412
rect 5172 38369 5181 38403
rect 5181 38369 5215 38403
rect 5215 38369 5224 38403
rect 5172 38360 5224 38369
rect 9864 38292 9916 38344
rect 24124 38360 24176 38412
rect 29092 38292 29144 38344
rect 27712 38199 27764 38208
rect 27712 38165 27721 38199
rect 27721 38165 27755 38199
rect 27755 38165 27764 38199
rect 27712 38156 27764 38165
rect 28080 38199 28132 38208
rect 28080 38165 28089 38199
rect 28089 38165 28123 38199
rect 28123 38165 28132 38199
rect 28080 38156 28132 38165
rect 29000 38156 29052 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 14246 38054 14298 38106
rect 14310 38054 14362 38106
rect 14374 38054 14426 38106
rect 14438 38054 14490 38106
rect 24246 38054 24298 38106
rect 24310 38054 24362 38106
rect 24374 38054 24426 38106
rect 24438 38054 24490 38106
rect 34246 38054 34298 38106
rect 34310 38054 34362 38106
rect 34374 38054 34426 38106
rect 34438 38054 34490 38106
rect 44246 38054 44298 38106
rect 44310 38054 44362 38106
rect 44374 38054 44426 38106
rect 44438 38054 44490 38106
rect 29092 37884 29144 37936
rect 42064 37884 42116 37936
rect 28080 37612 28132 37664
rect 39120 37612 39172 37664
rect 9246 37510 9298 37562
rect 9310 37510 9362 37562
rect 9374 37510 9426 37562
rect 9438 37510 9490 37562
rect 19246 37510 19298 37562
rect 19310 37510 19362 37562
rect 19374 37510 19426 37562
rect 19438 37510 19490 37562
rect 29246 37510 29298 37562
rect 29310 37510 29362 37562
rect 29374 37510 29426 37562
rect 29438 37510 29490 37562
rect 39246 37510 39298 37562
rect 39310 37510 39362 37562
rect 39374 37510 39426 37562
rect 39438 37510 39490 37562
rect 1860 37451 1912 37460
rect 1860 37417 1869 37451
rect 1869 37417 1903 37451
rect 1903 37417 1912 37451
rect 1860 37408 1912 37417
rect 38936 37272 38988 37324
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 14246 36966 14298 37018
rect 14310 36966 14362 37018
rect 14374 36966 14426 37018
rect 14438 36966 14490 37018
rect 24246 36966 24298 37018
rect 24310 36966 24362 37018
rect 24374 36966 24426 37018
rect 24438 36966 24490 37018
rect 34246 36966 34298 37018
rect 34310 36966 34362 37018
rect 34374 36966 34426 37018
rect 34438 36966 34490 37018
rect 44246 36966 44298 37018
rect 44310 36966 44362 37018
rect 44374 36966 44426 37018
rect 44438 36966 44490 37018
rect 11704 36796 11756 36848
rect 19984 36864 20036 36916
rect 13360 36567 13412 36576
rect 13360 36533 13369 36567
rect 13369 36533 13403 36567
rect 13403 36533 13412 36567
rect 13360 36524 13412 36533
rect 17040 36567 17092 36576
rect 17040 36533 17049 36567
rect 17049 36533 17083 36567
rect 17083 36533 17092 36567
rect 17040 36524 17092 36533
rect 9246 36422 9298 36474
rect 9310 36422 9362 36474
rect 9374 36422 9426 36474
rect 9438 36422 9490 36474
rect 19246 36422 19298 36474
rect 19310 36422 19362 36474
rect 19374 36422 19426 36474
rect 19438 36422 19490 36474
rect 29246 36422 29298 36474
rect 29310 36422 29362 36474
rect 29374 36422 29426 36474
rect 29438 36422 29490 36474
rect 39246 36422 39298 36474
rect 39310 36422 39362 36474
rect 39374 36422 39426 36474
rect 39438 36422 39490 36474
rect 9864 36320 9916 36372
rect 17040 36320 17092 36372
rect 35072 36320 35124 36372
rect 12532 36227 12584 36236
rect 12532 36193 12541 36227
rect 12541 36193 12575 36227
rect 12575 36193 12584 36227
rect 12532 36184 12584 36193
rect 13360 36184 13412 36236
rect 21364 36252 21416 36304
rect 24124 36116 24176 36168
rect 40776 35980 40828 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 14246 35878 14298 35930
rect 14310 35878 14362 35930
rect 14374 35878 14426 35930
rect 14438 35878 14490 35930
rect 24246 35878 24298 35930
rect 24310 35878 24362 35930
rect 24374 35878 24426 35930
rect 24438 35878 24490 35930
rect 34246 35878 34298 35930
rect 34310 35878 34362 35930
rect 34374 35878 34426 35930
rect 34438 35878 34490 35930
rect 44246 35878 44298 35930
rect 44310 35878 44362 35930
rect 44374 35878 44426 35930
rect 44438 35878 44490 35930
rect 47676 35615 47728 35624
rect 47676 35581 47685 35615
rect 47685 35581 47719 35615
rect 47719 35581 47728 35615
rect 47676 35572 47728 35581
rect 12532 35436 12584 35488
rect 21548 35436 21600 35488
rect 29000 35436 29052 35488
rect 39672 35436 39724 35488
rect 9246 35334 9298 35386
rect 9310 35334 9362 35386
rect 9374 35334 9426 35386
rect 9438 35334 9490 35386
rect 19246 35334 19298 35386
rect 19310 35334 19362 35386
rect 19374 35334 19426 35386
rect 19438 35334 19490 35386
rect 29246 35334 29298 35386
rect 29310 35334 29362 35386
rect 29374 35334 29426 35386
rect 29438 35334 29490 35386
rect 39246 35334 39298 35386
rect 39310 35334 39362 35386
rect 39374 35334 39426 35386
rect 39438 35334 39490 35386
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 14246 34790 14298 34842
rect 14310 34790 14362 34842
rect 14374 34790 14426 34842
rect 14438 34790 14490 34842
rect 24246 34790 24298 34842
rect 24310 34790 24362 34842
rect 24374 34790 24426 34842
rect 24438 34790 24490 34842
rect 34246 34790 34298 34842
rect 34310 34790 34362 34842
rect 34374 34790 34426 34842
rect 34438 34790 34490 34842
rect 44246 34790 44298 34842
rect 44310 34790 44362 34842
rect 44374 34790 44426 34842
rect 44438 34790 44490 34842
rect 39028 34484 39080 34536
rect 39672 34484 39724 34536
rect 9246 34246 9298 34298
rect 9310 34246 9362 34298
rect 9374 34246 9426 34298
rect 9438 34246 9490 34298
rect 19246 34246 19298 34298
rect 19310 34246 19362 34298
rect 19374 34246 19426 34298
rect 19438 34246 19490 34298
rect 29246 34246 29298 34298
rect 29310 34246 29362 34298
rect 29374 34246 29426 34298
rect 29438 34246 29490 34298
rect 39246 34246 39298 34298
rect 39310 34246 39362 34298
rect 39374 34246 39426 34298
rect 39438 34246 39490 34298
rect 10416 34051 10468 34060
rect 10416 34017 10425 34051
rect 10425 34017 10459 34051
rect 10459 34017 10468 34051
rect 10416 34008 10468 34017
rect 17408 33940 17460 33992
rect 38200 33847 38252 33856
rect 38200 33813 38209 33847
rect 38209 33813 38243 33847
rect 38243 33813 38252 33847
rect 38200 33804 38252 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 14246 33702 14298 33754
rect 14310 33702 14362 33754
rect 14374 33702 14426 33754
rect 14438 33702 14490 33754
rect 24246 33702 24298 33754
rect 24310 33702 24362 33754
rect 24374 33702 24426 33754
rect 24438 33702 24490 33754
rect 34246 33702 34298 33754
rect 34310 33702 34362 33754
rect 34374 33702 34426 33754
rect 34438 33702 34490 33754
rect 44246 33702 44298 33754
rect 44310 33702 44362 33754
rect 44374 33702 44426 33754
rect 44438 33702 44490 33754
rect 18328 33396 18380 33448
rect 39672 33464 39724 33516
rect 28264 33328 28316 33380
rect 38200 33328 38252 33380
rect 38292 33260 38344 33312
rect 39580 33303 39632 33312
rect 39580 33269 39589 33303
rect 39589 33269 39623 33303
rect 39623 33269 39632 33303
rect 39580 33260 39632 33269
rect 39672 33260 39724 33312
rect 47032 33303 47084 33312
rect 47032 33269 47041 33303
rect 47041 33269 47075 33303
rect 47075 33269 47084 33303
rect 47032 33260 47084 33269
rect 9246 33158 9298 33210
rect 9310 33158 9362 33210
rect 9374 33158 9426 33210
rect 9438 33158 9490 33210
rect 19246 33158 19298 33210
rect 19310 33158 19362 33210
rect 19374 33158 19426 33210
rect 19438 33158 19490 33210
rect 29246 33158 29298 33210
rect 29310 33158 29362 33210
rect 29374 33158 29426 33210
rect 29438 33158 29490 33210
rect 39246 33158 39298 33210
rect 39310 33158 39362 33210
rect 39374 33158 39426 33210
rect 39438 33158 39490 33210
rect 33140 33056 33192 33108
rect 29736 32920 29788 32972
rect 38476 32963 38528 32972
rect 38476 32929 38491 32963
rect 38491 32929 38525 32963
rect 38525 32929 38528 32963
rect 38476 32920 38528 32929
rect 47860 32963 47912 32972
rect 47860 32929 47869 32963
rect 47869 32929 47903 32963
rect 47903 32929 47912 32963
rect 47860 32920 47912 32929
rect 38016 32852 38068 32904
rect 39764 32852 39816 32904
rect 47032 32852 47084 32904
rect 42708 32784 42760 32836
rect 32404 32716 32456 32768
rect 38476 32716 38528 32768
rect 40500 32716 40552 32768
rect 46756 32716 46808 32768
rect 47584 32759 47636 32768
rect 47584 32725 47593 32759
rect 47593 32725 47627 32759
rect 47627 32725 47636 32759
rect 47584 32716 47636 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 14246 32614 14298 32666
rect 14310 32614 14362 32666
rect 14374 32614 14426 32666
rect 14438 32614 14490 32666
rect 24246 32614 24298 32666
rect 24310 32614 24362 32666
rect 24374 32614 24426 32666
rect 24438 32614 24490 32666
rect 34246 32614 34298 32666
rect 34310 32614 34362 32666
rect 34374 32614 34426 32666
rect 34438 32614 34490 32666
rect 44246 32614 44298 32666
rect 44310 32614 44362 32666
rect 44374 32614 44426 32666
rect 44438 32614 44490 32666
rect 24676 32512 24728 32564
rect 45560 32512 45612 32564
rect 47860 32512 47912 32564
rect 1768 32419 1820 32428
rect 1768 32385 1777 32419
rect 1777 32385 1811 32419
rect 1811 32385 1820 32419
rect 1768 32376 1820 32385
rect 40684 32419 40736 32428
rect 40684 32385 40693 32419
rect 40693 32385 40727 32419
rect 40727 32385 40736 32419
rect 40684 32376 40736 32385
rect 38752 32308 38804 32360
rect 37280 32172 37332 32224
rect 38016 32215 38068 32224
rect 38016 32181 38025 32215
rect 38025 32181 38059 32215
rect 38059 32181 38068 32215
rect 38016 32172 38068 32181
rect 38660 32215 38712 32224
rect 38660 32181 38669 32215
rect 38669 32181 38703 32215
rect 38703 32181 38712 32215
rect 38660 32172 38712 32181
rect 38752 32172 38804 32224
rect 39948 32172 40000 32224
rect 9246 32070 9298 32122
rect 9310 32070 9362 32122
rect 9374 32070 9426 32122
rect 9438 32070 9490 32122
rect 19246 32070 19298 32122
rect 19310 32070 19362 32122
rect 19374 32070 19426 32122
rect 19438 32070 19490 32122
rect 29246 32070 29298 32122
rect 29310 32070 29362 32122
rect 29374 32070 29426 32122
rect 29438 32070 29490 32122
rect 39246 32070 39298 32122
rect 39310 32070 39362 32122
rect 39374 32070 39426 32122
rect 39438 32070 39490 32122
rect 21548 32011 21600 32020
rect 21548 31977 21557 32011
rect 21557 31977 21591 32011
rect 21591 31977 21600 32011
rect 21548 31968 21600 31977
rect 41052 31968 41104 32020
rect 39120 31900 39172 31952
rect 38936 31875 38988 31884
rect 38936 31841 38945 31875
rect 38945 31841 38979 31875
rect 38979 31841 38988 31875
rect 38936 31832 38988 31841
rect 39856 31875 39908 31884
rect 39856 31841 39865 31875
rect 39865 31841 39899 31875
rect 39899 31841 39908 31875
rect 39856 31832 39908 31841
rect 3148 31807 3200 31816
rect 3148 31773 3157 31807
rect 3157 31773 3191 31807
rect 3191 31773 3200 31807
rect 3148 31764 3200 31773
rect 38292 31807 38344 31816
rect 38292 31773 38301 31807
rect 38301 31773 38335 31807
rect 38335 31773 38344 31807
rect 38292 31764 38344 31773
rect 39120 31807 39172 31816
rect 39120 31773 39129 31807
rect 39129 31773 39163 31807
rect 39163 31773 39172 31807
rect 39120 31764 39172 31773
rect 41236 31764 41288 31816
rect 1768 31628 1820 31680
rect 38660 31696 38712 31748
rect 39672 31696 39724 31748
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 14246 31526 14298 31578
rect 14310 31526 14362 31578
rect 14374 31526 14426 31578
rect 14438 31526 14490 31578
rect 24246 31526 24298 31578
rect 24310 31526 24362 31578
rect 24374 31526 24426 31578
rect 24438 31526 24490 31578
rect 34246 31526 34298 31578
rect 34310 31526 34362 31578
rect 34374 31526 34426 31578
rect 34438 31526 34490 31578
rect 44246 31526 44298 31578
rect 44310 31526 44362 31578
rect 44374 31526 44426 31578
rect 44438 31526 44490 31578
rect 1768 31467 1820 31476
rect 1768 31433 1777 31467
rect 1777 31433 1811 31467
rect 1811 31433 1820 31467
rect 1768 31424 1820 31433
rect 38936 31424 38988 31476
rect 3148 31356 3200 31408
rect 38384 31356 38436 31408
rect 40684 31356 40736 31408
rect 2228 31263 2280 31272
rect 2228 31229 2237 31263
rect 2237 31229 2271 31263
rect 2271 31229 2280 31263
rect 2228 31220 2280 31229
rect 4068 31220 4120 31272
rect 25688 31288 25740 31340
rect 15660 31220 15712 31272
rect 4068 31127 4120 31136
rect 4068 31093 4077 31127
rect 4077 31093 4111 31127
rect 4111 31093 4120 31127
rect 4068 31084 4120 31093
rect 39120 31152 39172 31204
rect 21916 31084 21968 31136
rect 9246 30982 9298 31034
rect 9310 30982 9362 31034
rect 9374 30982 9426 31034
rect 9438 30982 9490 31034
rect 19246 30982 19298 31034
rect 19310 30982 19362 31034
rect 19374 30982 19426 31034
rect 19438 30982 19490 31034
rect 29246 30982 29298 31034
rect 29310 30982 29362 31034
rect 29374 30982 29426 31034
rect 29438 30982 29490 31034
rect 39246 30982 39298 31034
rect 39310 30982 39362 31034
rect 39374 30982 39426 31034
rect 39438 30982 39490 31034
rect 4068 30880 4120 30932
rect 37464 30880 37516 30932
rect 15660 30855 15712 30864
rect 15660 30821 15669 30855
rect 15669 30821 15703 30855
rect 15703 30821 15712 30855
rect 15660 30812 15712 30821
rect 31852 30812 31904 30864
rect 2228 30540 2280 30592
rect 2964 30583 3016 30592
rect 2964 30549 2973 30583
rect 2973 30549 3007 30583
rect 3007 30549 3016 30583
rect 2964 30540 3016 30549
rect 47584 30744 47636 30796
rect 32404 30676 32456 30728
rect 38384 30676 38436 30728
rect 22744 30540 22796 30592
rect 33140 30540 33192 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 14246 30438 14298 30490
rect 14310 30438 14362 30490
rect 14374 30438 14426 30490
rect 14438 30438 14490 30490
rect 24246 30438 24298 30490
rect 24310 30438 24362 30490
rect 24374 30438 24426 30490
rect 24438 30438 24490 30490
rect 34246 30438 34298 30490
rect 34310 30438 34362 30490
rect 34374 30438 34426 30490
rect 34438 30438 34490 30490
rect 44246 30438 44298 30490
rect 44310 30438 44362 30490
rect 44374 30438 44426 30490
rect 44438 30438 44490 30490
rect 2964 30336 3016 30388
rect 18236 30336 18288 30388
rect 35072 30311 35124 30320
rect 35072 30277 35081 30311
rect 35081 30277 35115 30311
rect 35115 30277 35124 30311
rect 35072 30268 35124 30277
rect 35348 30311 35400 30320
rect 35348 30277 35357 30311
rect 35357 30277 35391 30311
rect 35391 30277 35400 30311
rect 35348 30268 35400 30277
rect 44088 30268 44140 30320
rect 33508 30243 33560 30252
rect 33508 30209 33517 30243
rect 33517 30209 33551 30243
rect 33551 30209 33560 30243
rect 33508 30200 33560 30209
rect 6920 29996 6972 30048
rect 31852 29996 31904 30048
rect 35624 30132 35676 30184
rect 39580 30200 39632 30252
rect 39764 30200 39816 30252
rect 43260 30200 43312 30252
rect 45008 30175 45060 30184
rect 45008 30141 45017 30175
rect 45017 30141 45051 30175
rect 45051 30141 45060 30175
rect 45008 30132 45060 30141
rect 39856 29996 39908 30048
rect 9246 29894 9298 29946
rect 9310 29894 9362 29946
rect 9374 29894 9426 29946
rect 9438 29894 9490 29946
rect 19246 29894 19298 29946
rect 19310 29894 19362 29946
rect 19374 29894 19426 29946
rect 19438 29894 19490 29946
rect 29246 29894 29298 29946
rect 29310 29894 29362 29946
rect 29374 29894 29426 29946
rect 29438 29894 29490 29946
rect 39246 29894 39298 29946
rect 39310 29894 39362 29946
rect 39374 29894 39426 29946
rect 39438 29894 39490 29946
rect 10692 29792 10744 29844
rect 33508 29792 33560 29844
rect 43996 29835 44048 29844
rect 43996 29801 44005 29835
rect 44005 29801 44039 29835
rect 44039 29801 44048 29835
rect 43996 29792 44048 29801
rect 10416 29656 10468 29708
rect 23112 29588 23164 29640
rect 25780 29631 25832 29640
rect 25780 29597 25789 29631
rect 25789 29597 25823 29631
rect 25823 29597 25832 29631
rect 25780 29588 25832 29597
rect 26056 29631 26108 29640
rect 26056 29597 26065 29631
rect 26065 29597 26099 29631
rect 26099 29597 26108 29631
rect 26056 29588 26108 29597
rect 37556 29588 37608 29640
rect 45008 29588 45060 29640
rect 42708 29520 42760 29572
rect 45192 29520 45244 29572
rect 30840 29452 30892 29504
rect 33784 29452 33836 29504
rect 35624 29452 35676 29504
rect 37280 29452 37332 29504
rect 44548 29452 44600 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 14246 29350 14298 29402
rect 14310 29350 14362 29402
rect 14374 29350 14426 29402
rect 14438 29350 14490 29402
rect 24246 29350 24298 29402
rect 24310 29350 24362 29402
rect 24374 29350 24426 29402
rect 24438 29350 24490 29402
rect 34246 29350 34298 29402
rect 34310 29350 34362 29402
rect 34374 29350 34426 29402
rect 34438 29350 34490 29402
rect 44246 29350 44298 29402
rect 44310 29350 44362 29402
rect 44374 29350 44426 29402
rect 44438 29350 44490 29402
rect 44088 29291 44140 29300
rect 44088 29257 44097 29291
rect 44097 29257 44131 29291
rect 44131 29257 44140 29291
rect 44088 29248 44140 29257
rect 43996 29180 44048 29232
rect 44088 29112 44140 29164
rect 35624 29044 35676 29096
rect 44180 29044 44232 29096
rect 44548 29044 44600 29096
rect 45192 29087 45244 29096
rect 25044 28976 25096 29028
rect 26056 28976 26108 29028
rect 30840 28976 30892 29028
rect 39580 28976 39632 29028
rect 45192 29053 45201 29087
rect 45201 29053 45235 29087
rect 45235 29053 45244 29087
rect 45192 29044 45244 29053
rect 41696 28908 41748 28960
rect 9246 28806 9298 28858
rect 9310 28806 9362 28858
rect 9374 28806 9426 28858
rect 9438 28806 9490 28858
rect 19246 28806 19298 28858
rect 19310 28806 19362 28858
rect 19374 28806 19426 28858
rect 19438 28806 19490 28858
rect 29246 28806 29298 28858
rect 29310 28806 29362 28858
rect 29374 28806 29426 28858
rect 29438 28806 29490 28858
rect 39246 28806 39298 28858
rect 39310 28806 39362 28858
rect 39374 28806 39426 28858
rect 39438 28806 39490 28858
rect 21364 28704 21416 28756
rect 22008 28704 22060 28756
rect 31852 28704 31904 28756
rect 38384 28704 38436 28756
rect 44180 28747 44232 28756
rect 44180 28713 44189 28747
rect 44189 28713 44223 28747
rect 44223 28713 44232 28747
rect 44180 28704 44232 28713
rect 23020 28568 23072 28620
rect 47032 28568 47084 28620
rect 32680 28500 32732 28552
rect 37372 28500 37424 28552
rect 38108 28543 38160 28552
rect 38108 28509 38117 28543
rect 38117 28509 38151 28543
rect 38151 28509 38160 28543
rect 38108 28500 38160 28509
rect 38384 28543 38436 28552
rect 38384 28509 38393 28543
rect 38393 28509 38427 28543
rect 38427 28509 38436 28543
rect 38384 28500 38436 28509
rect 29000 28432 29052 28484
rect 18236 28364 18288 28416
rect 24860 28364 24912 28416
rect 38016 28364 38068 28416
rect 38108 28364 38160 28416
rect 38568 28364 38620 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 14246 28262 14298 28314
rect 14310 28262 14362 28314
rect 14374 28262 14426 28314
rect 14438 28262 14490 28314
rect 24246 28262 24298 28314
rect 24310 28262 24362 28314
rect 24374 28262 24426 28314
rect 24438 28262 24490 28314
rect 34246 28262 34298 28314
rect 34310 28262 34362 28314
rect 34374 28262 34426 28314
rect 34438 28262 34490 28314
rect 44246 28262 44298 28314
rect 44310 28262 44362 28314
rect 44374 28262 44426 28314
rect 44438 28262 44490 28314
rect 22008 27956 22060 28008
rect 24124 28160 24176 28212
rect 24676 28160 24728 28212
rect 24768 28160 24820 28212
rect 32680 28160 32732 28212
rect 33232 28160 33284 28212
rect 43444 28092 43496 28144
rect 23020 27999 23072 28008
rect 23020 27965 23023 27999
rect 23023 27965 23072 27999
rect 23020 27956 23072 27965
rect 22652 27888 22704 27940
rect 24584 28024 24636 28076
rect 24860 28024 24912 28076
rect 31576 28024 31628 28076
rect 31852 28067 31904 28076
rect 31852 28033 31861 28067
rect 31861 28033 31895 28067
rect 31895 28033 31904 28067
rect 31852 28024 31904 28033
rect 31760 27999 31812 28008
rect 31760 27965 31769 27999
rect 31769 27965 31803 27999
rect 31803 27965 31812 27999
rect 33232 28024 33284 28076
rect 31760 27956 31812 27965
rect 24768 27820 24820 27872
rect 30932 27863 30984 27872
rect 30932 27829 30941 27863
rect 30941 27829 30975 27863
rect 30975 27829 30984 27863
rect 30932 27820 30984 27829
rect 31484 27863 31536 27872
rect 31484 27829 31493 27863
rect 31493 27829 31527 27863
rect 31527 27829 31536 27863
rect 31484 27820 31536 27829
rect 31576 27820 31628 27872
rect 38936 27820 38988 27872
rect 9246 27718 9298 27770
rect 9310 27718 9362 27770
rect 9374 27718 9426 27770
rect 9438 27718 9490 27770
rect 19246 27718 19298 27770
rect 19310 27718 19362 27770
rect 19374 27718 19426 27770
rect 19438 27718 19490 27770
rect 29246 27718 29298 27770
rect 29310 27718 29362 27770
rect 29374 27718 29426 27770
rect 29438 27718 29490 27770
rect 39246 27718 39298 27770
rect 39310 27718 39362 27770
rect 39374 27718 39426 27770
rect 39438 27718 39490 27770
rect 10600 27616 10652 27668
rect 30932 27616 30984 27668
rect 31852 27616 31904 27668
rect 32772 27616 32824 27668
rect 1768 27591 1820 27600
rect 1768 27557 1777 27591
rect 1777 27557 1811 27591
rect 1811 27557 1820 27591
rect 1768 27548 1820 27557
rect 4620 27548 4672 27600
rect 5172 27548 5224 27600
rect 17224 27548 17276 27600
rect 23020 27548 23072 27600
rect 28264 27480 28316 27532
rect 21916 27412 21968 27464
rect 31760 27412 31812 27464
rect 33048 27412 33100 27464
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 14246 27174 14298 27226
rect 14310 27174 14362 27226
rect 14374 27174 14426 27226
rect 14438 27174 14490 27226
rect 24246 27174 24298 27226
rect 24310 27174 24362 27226
rect 24374 27174 24426 27226
rect 24438 27174 24490 27226
rect 34246 27174 34298 27226
rect 34310 27174 34362 27226
rect 34374 27174 34426 27226
rect 34438 27174 34490 27226
rect 44246 27174 44298 27226
rect 44310 27174 44362 27226
rect 44374 27174 44426 27226
rect 44438 27174 44490 27226
rect 15936 27072 15988 27124
rect 33140 27072 33192 27124
rect 37280 27072 37332 27124
rect 33048 27004 33100 27056
rect 41604 27004 41656 27056
rect 17960 26936 18012 26988
rect 25780 26936 25832 26988
rect 2964 26868 3016 26920
rect 6736 26868 6788 26920
rect 17224 26868 17276 26920
rect 19984 26868 20036 26920
rect 30012 26911 30064 26920
rect 30012 26877 30021 26911
rect 30021 26877 30055 26911
rect 30055 26877 30064 26911
rect 30012 26868 30064 26877
rect 13636 26732 13688 26784
rect 31760 26775 31812 26784
rect 31760 26741 31769 26775
rect 31769 26741 31803 26775
rect 31803 26741 31812 26775
rect 32680 26775 32732 26784
rect 31760 26732 31812 26741
rect 32680 26741 32689 26775
rect 32689 26741 32723 26775
rect 32723 26741 32732 26775
rect 32680 26732 32732 26741
rect 37740 26732 37792 26784
rect 9246 26630 9298 26682
rect 9310 26630 9362 26682
rect 9374 26630 9426 26682
rect 9438 26630 9490 26682
rect 19246 26630 19298 26682
rect 19310 26630 19362 26682
rect 19374 26630 19426 26682
rect 19438 26630 19490 26682
rect 29246 26630 29298 26682
rect 29310 26630 29362 26682
rect 29374 26630 29426 26682
rect 29438 26630 29490 26682
rect 39246 26630 39298 26682
rect 39310 26630 39362 26682
rect 39374 26630 39426 26682
rect 39438 26630 39490 26682
rect 30012 26528 30064 26580
rect 32404 26528 32456 26580
rect 2964 26435 3016 26444
rect 2964 26401 2968 26435
rect 2968 26401 3002 26435
rect 3002 26401 3016 26435
rect 2964 26392 3016 26401
rect 2872 26256 2924 26308
rect 4620 26392 4672 26444
rect 17960 26324 18012 26376
rect 15936 26256 15988 26308
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 14246 26086 14298 26138
rect 14310 26086 14362 26138
rect 14374 26086 14426 26138
rect 14438 26086 14490 26138
rect 24246 26086 24298 26138
rect 24310 26086 24362 26138
rect 24374 26086 24426 26138
rect 24438 26086 24490 26138
rect 34246 26086 34298 26138
rect 34310 26086 34362 26138
rect 34374 26086 34426 26138
rect 34438 26086 34490 26138
rect 44246 26086 44298 26138
rect 44310 26086 44362 26138
rect 44374 26086 44426 26138
rect 44438 26086 44490 26138
rect 4620 25644 4672 25696
rect 18144 25644 18196 25696
rect 42064 25644 42116 25696
rect 45928 25687 45980 25696
rect 45928 25653 45937 25687
rect 45937 25653 45971 25687
rect 45971 25653 45980 25687
rect 45928 25644 45980 25653
rect 9246 25542 9298 25594
rect 9310 25542 9362 25594
rect 9374 25542 9426 25594
rect 9438 25542 9490 25594
rect 19246 25542 19298 25594
rect 19310 25542 19362 25594
rect 19374 25542 19426 25594
rect 19438 25542 19490 25594
rect 29246 25542 29298 25594
rect 29310 25542 29362 25594
rect 29374 25542 29426 25594
rect 29438 25542 29490 25594
rect 39246 25542 39298 25594
rect 39310 25542 39362 25594
rect 39374 25542 39426 25594
rect 39438 25542 39490 25594
rect 37372 25372 37424 25424
rect 38016 25372 38068 25424
rect 45652 25440 45704 25492
rect 46756 25440 46808 25492
rect 45928 25372 45980 25424
rect 45192 25304 45244 25356
rect 46572 25347 46624 25356
rect 46572 25313 46581 25347
rect 46581 25313 46615 25347
rect 46615 25313 46624 25347
rect 46572 25304 46624 25313
rect 46756 25347 46808 25356
rect 46756 25313 46765 25347
rect 46765 25313 46799 25347
rect 46799 25313 46808 25347
rect 46756 25304 46808 25313
rect 48136 25347 48188 25356
rect 48136 25313 48145 25347
rect 48145 25313 48179 25347
rect 48179 25313 48188 25347
rect 48136 25304 48188 25313
rect 45192 25143 45244 25152
rect 45192 25109 45201 25143
rect 45201 25109 45235 25143
rect 45235 25109 45244 25143
rect 45192 25100 45244 25109
rect 46204 25143 46256 25152
rect 46204 25109 46213 25143
rect 46213 25109 46247 25143
rect 46247 25109 46256 25143
rect 46204 25100 46256 25109
rect 47952 25143 48004 25152
rect 47952 25109 47961 25143
rect 47961 25109 47995 25143
rect 47995 25109 48004 25143
rect 47952 25100 48004 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 14246 24998 14298 25050
rect 14310 24998 14362 25050
rect 14374 24998 14426 25050
rect 14438 24998 14490 25050
rect 24246 24998 24298 25050
rect 24310 24998 24362 25050
rect 24374 24998 24426 25050
rect 24438 24998 24490 25050
rect 34246 24998 34298 25050
rect 34310 24998 34362 25050
rect 34374 24998 34426 25050
rect 34438 24998 34490 25050
rect 44246 24998 44298 25050
rect 44310 24998 44362 25050
rect 44374 24998 44426 25050
rect 44438 24998 44490 25050
rect 39764 24828 39816 24880
rect 42064 24828 42116 24880
rect 42616 24828 42668 24880
rect 38936 24760 38988 24812
rect 46572 24896 46624 24948
rect 39672 24692 39724 24744
rect 39856 24692 39908 24744
rect 45652 24692 45704 24744
rect 13728 24556 13780 24608
rect 39488 24624 39540 24676
rect 29736 24556 29788 24608
rect 9246 24454 9298 24506
rect 9310 24454 9362 24506
rect 9374 24454 9426 24506
rect 9438 24454 9490 24506
rect 19246 24454 19298 24506
rect 19310 24454 19362 24506
rect 19374 24454 19426 24506
rect 19438 24454 19490 24506
rect 29246 24454 29298 24506
rect 29310 24454 29362 24506
rect 29374 24454 29426 24506
rect 29438 24454 29490 24506
rect 39246 24454 39298 24506
rect 39310 24454 39362 24506
rect 39374 24454 39426 24506
rect 39438 24454 39490 24506
rect 19984 24352 20036 24404
rect 37556 24284 37608 24336
rect 35716 24259 35768 24268
rect 35716 24225 35725 24259
rect 35725 24225 35759 24259
rect 35759 24225 35768 24259
rect 35716 24216 35768 24225
rect 23480 24148 23532 24200
rect 17316 24012 17368 24064
rect 17500 24055 17552 24064
rect 17500 24021 17509 24055
rect 17509 24021 17543 24055
rect 17543 24021 17552 24055
rect 17500 24012 17552 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 14246 23910 14298 23962
rect 14310 23910 14362 23962
rect 14374 23910 14426 23962
rect 14438 23910 14490 23962
rect 24246 23910 24298 23962
rect 24310 23910 24362 23962
rect 24374 23910 24426 23962
rect 24438 23910 24490 23962
rect 34246 23910 34298 23962
rect 34310 23910 34362 23962
rect 34374 23910 34426 23962
rect 34438 23910 34490 23962
rect 44246 23910 44298 23962
rect 44310 23910 44362 23962
rect 44374 23910 44426 23962
rect 44438 23910 44490 23962
rect 17500 23808 17552 23860
rect 43536 23808 43588 23860
rect 31760 23740 31812 23792
rect 35716 23740 35768 23792
rect 9246 23366 9298 23418
rect 9310 23366 9362 23418
rect 9374 23366 9426 23418
rect 9438 23366 9490 23418
rect 19246 23366 19298 23418
rect 19310 23366 19362 23418
rect 19374 23366 19426 23418
rect 19438 23366 19490 23418
rect 29246 23366 29298 23418
rect 29310 23366 29362 23418
rect 29374 23366 29426 23418
rect 29438 23366 29490 23418
rect 39246 23366 39298 23418
rect 39310 23366 39362 23418
rect 39374 23366 39426 23418
rect 39438 23366 39490 23418
rect 25688 23264 25740 23316
rect 24676 23128 24728 23180
rect 39580 22924 39632 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 14246 22822 14298 22874
rect 14310 22822 14362 22874
rect 14374 22822 14426 22874
rect 14438 22822 14490 22874
rect 24246 22822 24298 22874
rect 24310 22822 24362 22874
rect 24374 22822 24426 22874
rect 24438 22822 24490 22874
rect 34246 22822 34298 22874
rect 34310 22822 34362 22874
rect 34374 22822 34426 22874
rect 34438 22822 34490 22874
rect 44246 22822 44298 22874
rect 44310 22822 44362 22874
rect 44374 22822 44426 22874
rect 44438 22822 44490 22874
rect 1768 22491 1820 22500
rect 1768 22457 1777 22491
rect 1777 22457 1811 22491
rect 1811 22457 1820 22491
rect 1768 22448 1820 22457
rect 11704 22380 11756 22432
rect 9246 22278 9298 22330
rect 9310 22278 9362 22330
rect 9374 22278 9426 22330
rect 9438 22278 9490 22330
rect 19246 22278 19298 22330
rect 19310 22278 19362 22330
rect 19374 22278 19426 22330
rect 19438 22278 19490 22330
rect 29246 22278 29298 22330
rect 29310 22278 29362 22330
rect 29374 22278 29426 22330
rect 29438 22278 29490 22330
rect 39246 22278 39298 22330
rect 39310 22278 39362 22330
rect 39374 22278 39426 22330
rect 39438 22278 39490 22330
rect 11704 22108 11756 22160
rect 12164 22108 12216 22160
rect 18420 21836 18472 21888
rect 28264 21904 28316 21956
rect 29552 21836 29604 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 14246 21734 14298 21786
rect 14310 21734 14362 21786
rect 14374 21734 14426 21786
rect 14438 21734 14490 21786
rect 24246 21734 24298 21786
rect 24310 21734 24362 21786
rect 24374 21734 24426 21786
rect 24438 21734 24490 21786
rect 34246 21734 34298 21786
rect 34310 21734 34362 21786
rect 34374 21734 34426 21786
rect 34438 21734 34490 21786
rect 44246 21734 44298 21786
rect 44310 21734 44362 21786
rect 44374 21734 44426 21786
rect 44438 21734 44490 21786
rect 9246 21190 9298 21242
rect 9310 21190 9362 21242
rect 9374 21190 9426 21242
rect 9438 21190 9490 21242
rect 19246 21190 19298 21242
rect 19310 21190 19362 21242
rect 19374 21190 19426 21242
rect 19438 21190 19490 21242
rect 29246 21190 29298 21242
rect 29310 21190 29362 21242
rect 29374 21190 29426 21242
rect 29438 21190 29490 21242
rect 39246 21190 39298 21242
rect 39310 21190 39362 21242
rect 39374 21190 39426 21242
rect 39438 21190 39490 21242
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 14246 20646 14298 20698
rect 14310 20646 14362 20698
rect 14374 20646 14426 20698
rect 14438 20646 14490 20698
rect 24246 20646 24298 20698
rect 24310 20646 24362 20698
rect 24374 20646 24426 20698
rect 24438 20646 24490 20698
rect 34246 20646 34298 20698
rect 34310 20646 34362 20698
rect 34374 20646 34426 20698
rect 34438 20646 34490 20698
rect 44246 20646 44298 20698
rect 44310 20646 44362 20698
rect 44374 20646 44426 20698
rect 44438 20646 44490 20698
rect 27252 20204 27304 20256
rect 44548 20204 44600 20256
rect 9246 20102 9298 20154
rect 9310 20102 9362 20154
rect 9374 20102 9426 20154
rect 9438 20102 9490 20154
rect 19246 20102 19298 20154
rect 19310 20102 19362 20154
rect 19374 20102 19426 20154
rect 19438 20102 19490 20154
rect 29246 20102 29298 20154
rect 29310 20102 29362 20154
rect 29374 20102 29426 20154
rect 29438 20102 29490 20154
rect 39246 20102 39298 20154
rect 39310 20102 39362 20154
rect 39374 20102 39426 20154
rect 39438 20102 39490 20154
rect 23480 20000 23532 20052
rect 27252 19975 27304 19984
rect 27252 19941 27261 19975
rect 27261 19941 27295 19975
rect 27295 19941 27304 19975
rect 27252 19932 27304 19941
rect 30840 19932 30892 19984
rect 31576 19932 31628 19984
rect 27528 19864 27580 19916
rect 29736 19907 29788 19916
rect 29736 19873 29745 19907
rect 29745 19873 29779 19907
rect 29779 19873 29788 19907
rect 29736 19864 29788 19873
rect 18144 19796 18196 19848
rect 33784 19864 33836 19916
rect 31760 19796 31812 19848
rect 27528 19660 27580 19712
rect 29552 19703 29604 19712
rect 29552 19669 29561 19703
rect 29561 19669 29595 19703
rect 29595 19669 29604 19703
rect 29552 19660 29604 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 14246 19558 14298 19610
rect 14310 19558 14362 19610
rect 14374 19558 14426 19610
rect 14438 19558 14490 19610
rect 24246 19558 24298 19610
rect 24310 19558 24362 19610
rect 24374 19558 24426 19610
rect 24438 19558 24490 19610
rect 34246 19558 34298 19610
rect 34310 19558 34362 19610
rect 34374 19558 34426 19610
rect 34438 19558 34490 19610
rect 44246 19558 44298 19610
rect 44310 19558 44362 19610
rect 44374 19558 44426 19610
rect 44438 19558 44490 19610
rect 3424 19295 3476 19304
rect 3424 19261 3433 19295
rect 3433 19261 3467 19295
rect 3467 19261 3476 19295
rect 3424 19252 3476 19261
rect 3608 19227 3660 19236
rect 3608 19193 3617 19227
rect 3617 19193 3651 19227
rect 3651 19193 3660 19227
rect 3608 19184 3660 19193
rect 13084 19252 13136 19304
rect 13360 19184 13412 19236
rect 17868 19184 17920 19236
rect 15108 19116 15160 19168
rect 9246 19014 9298 19066
rect 9310 19014 9362 19066
rect 9374 19014 9426 19066
rect 9438 19014 9490 19066
rect 39246 19014 39298 19066
rect 39310 19014 39362 19066
rect 39374 19014 39426 19066
rect 39438 19014 39490 19066
rect 3424 18572 3476 18624
rect 27528 18572 27580 18624
rect 37648 18572 37700 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 14246 18470 14298 18522
rect 14310 18470 14362 18522
rect 14374 18470 14426 18522
rect 14438 18470 14490 18522
rect 44246 18470 44298 18522
rect 44310 18470 44362 18522
rect 44374 18470 44426 18522
rect 44438 18470 44490 18522
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 9246 17926 9298 17978
rect 9310 17926 9362 17978
rect 9374 17926 9426 17978
rect 9438 17926 9490 17978
rect 39246 17926 39298 17978
rect 39310 17926 39362 17978
rect 39374 17926 39426 17978
rect 39438 17926 39490 17978
rect 12256 17867 12308 17876
rect 12256 17833 12265 17867
rect 12265 17833 12299 17867
rect 12299 17833 12308 17867
rect 12256 17824 12308 17833
rect 15108 17799 15160 17808
rect 15108 17765 15117 17799
rect 15117 17765 15151 17799
rect 15151 17765 15160 17799
rect 15108 17756 15160 17765
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 14188 17620 14240 17672
rect 1860 17527 1912 17536
rect 1860 17493 1869 17527
rect 1869 17493 1903 17527
rect 1903 17493 1912 17527
rect 1860 17484 1912 17493
rect 2596 17527 2648 17536
rect 2596 17493 2605 17527
rect 2605 17493 2639 17527
rect 2639 17493 2648 17527
rect 2596 17484 2648 17493
rect 39672 17620 39724 17672
rect 32312 17552 32364 17604
rect 32680 17552 32732 17604
rect 18052 17484 18104 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 14246 17382 14298 17434
rect 14310 17382 14362 17434
rect 14374 17382 14426 17434
rect 14438 17382 14490 17434
rect 44246 17382 44298 17434
rect 44310 17382 44362 17434
rect 44374 17382 44426 17434
rect 44438 17382 44490 17434
rect 2596 17280 2648 17332
rect 40500 17323 40552 17332
rect 40500 17289 40509 17323
rect 40509 17289 40543 17323
rect 40543 17289 40552 17323
rect 40500 17280 40552 17289
rect 18052 17212 18104 17264
rect 29552 17212 29604 17264
rect 12256 17144 12308 17196
rect 39672 17144 39724 17196
rect 13544 17008 13596 17060
rect 31484 17008 31536 17060
rect 29552 16940 29604 16992
rect 42708 17076 42760 17128
rect 41696 17008 41748 17060
rect 9246 16838 9298 16890
rect 9310 16838 9362 16890
rect 9374 16838 9426 16890
rect 9438 16838 9490 16890
rect 39246 16838 39298 16890
rect 39310 16838 39362 16890
rect 39374 16838 39426 16890
rect 39438 16838 39490 16890
rect 32312 16600 32364 16652
rect 37832 16600 37884 16652
rect 27712 16575 27764 16584
rect 27712 16541 27721 16575
rect 27721 16541 27755 16575
rect 27755 16541 27764 16575
rect 27712 16532 27764 16541
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 14246 16294 14298 16346
rect 14310 16294 14362 16346
rect 14374 16294 14426 16346
rect 14438 16294 14490 16346
rect 44246 16294 44298 16346
rect 44310 16294 44362 16346
rect 44374 16294 44426 16346
rect 44438 16294 44490 16346
rect 18144 16235 18196 16244
rect 18144 16201 18153 16235
rect 18153 16201 18187 16235
rect 18187 16201 18196 16235
rect 18144 16192 18196 16201
rect 43352 15988 43404 16040
rect 43996 15988 44048 16040
rect 17224 15852 17276 15904
rect 17868 15852 17920 15904
rect 42432 15852 42484 15904
rect 42708 15852 42760 15904
rect 9246 15750 9298 15802
rect 9310 15750 9362 15802
rect 9374 15750 9426 15802
rect 9438 15750 9490 15802
rect 39246 15750 39298 15802
rect 39310 15750 39362 15802
rect 39374 15750 39426 15802
rect 39438 15750 39490 15802
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 17960 15623 18012 15632
rect 17960 15589 17969 15623
rect 17969 15589 18003 15623
rect 18003 15589 18012 15623
rect 17960 15580 18012 15589
rect 32588 15648 32640 15700
rect 43352 15648 43404 15700
rect 17868 15555 17920 15564
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 18144 15512 18196 15564
rect 39580 15580 39632 15632
rect 47676 15512 47728 15564
rect 40776 15444 40828 15496
rect 42432 15487 42484 15496
rect 42432 15453 42441 15487
rect 42441 15453 42475 15487
rect 42475 15453 42484 15487
rect 42432 15444 42484 15453
rect 15384 15376 15436 15428
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 14246 15206 14298 15258
rect 14310 15206 14362 15258
rect 14374 15206 14426 15258
rect 14438 15206 14490 15258
rect 44246 15206 44298 15258
rect 44310 15206 44362 15258
rect 44374 15206 44426 15258
rect 44438 15206 44490 15258
rect 17960 15104 18012 15156
rect 40776 15104 40828 15156
rect 22560 15036 22612 15088
rect 14096 14832 14148 14884
rect 18144 14764 18196 14816
rect 9246 14662 9298 14714
rect 9310 14662 9362 14714
rect 9374 14662 9426 14714
rect 9438 14662 9490 14714
rect 39246 14662 39298 14714
rect 39310 14662 39362 14714
rect 39374 14662 39426 14714
rect 39438 14662 39490 14714
rect 15108 14560 15160 14612
rect 22652 14560 22704 14612
rect 17040 14424 17092 14476
rect 17684 14424 17736 14476
rect 44640 14560 44692 14612
rect 18512 14356 18564 14408
rect 13360 14220 13412 14272
rect 15384 14220 15436 14272
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 16856 14263 16908 14272
rect 16856 14229 16865 14263
rect 16865 14229 16899 14263
rect 16899 14229 16908 14263
rect 16856 14220 16908 14229
rect 24952 14220 25004 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 14246 14118 14298 14170
rect 14310 14118 14362 14170
rect 14374 14118 14426 14170
rect 14438 14118 14490 14170
rect 44246 14118 44298 14170
rect 44310 14118 44362 14170
rect 44374 14118 44426 14170
rect 44438 14118 44490 14170
rect 13084 14016 13136 14068
rect 18144 14016 18196 14068
rect 18512 14016 18564 14068
rect 14096 13991 14148 14000
rect 14096 13957 14105 13991
rect 14105 13957 14139 13991
rect 14139 13957 14148 13991
rect 14096 13948 14148 13957
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 16028 13948 16080 14000
rect 16396 13948 16448 14000
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 13360 13812 13412 13864
rect 17224 13880 17276 13932
rect 17684 13923 17736 13932
rect 17684 13889 17693 13923
rect 17693 13889 17727 13923
rect 17727 13889 17736 13923
rect 17684 13880 17736 13889
rect 42156 13880 42208 13932
rect 17776 13812 17828 13864
rect 16396 13744 16448 13796
rect 18236 13787 18288 13796
rect 18236 13753 18245 13787
rect 18245 13753 18279 13787
rect 18279 13753 18288 13787
rect 18236 13744 18288 13753
rect 9246 13574 9298 13626
rect 9310 13574 9362 13626
rect 9374 13574 9426 13626
rect 9438 13574 9490 13626
rect 39246 13574 39298 13626
rect 39310 13574 39362 13626
rect 39374 13574 39426 13626
rect 39438 13574 39490 13626
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 31668 13404 31720 13456
rect 11336 13268 11388 13320
rect 17408 13200 17460 13252
rect 38292 13200 38344 13252
rect 15108 13132 15160 13184
rect 17776 13132 17828 13184
rect 18236 13175 18288 13184
rect 18236 13141 18245 13175
rect 18245 13141 18279 13175
rect 18279 13141 18288 13175
rect 18236 13132 18288 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 14246 13030 14298 13082
rect 14310 13030 14362 13082
rect 14374 13030 14426 13082
rect 14438 13030 14490 13082
rect 44246 13030 44298 13082
rect 44310 13030 44362 13082
rect 44374 13030 44426 13082
rect 44438 13030 44490 13082
rect 39120 12928 39172 12980
rect 9246 12486 9298 12538
rect 9310 12486 9362 12538
rect 9374 12486 9426 12538
rect 9438 12486 9490 12538
rect 39246 12486 39298 12538
rect 39310 12486 39362 12538
rect 39374 12486 39426 12538
rect 39438 12486 39490 12538
rect 1860 12427 1912 12436
rect 1860 12393 1869 12427
rect 1869 12393 1903 12427
rect 1903 12393 1912 12427
rect 1860 12384 1912 12393
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 16856 12044 16908 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 14246 11942 14298 11994
rect 14310 11942 14362 11994
rect 14374 11942 14426 11994
rect 14438 11942 14490 11994
rect 44246 11942 44298 11994
rect 44310 11942 44362 11994
rect 44374 11942 44426 11994
rect 44438 11942 44490 11994
rect 12164 11840 12216 11892
rect 43444 11840 43496 11892
rect 10692 11772 10744 11824
rect 45560 11840 45612 11892
rect 12164 11636 12216 11688
rect 42432 11636 42484 11688
rect 43720 11636 43772 11688
rect 15108 11568 15160 11620
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 11336 11500 11388 11552
rect 9246 11398 9298 11450
rect 9310 11398 9362 11450
rect 9374 11398 9426 11450
rect 9438 11398 9490 11450
rect 39246 11398 39298 11450
rect 39310 11398 39362 11450
rect 39374 11398 39426 11450
rect 39438 11398 39490 11450
rect 10416 11296 10468 11348
rect 38752 11339 38804 11348
rect 37740 11228 37792 11280
rect 38752 11305 38761 11339
rect 38761 11305 38795 11339
rect 38795 11305 38804 11339
rect 38752 11296 38804 11305
rect 43720 11339 43772 11348
rect 43720 11305 43729 11339
rect 43729 11305 43763 11339
rect 43763 11305 43772 11339
rect 43720 11296 43772 11305
rect 37924 11135 37976 11144
rect 37924 11101 37933 11135
rect 37933 11101 37967 11135
rect 37967 11101 37976 11135
rect 37924 11092 37976 11101
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 14246 10854 14298 10906
rect 14310 10854 14362 10906
rect 14374 10854 14426 10906
rect 14438 10854 14490 10906
rect 44246 10854 44298 10906
rect 44310 10854 44362 10906
rect 44374 10854 44426 10906
rect 44438 10854 44490 10906
rect 37740 10752 37792 10804
rect 9246 10310 9298 10362
rect 9310 10310 9362 10362
rect 9374 10310 9426 10362
rect 9438 10310 9490 10362
rect 39246 10310 39298 10362
rect 39310 10310 39362 10362
rect 39374 10310 39426 10362
rect 39438 10310 39490 10362
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 14246 9766 14298 9818
rect 14310 9766 14362 9818
rect 14374 9766 14426 9818
rect 14438 9766 14490 9818
rect 44246 9766 44298 9818
rect 44310 9766 44362 9818
rect 44374 9766 44426 9818
rect 44438 9766 44490 9818
rect 32864 9324 32916 9376
rect 47952 9324 48004 9376
rect 9246 9222 9298 9274
rect 9310 9222 9362 9274
rect 9374 9222 9426 9274
rect 9438 9222 9490 9274
rect 24045 9215 25084 9277
rect 24045 9164 25085 9215
rect 25033 9163 25085 9164
rect 39246 9222 39298 9274
rect 39310 9222 39362 9274
rect 39374 9222 39426 9274
rect 39438 9222 39490 9274
rect 24046 9096 24098 9148
rect 24101 9096 24254 9148
rect 24257 9096 24408 9148
rect 24411 9096 24564 9148
rect 24567 9096 24720 9148
rect 24723 9096 24876 9148
rect 24879 9096 25030 9148
rect 25032 9095 25084 9147
rect 37280 9052 37332 9104
rect 45192 9052 45244 9104
rect 48136 9027 48188 9036
rect 48136 8993 48145 9027
rect 48145 8993 48179 9027
rect 48179 8993 48188 9027
rect 48136 8984 48188 8993
rect 22032 8955 22139 8956
rect 22032 8954 22251 8955
rect 22317 8954 22424 8955
rect 22032 8843 22424 8954
rect 22144 8842 22424 8843
rect 22260 8841 22312 8842
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 14246 8678 14298 8730
rect 14310 8678 14362 8730
rect 14374 8678 14426 8730
rect 14438 8678 14490 8730
rect 22033 8826 22140 8827
rect 22033 8825 22252 8826
rect 22318 8825 22425 8826
rect 22033 8664 22425 8825
rect 22145 8663 22425 8664
rect 47952 8823 48004 8832
rect 47952 8789 47961 8823
rect 47961 8789 47995 8823
rect 47995 8789 48004 8823
rect 47952 8780 48004 8789
rect 22261 8662 22313 8663
rect 44246 8678 44298 8730
rect 44310 8678 44362 8730
rect 44374 8678 44426 8730
rect 44438 8678 44490 8730
rect 22034 8647 22141 8648
rect 22262 8647 22314 8648
rect 22034 8596 22426 8647
rect 22035 8593 22426 8596
rect 22035 8481 22427 8593
rect 22147 8480 22254 8481
rect 22320 8480 22427 8481
rect 38292 8576 38344 8628
rect 38476 8576 38528 8628
rect 47952 8576 48004 8628
rect 17776 8304 17828 8356
rect 17960 8236 18012 8288
rect 18052 8236 18104 8288
rect 9246 8134 9298 8186
rect 9310 8134 9362 8186
rect 9374 8134 9426 8186
rect 9438 8134 9490 8186
rect 39246 8134 39298 8186
rect 39310 8134 39362 8186
rect 39374 8134 39426 8186
rect 39438 8134 39490 8186
rect 17408 8075 17460 8084
rect 17408 8041 17417 8075
rect 17417 8041 17451 8075
rect 17451 8041 17460 8075
rect 17408 8032 17460 8041
rect 34612 8032 34664 8084
rect 18052 7939 18104 7948
rect 18052 7905 18061 7939
rect 18061 7905 18095 7939
rect 18095 7905 18104 7939
rect 18052 7896 18104 7905
rect 37464 7964 37516 8016
rect 38108 8007 38160 8016
rect 38108 7973 38117 8007
rect 38117 7973 38151 8007
rect 38151 7973 38160 8007
rect 38108 7964 38160 7973
rect 38292 8075 38344 8084
rect 38292 8041 38301 8075
rect 38301 8041 38335 8075
rect 38335 8041 38344 8075
rect 38292 8032 38344 8041
rect 39948 8032 40000 8084
rect 42156 8075 42208 8084
rect 42156 8041 42165 8075
rect 42165 8041 42199 8075
rect 42199 8041 42208 8075
rect 42156 8032 42208 8041
rect 42616 8032 42668 8084
rect 39120 7964 39172 8016
rect 42432 7828 42484 7880
rect 11704 7760 11756 7812
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 14246 7590 14298 7642
rect 14310 7590 14362 7642
rect 14374 7590 14426 7642
rect 14438 7590 14490 7642
rect 44246 7590 44298 7642
rect 44310 7590 44362 7642
rect 44374 7590 44426 7642
rect 44438 7590 44490 7642
rect 38108 7488 38160 7540
rect 38292 7488 38344 7540
rect 1768 7463 1820 7472
rect 1768 7429 1777 7463
rect 1777 7429 1811 7463
rect 1811 7429 1820 7463
rect 1768 7420 1820 7429
rect 17868 7284 17920 7336
rect 11704 7216 11756 7268
rect 17960 7259 18012 7268
rect 17960 7225 17969 7259
rect 17969 7225 18003 7259
rect 18003 7225 18012 7259
rect 17960 7216 18012 7225
rect 21732 7216 21784 7268
rect 39028 7488 39080 7540
rect 42616 7488 42668 7540
rect 39764 7420 39816 7472
rect 42432 7463 42484 7472
rect 42432 7429 42441 7463
rect 42441 7429 42475 7463
rect 42475 7429 42484 7463
rect 42432 7420 42484 7429
rect 43260 7420 43312 7472
rect 39764 7327 39816 7336
rect 39764 7293 39773 7327
rect 39773 7293 39807 7327
rect 39807 7293 39816 7327
rect 39764 7284 39816 7293
rect 39120 7148 39172 7200
rect 39764 7148 39816 7200
rect 9246 7046 9298 7098
rect 9310 7046 9362 7098
rect 9374 7046 9426 7098
rect 9438 7046 9490 7098
rect 39246 7046 39298 7098
rect 39310 7046 39362 7098
rect 39374 7046 39426 7098
rect 39438 7046 39490 7098
rect 39120 6987 39172 6996
rect 39120 6953 39129 6987
rect 39129 6953 39163 6987
rect 39163 6953 39172 6987
rect 39120 6944 39172 6953
rect 39672 6987 39724 6996
rect 39672 6953 39681 6987
rect 39681 6953 39715 6987
rect 39715 6953 39724 6987
rect 39672 6944 39724 6953
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 18328 6604 18380 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 14246 6502 14298 6554
rect 14310 6502 14362 6554
rect 14374 6502 14426 6554
rect 14438 6502 14490 6554
rect 44246 6502 44298 6554
rect 44310 6502 44362 6554
rect 44374 6502 44426 6554
rect 44438 6502 44490 6554
rect 6920 6443 6972 6452
rect 6920 6409 6929 6443
rect 6929 6409 6963 6443
rect 6963 6409 6972 6443
rect 6920 6400 6972 6409
rect 15936 6400 15988 6452
rect 38016 6443 38068 6452
rect 38016 6409 38025 6443
rect 38025 6409 38059 6443
rect 38059 6409 38068 6443
rect 38016 6400 38068 6409
rect 17960 6060 18012 6112
rect 18328 6060 18380 6112
rect 32864 6060 32916 6112
rect 38476 6103 38528 6112
rect 38476 6069 38485 6103
rect 38485 6069 38519 6103
rect 38519 6069 38528 6103
rect 38476 6060 38528 6069
rect 9246 5958 9298 6010
rect 9310 5958 9362 6010
rect 9374 5958 9426 6010
rect 9438 5958 9490 6010
rect 39246 5958 39298 6010
rect 39310 5958 39362 6010
rect 39374 5958 39426 6010
rect 39438 5958 39490 6010
rect 18420 5856 18472 5908
rect 37648 5856 37700 5908
rect 18144 5788 18196 5840
rect 17960 5720 18012 5772
rect 18236 5720 18288 5772
rect 23940 5720 23992 5772
rect 33876 5720 33928 5772
rect 24952 5652 25004 5704
rect 17960 5627 18012 5636
rect 17960 5593 17969 5627
rect 17969 5593 18003 5627
rect 18003 5593 18012 5627
rect 17960 5584 18012 5593
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 14246 5414 14298 5466
rect 14310 5414 14362 5466
rect 14374 5414 14426 5466
rect 14438 5414 14490 5466
rect 44246 5414 44298 5466
rect 44310 5414 44362 5466
rect 44374 5414 44426 5466
rect 44438 5414 44490 5466
rect 38568 5312 38620 5364
rect 18052 5244 18104 5296
rect 23756 5244 23808 5296
rect 37280 5176 37332 5228
rect 38016 5108 38068 5160
rect 38108 5151 38160 5160
rect 38108 5117 38117 5151
rect 38117 5117 38151 5151
rect 38151 5117 38160 5151
rect 38292 5151 38344 5160
rect 38108 5108 38160 5117
rect 38292 5117 38301 5151
rect 38301 5117 38335 5151
rect 38335 5117 38344 5151
rect 38292 5108 38344 5117
rect 38844 5040 38896 5092
rect 17960 4972 18012 5024
rect 35256 4972 35308 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 9246 4870 9298 4922
rect 9310 4870 9362 4922
rect 9374 4870 9426 4922
rect 9438 4870 9490 4922
rect 39246 4870 39298 4922
rect 39310 4870 39362 4922
rect 39374 4870 39426 4922
rect 39438 4870 39490 4922
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 38108 4768 38160 4820
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 14246 4326 14298 4378
rect 14310 4326 14362 4378
rect 14374 4326 14426 4378
rect 14438 4326 14490 4378
rect 44246 4326 44298 4378
rect 44310 4326 44362 4378
rect 44374 4326 44426 4378
rect 44438 4326 44490 4378
rect 38292 4224 38344 4276
rect 43536 4131 43588 4140
rect 43536 4097 43545 4131
rect 43545 4097 43579 4131
rect 43579 4097 43588 4131
rect 43536 4088 43588 4097
rect 44640 4088 44692 4140
rect 9246 3782 9298 3834
rect 9310 3782 9362 3834
rect 9374 3782 9426 3834
rect 9438 3782 9490 3834
rect 18328 3544 18380 3596
rect 42340 3952 42392 4004
rect 39246 3782 39298 3834
rect 39310 3782 39362 3834
rect 39374 3782 39426 3834
rect 39438 3782 39490 3834
rect 41052 3723 41104 3732
rect 41052 3689 41061 3723
rect 41061 3689 41095 3723
rect 41095 3689 41104 3723
rect 41052 3680 41104 3689
rect 41604 3723 41656 3732
rect 41604 3689 41613 3723
rect 41613 3689 41647 3723
rect 41647 3689 41656 3723
rect 41604 3680 41656 3689
rect 42524 3680 42576 3732
rect 42800 3723 42852 3732
rect 42800 3689 42809 3723
rect 42809 3689 42843 3723
rect 42843 3689 42852 3723
rect 42800 3680 42852 3689
rect 43352 3723 43404 3732
rect 43352 3689 43361 3723
rect 43361 3689 43395 3723
rect 43395 3689 43404 3723
rect 43352 3680 43404 3689
rect 44548 3680 44600 3732
rect 41236 3544 41288 3596
rect 42340 3587 42392 3596
rect 42340 3553 42349 3587
rect 42349 3553 42383 3587
rect 42383 3553 42392 3587
rect 42340 3544 42392 3553
rect 42524 3587 42576 3596
rect 42524 3553 42533 3587
rect 42533 3553 42567 3587
rect 42567 3553 42576 3587
rect 42524 3544 42576 3553
rect 43536 3612 43588 3664
rect 44640 3587 44692 3596
rect 44640 3553 44649 3587
rect 44649 3553 44683 3587
rect 44683 3553 44692 3587
rect 44640 3544 44692 3553
rect 12440 3476 12492 3528
rect 13728 3476 13780 3528
rect 35256 3476 35308 3528
rect 42432 3451 42484 3460
rect 42432 3417 42441 3451
rect 42441 3417 42475 3451
rect 42475 3417 42484 3451
rect 42432 3408 42484 3417
rect 43352 3408 43404 3460
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 14246 3238 14298 3290
rect 14310 3238 14362 3290
rect 14374 3238 14426 3290
rect 14438 3238 14490 3290
rect 44246 3238 44298 3290
rect 44310 3238 44362 3290
rect 44374 3238 44426 3290
rect 44438 3238 44490 3290
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 41236 3179 41288 3188
rect 41236 3145 41245 3179
rect 41245 3145 41279 3179
rect 41279 3145 41288 3179
rect 41236 3136 41288 3145
rect 32956 3068 33008 3120
rect 42432 3068 42484 3120
rect 10876 2932 10928 2984
rect 39028 3000 39080 3052
rect 46204 3000 46256 3052
rect 43260 2932 43312 2984
rect 37924 2839 37976 2848
rect 37924 2805 37933 2839
rect 37933 2805 37967 2839
rect 37967 2805 37976 2839
rect 37924 2796 37976 2805
rect 9246 2694 9298 2746
rect 9310 2694 9362 2746
rect 9374 2694 9426 2746
rect 9438 2694 9490 2746
rect 39246 2694 39298 2746
rect 39310 2694 39362 2746
rect 39374 2694 39426 2746
rect 39438 2694 39490 2746
rect 3608 2592 3660 2644
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 37832 2592 37884 2644
rect 43260 2635 43312 2644
rect 43260 2601 43269 2635
rect 43269 2601 43303 2635
rect 43303 2601 43312 2635
rect 43260 2592 43312 2601
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 37372 2456 37424 2508
rect 37924 2499 37976 2508
rect 37924 2465 37933 2499
rect 37933 2465 37967 2499
rect 37967 2465 37976 2499
rect 37924 2456 37976 2465
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 14246 2150 14298 2202
rect 14310 2150 14362 2202
rect 14374 2150 14426 2202
rect 14438 2150 14490 2202
rect 44246 2150 44298 2202
rect 44310 2150 44362 2202
rect 44374 2150 44426 2202
rect 44438 2150 44490 2202
<< metal2 >>
rect 1858 47560 1914 47569
rect 1858 47495 1914 47504
rect 1872 47258 1900 47495
rect 9220 47356 9516 47376
rect 9276 47354 9300 47356
rect 9356 47354 9380 47356
rect 9436 47354 9460 47356
rect 9298 47302 9300 47354
rect 9362 47302 9374 47354
rect 9436 47302 9438 47354
rect 9276 47300 9300 47302
rect 9356 47300 9380 47302
rect 9436 47300 9460 47302
rect 9220 47280 9516 47300
rect 19220 47356 19516 47376
rect 19276 47354 19300 47356
rect 19356 47354 19380 47356
rect 19436 47354 19460 47356
rect 19298 47302 19300 47354
rect 19362 47302 19374 47354
rect 19436 47302 19438 47354
rect 19276 47300 19300 47302
rect 19356 47300 19380 47302
rect 19436 47300 19460 47302
rect 19220 47280 19516 47300
rect 29220 47356 29516 47376
rect 29276 47354 29300 47356
rect 29356 47354 29380 47356
rect 29436 47354 29460 47356
rect 29298 47302 29300 47354
rect 29362 47302 29374 47354
rect 29436 47302 29438 47354
rect 29276 47300 29300 47302
rect 29356 47300 29380 47302
rect 29436 47300 29460 47302
rect 29220 47280 29516 47300
rect 39220 47356 39516 47376
rect 39276 47354 39300 47356
rect 39356 47354 39380 47356
rect 39436 47354 39460 47356
rect 39298 47302 39300 47354
rect 39362 47302 39374 47354
rect 39436 47302 39438 47354
rect 39276 47300 39300 47302
rect 39356 47300 39380 47302
rect 39436 47300 39460 47302
rect 39220 47280 39516 47300
rect 1860 47252 1912 47258
rect 1860 47194 1912 47200
rect 17316 47116 17368 47122
rect 17316 47058 17368 47064
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 14220 46812 14516 46832
rect 14276 46810 14300 46812
rect 14356 46810 14380 46812
rect 14436 46810 14460 46812
rect 14298 46758 14300 46810
rect 14362 46758 14374 46810
rect 14436 46758 14438 46810
rect 14276 46756 14300 46758
rect 14356 46756 14380 46758
rect 14436 46756 14460 46758
rect 14220 46736 14516 46756
rect 9220 46268 9516 46288
rect 9276 46266 9300 46268
rect 9356 46266 9380 46268
rect 9436 46266 9460 46268
rect 9298 46214 9300 46266
rect 9362 46214 9374 46266
rect 9436 46214 9438 46266
rect 9276 46212 9300 46214
rect 9356 46212 9380 46214
rect 9436 46212 9460 46214
rect 9220 46192 9516 46212
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 14220 45724 14516 45744
rect 14276 45722 14300 45724
rect 14356 45722 14380 45724
rect 14436 45722 14460 45724
rect 14298 45670 14300 45722
rect 14362 45670 14374 45722
rect 14436 45670 14438 45722
rect 14276 45668 14300 45670
rect 14356 45668 14380 45670
rect 14436 45668 14460 45670
rect 14220 45648 14516 45668
rect 2872 45280 2924 45286
rect 2872 45222 2924 45228
rect 1860 42560 1912 42566
rect 1858 42528 1860 42537
rect 1912 42528 1914 42537
rect 1858 42463 1914 42472
rect 1858 37496 1914 37505
rect 1858 37431 1860 37440
rect 1912 37431 1914 37440
rect 1860 37402 1912 37408
rect 1766 32464 1822 32473
rect 1766 32399 1768 32408
rect 1820 32399 1822 32408
rect 1768 32370 1820 32376
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1780 31482 1808 31622
rect 1768 31476 1820 31482
rect 1768 31418 1820 31424
rect 2228 31272 2280 31278
rect 2228 31214 2280 31220
rect 2240 30598 2268 31214
rect 2228 30592 2280 30598
rect 2228 30534 2280 30540
rect 1768 27600 1820 27606
rect 1766 27568 1768 27577
rect 1820 27568 1822 27577
rect 1766 27503 1822 27512
rect 2884 26314 2912 45222
rect 9220 45180 9516 45200
rect 9276 45178 9300 45180
rect 9356 45178 9380 45180
rect 9436 45178 9460 45180
rect 9298 45126 9300 45178
rect 9362 45126 9374 45178
rect 9436 45126 9438 45178
rect 9276 45124 9300 45126
rect 9356 45124 9380 45126
rect 9436 45124 9460 45126
rect 9220 45104 9516 45124
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 14220 44636 14516 44656
rect 14276 44634 14300 44636
rect 14356 44634 14380 44636
rect 14436 44634 14460 44636
rect 14298 44582 14300 44634
rect 14362 44582 14374 44634
rect 14436 44582 14438 44634
rect 14276 44580 14300 44582
rect 14356 44580 14380 44582
rect 14436 44580 14460 44582
rect 14220 44560 14516 44580
rect 9220 44092 9516 44112
rect 9276 44090 9300 44092
rect 9356 44090 9380 44092
rect 9436 44090 9460 44092
rect 9298 44038 9300 44090
rect 9362 44038 9374 44090
rect 9436 44038 9438 44090
rect 9276 44036 9300 44038
rect 9356 44036 9380 44038
rect 9436 44036 9460 44038
rect 9220 44016 9516 44036
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 14220 43548 14516 43568
rect 14276 43546 14300 43548
rect 14356 43546 14380 43548
rect 14436 43546 14460 43548
rect 14298 43494 14300 43546
rect 14362 43494 14374 43546
rect 14436 43494 14438 43546
rect 14276 43492 14300 43494
rect 14356 43492 14380 43494
rect 14436 43492 14460 43494
rect 14220 43472 14516 43492
rect 9220 43004 9516 43024
rect 9276 43002 9300 43004
rect 9356 43002 9380 43004
rect 9436 43002 9460 43004
rect 9298 42950 9300 43002
rect 9362 42950 9374 43002
rect 9436 42950 9438 43002
rect 9276 42948 9300 42950
rect 9356 42948 9380 42950
rect 9436 42948 9460 42950
rect 9220 42928 9516 42948
rect 12256 42560 12308 42566
rect 12256 42502 12308 42508
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 9220 41916 9516 41936
rect 9276 41914 9300 41916
rect 9356 41914 9380 41916
rect 9436 41914 9460 41916
rect 9298 41862 9300 41914
rect 9362 41862 9374 41914
rect 9436 41862 9438 41914
rect 9276 41860 9300 41862
rect 9356 41860 9380 41862
rect 9436 41860 9460 41862
rect 9220 41840 9516 41860
rect 6736 41472 6788 41478
rect 6736 41414 6788 41420
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 5172 38412 5224 38418
rect 5172 38354 5224 38360
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 3160 31414 3188 31758
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 3148 31408 3200 31414
rect 3148 31350 3200 31356
rect 4068 31272 4120 31278
rect 4068 31214 4120 31220
rect 4080 31142 4108 31214
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30938 4108 31078
rect 4068 30932 4120 30938
rect 4068 30874 4120 30880
rect 2964 30592 3016 30598
rect 2964 30534 3016 30540
rect 2976 30394 3004 30534
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 2964 30388 3016 30394
rect 2964 30330 3016 30336
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 5184 27606 5212 38354
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 2964 26920 3016 26926
rect 2964 26862 3016 26868
rect 2976 26450 3004 26862
rect 4632 26450 4660 27542
rect 6748 26926 6776 41414
rect 9220 40828 9516 40848
rect 9276 40826 9300 40828
rect 9356 40826 9380 40828
rect 9436 40826 9460 40828
rect 9298 40774 9300 40826
rect 9362 40774 9374 40826
rect 9436 40774 9438 40826
rect 9276 40772 9300 40774
rect 9356 40772 9380 40774
rect 9436 40772 9460 40774
rect 9220 40752 9516 40772
rect 9220 39740 9516 39760
rect 9276 39738 9300 39740
rect 9356 39738 9380 39740
rect 9436 39738 9460 39740
rect 9298 39686 9300 39738
rect 9362 39686 9374 39738
rect 9436 39686 9438 39738
rect 9276 39684 9300 39686
rect 9356 39684 9380 39686
rect 9436 39684 9460 39686
rect 9220 39664 9516 39684
rect 9220 38652 9516 38672
rect 9276 38650 9300 38652
rect 9356 38650 9380 38652
rect 9436 38650 9460 38652
rect 9298 38598 9300 38650
rect 9362 38598 9374 38650
rect 9436 38598 9438 38650
rect 9276 38596 9300 38598
rect 9356 38596 9380 38598
rect 9436 38596 9460 38598
rect 9220 38576 9516 38596
rect 9864 38344 9916 38350
rect 9864 38286 9916 38292
rect 9220 37564 9516 37584
rect 9276 37562 9300 37564
rect 9356 37562 9380 37564
rect 9436 37562 9460 37564
rect 9298 37510 9300 37562
rect 9362 37510 9374 37562
rect 9436 37510 9438 37562
rect 9276 37508 9300 37510
rect 9356 37508 9380 37510
rect 9436 37508 9460 37510
rect 9220 37488 9516 37508
rect 9220 36476 9516 36496
rect 9276 36474 9300 36476
rect 9356 36474 9380 36476
rect 9436 36474 9460 36476
rect 9298 36422 9300 36474
rect 9362 36422 9374 36474
rect 9436 36422 9438 36474
rect 9276 36420 9300 36422
rect 9356 36420 9380 36422
rect 9436 36420 9460 36422
rect 9220 36400 9516 36420
rect 9876 36378 9904 38286
rect 11704 36848 11756 36854
rect 11704 36790 11756 36796
rect 9864 36372 9916 36378
rect 9864 36314 9916 36320
rect 9220 35388 9516 35408
rect 9276 35386 9300 35388
rect 9356 35386 9380 35388
rect 9436 35386 9460 35388
rect 9298 35334 9300 35386
rect 9362 35334 9374 35386
rect 9436 35334 9438 35386
rect 9276 35332 9300 35334
rect 9356 35332 9380 35334
rect 9436 35332 9460 35334
rect 9220 35312 9516 35332
rect 9220 34300 9516 34320
rect 9276 34298 9300 34300
rect 9356 34298 9380 34300
rect 9436 34298 9460 34300
rect 9298 34246 9300 34298
rect 9362 34246 9374 34298
rect 9436 34246 9438 34298
rect 9276 34244 9300 34246
rect 9356 34244 9380 34246
rect 9436 34244 9460 34246
rect 9220 34224 9516 34244
rect 10416 34060 10468 34066
rect 10416 34002 10468 34008
rect 9220 33212 9516 33232
rect 9276 33210 9300 33212
rect 9356 33210 9380 33212
rect 9436 33210 9460 33212
rect 9298 33158 9300 33210
rect 9362 33158 9374 33210
rect 9436 33158 9438 33210
rect 9276 33156 9300 33158
rect 9356 33156 9380 33158
rect 9436 33156 9460 33158
rect 9220 33136 9516 33156
rect 9220 32124 9516 32144
rect 9276 32122 9300 32124
rect 9356 32122 9380 32124
rect 9436 32122 9460 32124
rect 9298 32070 9300 32122
rect 9362 32070 9374 32122
rect 9436 32070 9438 32122
rect 9276 32068 9300 32070
rect 9356 32068 9380 32070
rect 9436 32068 9460 32070
rect 9220 32048 9516 32068
rect 9220 31036 9516 31056
rect 9276 31034 9300 31036
rect 9356 31034 9380 31036
rect 9436 31034 9460 31036
rect 9298 30982 9300 31034
rect 9362 30982 9374 31034
rect 9436 30982 9438 31034
rect 9276 30980 9300 30982
rect 9356 30980 9380 30982
rect 9436 30980 9460 30982
rect 9220 30960 9516 30980
rect 6920 30048 6972 30054
rect 6920 29990 6972 29996
rect 6736 26920 6788 26926
rect 6736 26862 6788 26868
rect 2964 26444 3016 26450
rect 2964 26386 3016 26392
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 2872 26308 2924 26314
rect 2872 26250 2924 26256
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4632 25702 4660 26386
rect 4620 25696 4672 25702
rect 4620 25638 4672 25644
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 1766 22536 1822 22545
rect 1766 22471 1768 22480
rect 1820 22471 1822 22480
rect 1768 22442 1820 22448
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3436 18630 3464 19246
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 1860 17536 1912 17542
rect 1858 17504 1860 17513
rect 2596 17536 2648 17542
rect 1912 17504 1914 17513
rect 2596 17478 2648 17484
rect 1858 17439 1914 17448
rect 2608 17338 2636 17478
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 1858 12472 1914 12481
rect 1858 12407 1860 12416
rect 1912 12407 1914 12416
rect 1860 12378 1912 12384
rect 1768 7472 1820 7478
rect 1766 7440 1768 7449
rect 1820 7440 1822 7449
rect 1766 7375 1822 7384
rect 3620 2650 3648 19178
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 6932 6458 6960 29990
rect 9220 29948 9516 29968
rect 9276 29946 9300 29948
rect 9356 29946 9380 29948
rect 9436 29946 9460 29948
rect 9298 29894 9300 29946
rect 9362 29894 9374 29946
rect 9436 29894 9438 29946
rect 9276 29892 9300 29894
rect 9356 29892 9380 29894
rect 9436 29892 9460 29894
rect 9220 29872 9516 29892
rect 10428 29714 10456 34002
rect 10692 29844 10744 29850
rect 10692 29786 10744 29792
rect 10416 29708 10468 29714
rect 10416 29650 10468 29656
rect 9220 28860 9516 28880
rect 9276 28858 9300 28860
rect 9356 28858 9380 28860
rect 9436 28858 9460 28860
rect 9298 28806 9300 28858
rect 9362 28806 9374 28858
rect 9436 28806 9438 28858
rect 9276 28804 9300 28806
rect 9356 28804 9380 28806
rect 9436 28804 9460 28806
rect 9220 28784 9516 28804
rect 9220 27772 9516 27792
rect 9276 27770 9300 27772
rect 9356 27770 9380 27772
rect 9436 27770 9460 27772
rect 9298 27718 9300 27770
rect 9362 27718 9374 27770
rect 9436 27718 9438 27770
rect 9276 27716 9300 27718
rect 9356 27716 9380 27718
rect 9436 27716 9460 27718
rect 9220 27696 9516 27716
rect 9220 26684 9516 26704
rect 9276 26682 9300 26684
rect 9356 26682 9380 26684
rect 9436 26682 9460 26684
rect 9298 26630 9300 26682
rect 9362 26630 9374 26682
rect 9436 26630 9438 26682
rect 9276 26628 9300 26630
rect 9356 26628 9380 26630
rect 9436 26628 9460 26630
rect 9220 26608 9516 26628
rect 9220 25596 9516 25616
rect 9276 25594 9300 25596
rect 9356 25594 9380 25596
rect 9436 25594 9460 25596
rect 9298 25542 9300 25594
rect 9362 25542 9374 25594
rect 9436 25542 9438 25594
rect 9276 25540 9300 25542
rect 9356 25540 9380 25542
rect 9436 25540 9460 25542
rect 9220 25520 9516 25540
rect 9220 24508 9516 24528
rect 9276 24506 9300 24508
rect 9356 24506 9380 24508
rect 9436 24506 9460 24508
rect 9298 24454 9300 24506
rect 9362 24454 9374 24506
rect 9436 24454 9438 24506
rect 9276 24452 9300 24454
rect 9356 24452 9380 24454
rect 9436 24452 9460 24454
rect 9220 24432 9516 24452
rect 9220 23420 9516 23440
rect 9276 23418 9300 23420
rect 9356 23418 9380 23420
rect 9436 23418 9460 23420
rect 9298 23366 9300 23418
rect 9362 23366 9374 23418
rect 9436 23366 9438 23418
rect 9276 23364 9300 23366
rect 9356 23364 9380 23366
rect 9436 23364 9460 23366
rect 9220 23344 9516 23364
rect 9220 22332 9516 22352
rect 9276 22330 9300 22332
rect 9356 22330 9380 22332
rect 9436 22330 9460 22332
rect 9298 22278 9300 22330
rect 9362 22278 9374 22330
rect 9436 22278 9438 22330
rect 9276 22276 9300 22278
rect 9356 22276 9380 22278
rect 9436 22276 9460 22278
rect 9220 22256 9516 22276
rect 9220 21244 9516 21264
rect 9276 21242 9300 21244
rect 9356 21242 9380 21244
rect 9436 21242 9460 21244
rect 9298 21190 9300 21242
rect 9362 21190 9374 21242
rect 9436 21190 9438 21242
rect 9276 21188 9300 21190
rect 9356 21188 9380 21190
rect 9436 21188 9460 21190
rect 9220 21168 9516 21188
rect 9220 20156 9516 20176
rect 9276 20154 9300 20156
rect 9356 20154 9380 20156
rect 9436 20154 9460 20156
rect 9298 20102 9300 20154
rect 9362 20102 9374 20154
rect 9436 20102 9438 20154
rect 9276 20100 9300 20102
rect 9356 20100 9380 20102
rect 9436 20100 9460 20102
rect 9220 20080 9516 20100
rect 9220 19068 9516 19088
rect 9276 19066 9300 19068
rect 9356 19066 9380 19068
rect 9436 19066 9460 19068
rect 9298 19014 9300 19066
rect 9362 19014 9374 19066
rect 9436 19014 9438 19066
rect 9276 19012 9300 19014
rect 9356 19012 9380 19014
rect 9436 19012 9460 19014
rect 9220 18992 9516 19012
rect 9220 17980 9516 18000
rect 9276 17978 9300 17980
rect 9356 17978 9380 17980
rect 9436 17978 9460 17980
rect 9298 17926 9300 17978
rect 9362 17926 9374 17978
rect 9436 17926 9438 17978
rect 9276 17924 9300 17926
rect 9356 17924 9380 17926
rect 9436 17924 9460 17926
rect 9220 17904 9516 17924
rect 9220 16892 9516 16912
rect 9276 16890 9300 16892
rect 9356 16890 9380 16892
rect 9436 16890 9460 16892
rect 9298 16838 9300 16890
rect 9362 16838 9374 16890
rect 9436 16838 9438 16890
rect 9276 16836 9300 16838
rect 9356 16836 9380 16838
rect 9436 16836 9460 16838
rect 9220 16816 9516 16836
rect 9220 15804 9516 15824
rect 9276 15802 9300 15804
rect 9356 15802 9380 15804
rect 9436 15802 9460 15804
rect 9298 15750 9300 15802
rect 9362 15750 9374 15802
rect 9436 15750 9438 15802
rect 9276 15748 9300 15750
rect 9356 15748 9380 15750
rect 9436 15748 9460 15750
rect 9220 15728 9516 15748
rect 9220 14716 9516 14736
rect 9276 14714 9300 14716
rect 9356 14714 9380 14716
rect 9436 14714 9460 14716
rect 9298 14662 9300 14714
rect 9362 14662 9374 14714
rect 9436 14662 9438 14714
rect 9276 14660 9300 14662
rect 9356 14660 9380 14662
rect 9436 14660 9460 14662
rect 9220 14640 9516 14660
rect 9220 13628 9516 13648
rect 9276 13626 9300 13628
rect 9356 13626 9380 13628
rect 9436 13626 9460 13628
rect 9298 13574 9300 13626
rect 9362 13574 9374 13626
rect 9436 13574 9438 13626
rect 9276 13572 9300 13574
rect 9356 13572 9380 13574
rect 9436 13572 9460 13574
rect 9220 13552 9516 13572
rect 9220 12540 9516 12560
rect 9276 12538 9300 12540
rect 9356 12538 9380 12540
rect 9436 12538 9460 12540
rect 9298 12486 9300 12538
rect 9362 12486 9374 12538
rect 9436 12486 9438 12538
rect 9276 12484 9300 12486
rect 9356 12484 9380 12486
rect 9436 12484 9460 12486
rect 9220 12464 9516 12484
rect 10428 11558 10456 29650
rect 10600 27668 10652 27674
rect 10600 27610 10652 27616
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 9220 11452 9516 11472
rect 9276 11450 9300 11452
rect 9356 11450 9380 11452
rect 9436 11450 9460 11452
rect 9298 11398 9300 11450
rect 9362 11398 9374 11450
rect 9436 11398 9438 11450
rect 9276 11396 9300 11398
rect 9356 11396 9380 11398
rect 9436 11396 9460 11398
rect 9220 11376 9516 11396
rect 10428 11354 10456 11494
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 9220 10364 9516 10384
rect 9276 10362 9300 10364
rect 9356 10362 9380 10364
rect 9436 10362 9460 10364
rect 9298 10310 9300 10362
rect 9362 10310 9374 10362
rect 9436 10310 9438 10362
rect 9276 10308 9300 10310
rect 9356 10308 9380 10310
rect 9436 10308 9460 10310
rect 9220 10288 9516 10308
rect 9220 9276 9516 9296
rect 9276 9274 9300 9276
rect 9356 9274 9380 9276
rect 9436 9274 9460 9276
rect 9298 9222 9300 9274
rect 9362 9222 9374 9274
rect 9436 9222 9438 9274
rect 9276 9220 9300 9222
rect 9356 9220 9380 9222
rect 9436 9220 9460 9222
rect 9220 9200 9516 9220
rect 9220 8188 9516 8208
rect 9276 8186 9300 8188
rect 9356 8186 9380 8188
rect 9436 8186 9460 8188
rect 9298 8134 9300 8186
rect 9362 8134 9374 8186
rect 9436 8134 9438 8186
rect 9276 8132 9300 8134
rect 9356 8132 9380 8134
rect 9436 8132 9460 8134
rect 9220 8112 9516 8132
rect 9220 7100 9516 7120
rect 9276 7098 9300 7100
rect 9356 7098 9380 7100
rect 9436 7098 9460 7100
rect 9298 7046 9300 7098
rect 9362 7046 9374 7098
rect 9436 7046 9438 7098
rect 9276 7044 9300 7046
rect 9356 7044 9380 7046
rect 9436 7044 9460 7046
rect 9220 7024 9516 7044
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 9220 6012 9516 6032
rect 9276 6010 9300 6012
rect 9356 6010 9380 6012
rect 9436 6010 9460 6012
rect 9298 5958 9300 6010
rect 9362 5958 9374 6010
rect 9436 5958 9438 6010
rect 9276 5956 9300 5958
rect 9356 5956 9380 5958
rect 9436 5956 9460 5958
rect 9220 5936 9516 5956
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 9220 4924 9516 4944
rect 9276 4922 9300 4924
rect 9356 4922 9380 4924
rect 9436 4922 9460 4924
rect 9298 4870 9300 4922
rect 9362 4870 9374 4922
rect 9436 4870 9438 4922
rect 9276 4868 9300 4870
rect 9356 4868 9380 4870
rect 9436 4868 9460 4870
rect 9220 4848 9516 4868
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 9220 3836 9516 3856
rect 9276 3834 9300 3836
rect 9356 3834 9380 3836
rect 9436 3834 9460 3836
rect 9298 3782 9300 3834
rect 9362 3782 9374 3834
rect 9436 3782 9438 3834
rect 9276 3780 9300 3782
rect 9356 3780 9380 3782
rect 9436 3780 9460 3782
rect 9220 3760 9516 3780
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 10612 3194 10640 27610
rect 10704 11830 10732 29786
rect 11716 22438 11744 36790
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11716 22166 11744 22374
rect 11704 22160 11756 22166
rect 11704 22102 11756 22108
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11348 12442 11376 13262
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 11348 11558 11376 12378
rect 12176 11898 12204 22102
rect 12268 17882 12296 42502
rect 14220 42460 14516 42480
rect 14276 42458 14300 42460
rect 14356 42458 14380 42460
rect 14436 42458 14460 42460
rect 14298 42406 14300 42458
rect 14362 42406 14374 42458
rect 14436 42406 14438 42458
rect 14276 42404 14300 42406
rect 14356 42404 14380 42406
rect 14436 42404 14460 42406
rect 14220 42384 14516 42404
rect 13084 41676 13136 41682
rect 13084 41618 13136 41624
rect 13096 40934 13124 41618
rect 13636 41608 13688 41614
rect 13636 41550 13688 41556
rect 13084 40928 13136 40934
rect 13084 40870 13136 40876
rect 12532 36236 12584 36242
rect 12532 36178 12584 36184
rect 12544 35494 12572 36178
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 13096 19310 13124 40870
rect 13360 36576 13412 36582
rect 13360 36518 13412 36524
rect 13372 36242 13400 36518
rect 13360 36236 13412 36242
rect 13360 36178 13412 36184
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12268 17202 12296 17818
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 13096 14074 13124 19246
rect 13372 19242 13400 36178
rect 13648 26790 13676 41550
rect 15108 41540 15160 41546
rect 15108 41482 15160 41488
rect 14220 41372 14516 41392
rect 14276 41370 14300 41372
rect 14356 41370 14380 41372
rect 14436 41370 14460 41372
rect 14298 41318 14300 41370
rect 14362 41318 14374 41370
rect 14436 41318 14438 41370
rect 14276 41316 14300 41318
rect 14356 41316 14380 41318
rect 14436 41316 14460 41318
rect 14220 41296 14516 41316
rect 14220 40284 14516 40304
rect 14276 40282 14300 40284
rect 14356 40282 14380 40284
rect 14436 40282 14460 40284
rect 14298 40230 14300 40282
rect 14362 40230 14374 40282
rect 14436 40230 14438 40282
rect 14276 40228 14300 40230
rect 14356 40228 14380 40230
rect 14436 40228 14460 40230
rect 14220 40208 14516 40228
rect 15120 39574 15148 41482
rect 15108 39568 15160 39574
rect 15108 39510 15160 39516
rect 14220 39196 14516 39216
rect 14276 39194 14300 39196
rect 14356 39194 14380 39196
rect 14436 39194 14460 39196
rect 14298 39142 14300 39194
rect 14362 39142 14374 39194
rect 14436 39142 14438 39194
rect 14276 39140 14300 39142
rect 14356 39140 14380 39142
rect 14436 39140 14460 39142
rect 14220 39120 14516 39140
rect 16948 38480 17000 38486
rect 16948 38422 17000 38428
rect 14220 38108 14516 38128
rect 14276 38106 14300 38108
rect 14356 38106 14380 38108
rect 14436 38106 14460 38108
rect 14298 38054 14300 38106
rect 14362 38054 14374 38106
rect 14436 38054 14438 38106
rect 14276 38052 14300 38054
rect 14356 38052 14380 38054
rect 14436 38052 14460 38054
rect 14220 38032 14516 38052
rect 14220 37020 14516 37040
rect 14276 37018 14300 37020
rect 14356 37018 14380 37020
rect 14436 37018 14460 37020
rect 14298 36966 14300 37018
rect 14362 36966 14374 37018
rect 14436 36966 14438 37018
rect 14276 36964 14300 36966
rect 14356 36964 14380 36966
rect 14436 36964 14460 36966
rect 14220 36944 14516 36964
rect 14220 35932 14516 35952
rect 14276 35930 14300 35932
rect 14356 35930 14380 35932
rect 14436 35930 14460 35932
rect 14298 35878 14300 35930
rect 14362 35878 14374 35930
rect 14436 35878 14438 35930
rect 14276 35876 14300 35878
rect 14356 35876 14380 35878
rect 14436 35876 14460 35878
rect 14220 35856 14516 35876
rect 16960 35894 16988 38422
rect 17040 36576 17092 36582
rect 17040 36518 17092 36524
rect 17052 36378 17080 36518
rect 17040 36372 17092 36378
rect 17040 36314 17092 36320
rect 16960 35866 17080 35894
rect 14220 34844 14516 34864
rect 14276 34842 14300 34844
rect 14356 34842 14380 34844
rect 14436 34842 14460 34844
rect 14298 34790 14300 34842
rect 14362 34790 14374 34842
rect 14436 34790 14438 34842
rect 14276 34788 14300 34790
rect 14356 34788 14380 34790
rect 14436 34788 14460 34790
rect 14220 34768 14516 34788
rect 14220 33756 14516 33776
rect 14276 33754 14300 33756
rect 14356 33754 14380 33756
rect 14436 33754 14460 33756
rect 14298 33702 14300 33754
rect 14362 33702 14374 33754
rect 14436 33702 14438 33754
rect 14276 33700 14300 33702
rect 14356 33700 14380 33702
rect 14436 33700 14460 33702
rect 14220 33680 14516 33700
rect 14220 32668 14516 32688
rect 14276 32666 14300 32668
rect 14356 32666 14380 32668
rect 14436 32666 14460 32668
rect 14298 32614 14300 32666
rect 14362 32614 14374 32666
rect 14436 32614 14438 32666
rect 14276 32612 14300 32614
rect 14356 32612 14380 32614
rect 14436 32612 14460 32614
rect 14220 32592 14516 32612
rect 14220 31580 14516 31600
rect 14276 31578 14300 31580
rect 14356 31578 14380 31580
rect 14436 31578 14460 31580
rect 14298 31526 14300 31578
rect 14362 31526 14374 31578
rect 14436 31526 14438 31578
rect 14276 31524 14300 31526
rect 14356 31524 14380 31526
rect 14436 31524 14460 31526
rect 14220 31504 14516 31524
rect 15660 31272 15712 31278
rect 15660 31214 15712 31220
rect 15672 30870 15700 31214
rect 15660 30864 15712 30870
rect 15660 30806 15712 30812
rect 14220 30492 14516 30512
rect 14276 30490 14300 30492
rect 14356 30490 14380 30492
rect 14436 30490 14460 30492
rect 14298 30438 14300 30490
rect 14362 30438 14374 30490
rect 14436 30438 14438 30490
rect 14276 30436 14300 30438
rect 14356 30436 14380 30438
rect 14436 30436 14460 30438
rect 14220 30416 14516 30436
rect 14220 29404 14516 29424
rect 14276 29402 14300 29404
rect 14356 29402 14380 29404
rect 14436 29402 14460 29404
rect 14298 29350 14300 29402
rect 14362 29350 14374 29402
rect 14436 29350 14438 29402
rect 14276 29348 14300 29350
rect 14356 29348 14380 29350
rect 14436 29348 14460 29350
rect 14220 29328 14516 29348
rect 14220 28316 14516 28336
rect 14276 28314 14300 28316
rect 14356 28314 14380 28316
rect 14436 28314 14460 28316
rect 14298 28262 14300 28314
rect 14362 28262 14374 28314
rect 14436 28262 14438 28314
rect 14276 28260 14300 28262
rect 14356 28260 14380 28262
rect 14436 28260 14460 28262
rect 14220 28240 14516 28260
rect 14220 27228 14516 27248
rect 14276 27226 14300 27228
rect 14356 27226 14380 27228
rect 14436 27226 14460 27228
rect 14298 27174 14300 27226
rect 14362 27174 14374 27226
rect 14436 27174 14438 27226
rect 14276 27172 14300 27174
rect 14356 27172 14380 27174
rect 14436 27172 14460 27174
rect 14220 27152 14516 27172
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 15948 26314 15976 27066
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 14220 26140 14516 26160
rect 14276 26138 14300 26140
rect 14356 26138 14380 26140
rect 14436 26138 14460 26140
rect 14298 26086 14300 26138
rect 14362 26086 14374 26138
rect 14436 26086 14438 26138
rect 14276 26084 14300 26086
rect 14356 26084 14380 26086
rect 14436 26084 14460 26086
rect 14220 26064 14516 26084
rect 14220 25052 14516 25072
rect 14276 25050 14300 25052
rect 14356 25050 14380 25052
rect 14436 25050 14460 25052
rect 14298 24998 14300 25050
rect 14362 24998 14374 25050
rect 14436 24998 14438 25050
rect 14276 24996 14300 24998
rect 14356 24996 14380 24998
rect 14436 24996 14460 24998
rect 14220 24976 14516 24996
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13556 17066 13584 17614
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13372 13870 13400 14214
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12176 11694 12204 11834
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11716 7274 11744 7754
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 13740 3534 13768 24550
rect 14220 23964 14516 23984
rect 14276 23962 14300 23964
rect 14356 23962 14380 23964
rect 14436 23962 14460 23964
rect 14298 23910 14300 23962
rect 14362 23910 14374 23962
rect 14436 23910 14438 23962
rect 14276 23908 14300 23910
rect 14356 23908 14380 23910
rect 14436 23908 14460 23910
rect 14220 23888 14516 23908
rect 14220 22876 14516 22896
rect 14276 22874 14300 22876
rect 14356 22874 14380 22876
rect 14436 22874 14460 22876
rect 14298 22822 14300 22874
rect 14362 22822 14374 22874
rect 14436 22822 14438 22874
rect 14276 22820 14300 22822
rect 14356 22820 14380 22822
rect 14436 22820 14460 22822
rect 14220 22800 14516 22820
rect 14220 21788 14516 21808
rect 14276 21786 14300 21788
rect 14356 21786 14380 21788
rect 14436 21786 14460 21788
rect 14298 21734 14300 21786
rect 14362 21734 14374 21786
rect 14436 21734 14438 21786
rect 14276 21732 14300 21734
rect 14356 21732 14380 21734
rect 14436 21732 14460 21734
rect 14220 21712 14516 21732
rect 14220 20700 14516 20720
rect 14276 20698 14300 20700
rect 14356 20698 14380 20700
rect 14436 20698 14460 20700
rect 14298 20646 14300 20698
rect 14362 20646 14374 20698
rect 14436 20646 14438 20698
rect 14276 20644 14300 20646
rect 14356 20644 14380 20646
rect 14436 20644 14460 20646
rect 14220 20624 14516 20644
rect 14220 19612 14516 19632
rect 14276 19610 14300 19612
rect 14356 19610 14380 19612
rect 14436 19610 14460 19612
rect 14298 19558 14300 19610
rect 14362 19558 14374 19610
rect 14436 19558 14438 19610
rect 14276 19556 14300 19558
rect 14356 19556 14380 19558
rect 14436 19556 14460 19558
rect 14220 19536 14516 19556
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 14220 18524 14516 18544
rect 14276 18522 14300 18524
rect 14356 18522 14380 18524
rect 14436 18522 14460 18524
rect 14298 18470 14300 18522
rect 14362 18470 14374 18522
rect 14436 18470 14438 18522
rect 14276 18468 14300 18470
rect 14356 18468 14380 18470
rect 14436 18468 14460 18470
rect 14220 18448 14516 18468
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17678 14228 18022
rect 15120 17814 15148 19110
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14220 17436 14516 17456
rect 14276 17434 14300 17436
rect 14356 17434 14380 17436
rect 14436 17434 14460 17436
rect 14298 17382 14300 17434
rect 14362 17382 14374 17434
rect 14436 17382 14438 17434
rect 14276 17380 14300 17382
rect 14356 17380 14380 17382
rect 14436 17380 14460 17382
rect 14220 17360 14516 17380
rect 14220 16348 14516 16368
rect 14276 16346 14300 16348
rect 14356 16346 14380 16348
rect 14436 16346 14460 16348
rect 14298 16294 14300 16346
rect 14362 16294 14374 16346
rect 14436 16294 14438 16346
rect 14276 16292 14300 16294
rect 14356 16292 14380 16294
rect 14436 16292 14460 16294
rect 14220 16272 14516 16292
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 14220 15260 14516 15280
rect 14276 15258 14300 15260
rect 14356 15258 14380 15260
rect 14436 15258 14460 15260
rect 14298 15206 14300 15258
rect 14362 15206 14374 15258
rect 14436 15206 14438 15258
rect 14276 15204 14300 15206
rect 14356 15204 14380 15206
rect 14436 15204 14460 15206
rect 14220 15184 14516 15204
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14006 14136 14826
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 14220 14172 14516 14192
rect 14276 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14298 14118 14300 14170
rect 14362 14118 14374 14170
rect 14436 14118 14438 14170
rect 14276 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14220 14096 14516 14116
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 15120 13938 15148 14554
rect 15396 14278 15424 15370
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15948 13938 15976 26250
rect 17052 14482 17080 35866
rect 17224 27600 17276 27606
rect 17224 27542 17276 27548
rect 17236 26926 17264 27542
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17236 15910 17264 26862
rect 17328 24070 17356 47058
rect 24220 46812 24516 46832
rect 24276 46810 24300 46812
rect 24356 46810 24380 46812
rect 24436 46810 24460 46812
rect 24298 46758 24300 46810
rect 24362 46758 24374 46810
rect 24436 46758 24438 46810
rect 24276 46756 24300 46758
rect 24356 46756 24380 46758
rect 24436 46756 24460 46758
rect 24220 46736 24516 46756
rect 34220 46812 34516 46832
rect 34276 46810 34300 46812
rect 34356 46810 34380 46812
rect 34436 46810 34460 46812
rect 34298 46758 34300 46810
rect 34362 46758 34374 46810
rect 34436 46758 34438 46810
rect 34276 46756 34300 46758
rect 34356 46756 34380 46758
rect 34436 46756 34460 46758
rect 34220 46736 34516 46756
rect 44220 46812 44516 46832
rect 44276 46810 44300 46812
rect 44356 46810 44380 46812
rect 44436 46810 44460 46812
rect 44298 46758 44300 46810
rect 44362 46758 44374 46810
rect 44436 46758 44438 46810
rect 44276 46756 44300 46758
rect 44356 46756 44380 46758
rect 44436 46756 44460 46758
rect 44220 46736 44516 46756
rect 19220 46268 19516 46288
rect 19276 46266 19300 46268
rect 19356 46266 19380 46268
rect 19436 46266 19460 46268
rect 19298 46214 19300 46266
rect 19362 46214 19374 46266
rect 19436 46214 19438 46266
rect 19276 46212 19300 46214
rect 19356 46212 19380 46214
rect 19436 46212 19460 46214
rect 19220 46192 19516 46212
rect 29220 46268 29516 46288
rect 29276 46266 29300 46268
rect 29356 46266 29380 46268
rect 29436 46266 29460 46268
rect 29298 46214 29300 46266
rect 29362 46214 29374 46266
rect 29436 46214 29438 46266
rect 29276 46212 29300 46214
rect 29356 46212 29380 46214
rect 29436 46212 29460 46214
rect 29220 46192 29516 46212
rect 39220 46268 39516 46288
rect 39276 46266 39300 46268
rect 39356 46266 39380 46268
rect 39436 46266 39460 46268
rect 39298 46214 39300 46266
rect 39362 46214 39374 46266
rect 39436 46214 39438 46266
rect 39276 46212 39300 46214
rect 39356 46212 39380 46214
rect 39436 46212 39460 46214
rect 39220 46192 39516 46212
rect 24220 45724 24516 45744
rect 24276 45722 24300 45724
rect 24356 45722 24380 45724
rect 24436 45722 24460 45724
rect 24298 45670 24300 45722
rect 24362 45670 24374 45722
rect 24436 45670 24438 45722
rect 24276 45668 24300 45670
rect 24356 45668 24380 45670
rect 24436 45668 24460 45670
rect 24220 45648 24516 45668
rect 34220 45724 34516 45744
rect 34276 45722 34300 45724
rect 34356 45722 34380 45724
rect 34436 45722 34460 45724
rect 34298 45670 34300 45722
rect 34362 45670 34374 45722
rect 34436 45670 34438 45722
rect 34276 45668 34300 45670
rect 34356 45668 34380 45670
rect 34436 45668 34460 45670
rect 34220 45648 34516 45668
rect 44220 45724 44516 45744
rect 44276 45722 44300 45724
rect 44356 45722 44380 45724
rect 44436 45722 44460 45724
rect 44298 45670 44300 45722
rect 44362 45670 44374 45722
rect 44436 45670 44438 45722
rect 44276 45668 44300 45670
rect 44356 45668 44380 45670
rect 44436 45668 44460 45670
rect 44220 45648 44516 45668
rect 19984 45484 20036 45490
rect 19984 45426 20036 45432
rect 19220 45180 19516 45200
rect 19276 45178 19300 45180
rect 19356 45178 19380 45180
rect 19436 45178 19460 45180
rect 19298 45126 19300 45178
rect 19362 45126 19374 45178
rect 19436 45126 19438 45178
rect 19276 45124 19300 45126
rect 19356 45124 19380 45126
rect 19436 45124 19460 45126
rect 19220 45104 19516 45124
rect 19220 44092 19516 44112
rect 19276 44090 19300 44092
rect 19356 44090 19380 44092
rect 19436 44090 19460 44092
rect 19298 44038 19300 44090
rect 19362 44038 19374 44090
rect 19436 44038 19438 44090
rect 19276 44036 19300 44038
rect 19356 44036 19380 44038
rect 19436 44036 19460 44038
rect 19220 44016 19516 44036
rect 19220 43004 19516 43024
rect 19276 43002 19300 43004
rect 19356 43002 19380 43004
rect 19436 43002 19460 43004
rect 19298 42950 19300 43002
rect 19362 42950 19374 43002
rect 19436 42950 19438 43002
rect 19276 42948 19300 42950
rect 19356 42948 19380 42950
rect 19436 42948 19460 42950
rect 19220 42928 19516 42948
rect 19220 41916 19516 41936
rect 19276 41914 19300 41916
rect 19356 41914 19380 41916
rect 19436 41914 19460 41916
rect 19298 41862 19300 41914
rect 19362 41862 19374 41914
rect 19436 41862 19438 41914
rect 19276 41860 19300 41862
rect 19356 41860 19380 41862
rect 19436 41860 19460 41862
rect 19220 41840 19516 41860
rect 19220 40828 19516 40848
rect 19276 40826 19300 40828
rect 19356 40826 19380 40828
rect 19436 40826 19460 40828
rect 19298 40774 19300 40826
rect 19362 40774 19374 40826
rect 19436 40774 19438 40826
rect 19276 40772 19300 40774
rect 19356 40772 19380 40774
rect 19436 40772 19460 40774
rect 19220 40752 19516 40772
rect 19220 39740 19516 39760
rect 19276 39738 19300 39740
rect 19356 39738 19380 39740
rect 19436 39738 19460 39740
rect 19298 39686 19300 39738
rect 19362 39686 19374 39738
rect 19436 39686 19438 39738
rect 19276 39684 19300 39686
rect 19356 39684 19380 39686
rect 19436 39684 19460 39686
rect 19220 39664 19516 39684
rect 19220 38652 19516 38672
rect 19276 38650 19300 38652
rect 19356 38650 19380 38652
rect 19436 38650 19460 38652
rect 19298 38598 19300 38650
rect 19362 38598 19374 38650
rect 19436 38598 19438 38650
rect 19276 38596 19300 38598
rect 19356 38596 19380 38598
rect 19436 38596 19460 38598
rect 19220 38576 19516 38596
rect 19220 37564 19516 37584
rect 19276 37562 19300 37564
rect 19356 37562 19380 37564
rect 19436 37562 19460 37564
rect 19298 37510 19300 37562
rect 19362 37510 19374 37562
rect 19436 37510 19438 37562
rect 19276 37508 19300 37510
rect 19356 37508 19380 37510
rect 19436 37508 19460 37510
rect 19220 37488 19516 37508
rect 19996 36922 20024 45426
rect 25780 45348 25832 45354
rect 25780 45290 25832 45296
rect 24220 44636 24516 44656
rect 24276 44634 24300 44636
rect 24356 44634 24380 44636
rect 24436 44634 24460 44636
rect 24298 44582 24300 44634
rect 24362 44582 24374 44634
rect 24436 44582 24438 44634
rect 24276 44580 24300 44582
rect 24356 44580 24380 44582
rect 24436 44580 24460 44582
rect 24220 44560 24516 44580
rect 24220 43548 24516 43568
rect 24276 43546 24300 43548
rect 24356 43546 24380 43548
rect 24436 43546 24460 43548
rect 24298 43494 24300 43546
rect 24362 43494 24374 43546
rect 24436 43494 24438 43546
rect 24276 43492 24300 43494
rect 24356 43492 24380 43494
rect 24436 43492 24460 43494
rect 24220 43472 24516 43492
rect 24220 42460 24516 42480
rect 24276 42458 24300 42460
rect 24356 42458 24380 42460
rect 24436 42458 24460 42460
rect 24298 42406 24300 42458
rect 24362 42406 24374 42458
rect 24436 42406 24438 42458
rect 24276 42404 24300 42406
rect 24356 42404 24380 42406
rect 24436 42404 24460 42406
rect 24220 42384 24516 42404
rect 24220 41372 24516 41392
rect 24276 41370 24300 41372
rect 24356 41370 24380 41372
rect 24436 41370 24460 41372
rect 24298 41318 24300 41370
rect 24362 41318 24374 41370
rect 24436 41318 24438 41370
rect 24276 41316 24300 41318
rect 24356 41316 24380 41318
rect 24436 41316 24460 41318
rect 24220 41296 24516 41316
rect 24220 40284 24516 40304
rect 24276 40282 24300 40284
rect 24356 40282 24380 40284
rect 24436 40282 24460 40284
rect 24298 40230 24300 40282
rect 24362 40230 24374 40282
rect 24436 40230 24438 40282
rect 24276 40228 24300 40230
rect 24356 40228 24380 40230
rect 24436 40228 24460 40230
rect 24220 40208 24516 40228
rect 23112 39500 23164 39506
rect 23112 39442 23164 39448
rect 21916 39432 21968 39438
rect 21916 39374 21968 39380
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19220 36476 19516 36496
rect 19276 36474 19300 36476
rect 19356 36474 19380 36476
rect 19436 36474 19460 36476
rect 19298 36422 19300 36474
rect 19362 36422 19374 36474
rect 19436 36422 19438 36474
rect 19276 36420 19300 36422
rect 19356 36420 19380 36422
rect 19436 36420 19460 36422
rect 19220 36400 19516 36420
rect 19220 35388 19516 35408
rect 19276 35386 19300 35388
rect 19356 35386 19380 35388
rect 19436 35386 19460 35388
rect 19298 35334 19300 35386
rect 19362 35334 19374 35386
rect 19436 35334 19438 35386
rect 19276 35332 19300 35334
rect 19356 35332 19380 35334
rect 19436 35332 19460 35334
rect 19220 35312 19516 35332
rect 19220 34300 19516 34320
rect 19276 34298 19300 34300
rect 19356 34298 19380 34300
rect 19436 34298 19460 34300
rect 19298 34246 19300 34298
rect 19362 34246 19374 34298
rect 19436 34246 19438 34298
rect 19276 34244 19300 34246
rect 19356 34244 19380 34246
rect 19436 34244 19460 34246
rect 19220 34224 19516 34244
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16040 14006 16068 14214
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15120 13190 15148 13874
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 14220 13084 14516 13104
rect 14276 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14298 13030 14300 13082
rect 14362 13030 14374 13082
rect 14436 13030 14438 13082
rect 14276 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14220 13008 14516 13028
rect 14220 11996 14516 12016
rect 14276 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14298 11942 14300 11994
rect 14362 11942 14374 11994
rect 14436 11942 14438 11994
rect 14276 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14220 11920 14516 11940
rect 15120 11626 15148 13126
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 14220 10908 14516 10928
rect 14276 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14298 10854 14300 10906
rect 14362 10854 14374 10906
rect 14436 10854 14438 10906
rect 14276 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14220 10832 14516 10852
rect 14220 9820 14516 9840
rect 14276 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14298 9766 14300 9818
rect 14362 9766 14374 9818
rect 14436 9766 14438 9818
rect 14276 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14220 9744 14516 9764
rect 14220 8732 14516 8752
rect 14276 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14298 8678 14300 8730
rect 14362 8678 14374 8730
rect 14436 8678 14438 8730
rect 14276 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14220 8656 14516 8676
rect 14220 7644 14516 7664
rect 14276 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14298 7590 14300 7642
rect 14362 7590 14374 7642
rect 14436 7590 14438 7642
rect 14276 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14220 7568 14516 7588
rect 14220 6556 14516 6576
rect 14276 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14298 6502 14300 6554
rect 14362 6502 14374 6554
rect 14436 6502 14438 6554
rect 14276 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14220 6480 14516 6500
rect 15948 6458 15976 13874
rect 16040 11121 16068 13942
rect 16408 13802 16436 13942
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16408 13530 16436 13738
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16868 12102 16896 14214
rect 17236 13938 17264 15642
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17420 13258 17448 33934
rect 18328 33448 18380 33454
rect 18328 33390 18380 33396
rect 18236 30388 18288 30394
rect 18236 30330 18288 30336
rect 18248 28422 18276 30330
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17972 26382 18000 26930
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17512 23866 17540 24006
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17868 19236 17920 19242
rect 17868 19178 17920 19184
rect 17880 16574 17908 19178
rect 17788 16546 17908 16574
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17696 13938 17724 14418
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17788 13870 17816 16546
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15570 17908 15846
rect 17972 15638 18000 26318
rect 18144 25696 18196 25702
rect 18144 25638 18196 25644
rect 18156 19854 18184 25638
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18064 17270 18092 17478
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16026 11112 16082 11121
rect 16026 11047 16082 11056
rect 17420 8090 17448 13194
rect 17788 13190 17816 13806
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 8362 17816 13126
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17880 7342 17908 15506
rect 17972 15162 18000 15574
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18064 14906 18092 17206
rect 18156 16250 18184 19790
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18156 15570 18184 16186
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18064 14878 18184 14906
rect 18156 14822 18184 14878
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18156 14074 18184 14758
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17972 7274 18000 8230
rect 18064 7954 18092 8230
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 18064 7041 18092 7890
rect 18050 7032 18106 7041
rect 18050 6967 18106 6976
rect 18156 6914 18184 14010
rect 18248 13802 18276 28358
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18248 13190 18276 13738
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18064 6886 18184 6914
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17972 5778 18000 6054
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 14220 5468 14516 5488
rect 14276 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14298 5414 14300 5466
rect 14362 5414 14374 5466
rect 14436 5414 14438 5466
rect 14276 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14220 5392 14516 5412
rect 17972 5030 18000 5578
rect 18064 5302 18092 6886
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 5846 18184 6598
rect 18248 6474 18276 13126
rect 18340 6662 18368 33390
rect 19220 33212 19516 33232
rect 19276 33210 19300 33212
rect 19356 33210 19380 33212
rect 19436 33210 19460 33212
rect 19298 33158 19300 33210
rect 19362 33158 19374 33210
rect 19436 33158 19438 33210
rect 19276 33156 19300 33158
rect 19356 33156 19380 33158
rect 19436 33156 19460 33158
rect 19220 33136 19516 33156
rect 19220 32124 19516 32144
rect 19276 32122 19300 32124
rect 19356 32122 19380 32124
rect 19436 32122 19460 32124
rect 19298 32070 19300 32122
rect 19362 32070 19374 32122
rect 19436 32070 19438 32122
rect 19276 32068 19300 32070
rect 19356 32068 19380 32070
rect 19436 32068 19460 32070
rect 19220 32048 19516 32068
rect 19220 31036 19516 31056
rect 19276 31034 19300 31036
rect 19356 31034 19380 31036
rect 19436 31034 19460 31036
rect 19298 30982 19300 31034
rect 19362 30982 19374 31034
rect 19436 30982 19438 31034
rect 19276 30980 19300 30982
rect 19356 30980 19380 30982
rect 19436 30980 19460 30982
rect 19220 30960 19516 30980
rect 19220 29948 19516 29968
rect 19276 29946 19300 29948
rect 19356 29946 19380 29948
rect 19436 29946 19460 29948
rect 19298 29894 19300 29946
rect 19362 29894 19374 29946
rect 19436 29894 19438 29946
rect 19276 29892 19300 29894
rect 19356 29892 19380 29894
rect 19436 29892 19460 29894
rect 19220 29872 19516 29892
rect 19220 28860 19516 28880
rect 19276 28858 19300 28860
rect 19356 28858 19380 28860
rect 19436 28858 19460 28860
rect 19298 28806 19300 28858
rect 19362 28806 19374 28858
rect 19436 28806 19438 28858
rect 19276 28804 19300 28806
rect 19356 28804 19380 28806
rect 19436 28804 19460 28806
rect 19220 28784 19516 28804
rect 19220 27772 19516 27792
rect 19276 27770 19300 27772
rect 19356 27770 19380 27772
rect 19436 27770 19460 27772
rect 19298 27718 19300 27770
rect 19362 27718 19374 27770
rect 19436 27718 19438 27770
rect 19276 27716 19300 27718
rect 19356 27716 19380 27718
rect 19436 27716 19460 27718
rect 19220 27696 19516 27716
rect 19996 26926 20024 36858
rect 21364 36304 21416 36310
rect 21364 36246 21416 36252
rect 21376 28762 21404 36246
rect 21548 35488 21600 35494
rect 21548 35430 21600 35436
rect 21560 32026 21588 35430
rect 21548 32020 21600 32026
rect 21548 31962 21600 31968
rect 21928 31142 21956 39374
rect 22744 39364 22796 39370
rect 22744 39306 22796 39312
rect 22560 39296 22612 39302
rect 22560 39238 22612 39244
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21364 28756 21416 28762
rect 21364 28698 21416 28704
rect 21928 27470 21956 31078
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 22020 28014 22048 28698
rect 22008 28008 22060 28014
rect 22008 27950 22060 27956
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 19984 26920 20036 26926
rect 19984 26862 20036 26868
rect 19220 26684 19516 26704
rect 19276 26682 19300 26684
rect 19356 26682 19380 26684
rect 19436 26682 19460 26684
rect 19298 26630 19300 26682
rect 19362 26630 19374 26682
rect 19436 26630 19438 26682
rect 19276 26628 19300 26630
rect 19356 26628 19380 26630
rect 19436 26628 19460 26630
rect 19220 26608 19516 26628
rect 19220 25596 19516 25616
rect 19276 25594 19300 25596
rect 19356 25594 19380 25596
rect 19436 25594 19460 25596
rect 19298 25542 19300 25594
rect 19362 25542 19374 25594
rect 19436 25542 19438 25594
rect 19276 25540 19300 25542
rect 19356 25540 19380 25542
rect 19436 25540 19460 25542
rect 19220 25520 19516 25540
rect 19220 24508 19516 24528
rect 19276 24506 19300 24508
rect 19356 24506 19380 24508
rect 19436 24506 19460 24508
rect 19298 24454 19300 24506
rect 19362 24454 19374 24506
rect 19436 24454 19438 24506
rect 19276 24452 19300 24454
rect 19356 24452 19380 24454
rect 19436 24452 19460 24454
rect 19220 24432 19516 24452
rect 19996 24410 20024 26862
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19220 23420 19516 23440
rect 19276 23418 19300 23420
rect 19356 23418 19380 23420
rect 19436 23418 19460 23420
rect 19298 23366 19300 23418
rect 19362 23366 19374 23418
rect 19436 23366 19438 23418
rect 19276 23364 19300 23366
rect 19356 23364 19380 23366
rect 19436 23364 19460 23366
rect 19220 23344 19516 23364
rect 19220 22332 19516 22352
rect 19276 22330 19300 22332
rect 19356 22330 19380 22332
rect 19436 22330 19460 22332
rect 19298 22278 19300 22330
rect 19362 22278 19374 22330
rect 19436 22278 19438 22330
rect 19276 22276 19300 22278
rect 19356 22276 19380 22278
rect 19436 22276 19460 22278
rect 19220 22256 19516 22276
rect 18420 21888 18472 21894
rect 18420 21830 18472 21836
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18248 6446 18368 6474
rect 18340 6118 18368 6446
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 18248 4826 18276 5714
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 14220 4380 14516 4400
rect 14276 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14298 4326 14300 4378
rect 14362 4326 14374 4378
rect 14436 4326 14438 4378
rect 14276 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14220 4304 14516 4324
rect 18340 3602 18368 6054
rect 18432 5914 18460 21830
rect 19220 21244 19516 21264
rect 19276 21242 19300 21244
rect 19356 21242 19380 21244
rect 19436 21242 19460 21244
rect 19298 21190 19300 21242
rect 19362 21190 19374 21242
rect 19436 21190 19438 21242
rect 19276 21188 19300 21190
rect 19356 21188 19380 21190
rect 19436 21188 19460 21190
rect 19220 21168 19516 21188
rect 19220 20156 19516 20176
rect 19276 20154 19300 20156
rect 19356 20154 19380 20156
rect 19436 20154 19460 20156
rect 19298 20102 19300 20154
rect 19362 20102 19374 20154
rect 19436 20102 19438 20154
rect 19276 20100 19300 20102
rect 19356 20100 19380 20102
rect 19436 20100 19460 20102
rect 19220 20080 19516 20100
rect 22572 15094 22600 39238
rect 22756 38758 22784 39306
rect 22744 38752 22796 38758
rect 22744 38694 22796 38700
rect 22756 30598 22784 38694
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 23124 29646 23152 39442
rect 23664 39296 23716 39302
rect 23664 39238 23716 39244
rect 24584 39296 24636 39302
rect 24584 39238 24636 39244
rect 24768 39296 24820 39302
rect 24768 39238 24820 39244
rect 23676 39030 23704 39238
rect 24220 39196 24516 39216
rect 24276 39194 24300 39196
rect 24356 39194 24380 39196
rect 24436 39194 24460 39196
rect 24298 39142 24300 39194
rect 24362 39142 24374 39194
rect 24436 39142 24438 39194
rect 24276 39140 24300 39142
rect 24356 39140 24380 39142
rect 24436 39140 24460 39142
rect 24220 39120 24516 39140
rect 24596 39098 24624 39238
rect 24584 39092 24636 39098
rect 24584 39034 24636 39040
rect 23664 39024 23716 39030
rect 23664 38966 23716 38972
rect 24676 38888 24728 38894
rect 24676 38830 24728 38836
rect 23940 38752 23992 38758
rect 23940 38694 23992 38700
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23020 28620 23072 28626
rect 23020 28562 23072 28568
rect 23032 28014 23060 28562
rect 23020 28008 23072 28014
rect 23020 27950 23072 27956
rect 22652 27940 22704 27946
rect 22652 27882 22704 27888
rect 22560 15088 22612 15094
rect 22560 15030 22612 15036
rect 22664 14618 22692 27882
rect 23032 27606 23060 27950
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23492 20058 23520 24142
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18524 14074 18552 14350
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21744 6225 21772 7210
rect 21822 7032 21878 7041
rect 21822 6967 21878 6976
rect 21836 6361 21864 6967
rect 21822 6352 21878 6361
rect 21822 6287 21878 6296
rect 21730 6216 21786 6225
rect 21730 6151 21786 6160
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 23952 5778 23980 38694
rect 24124 38412 24176 38418
rect 24124 38354 24176 38360
rect 24136 36174 24164 38354
rect 24220 38108 24516 38128
rect 24276 38106 24300 38108
rect 24356 38106 24380 38108
rect 24436 38106 24460 38108
rect 24298 38054 24300 38106
rect 24362 38054 24374 38106
rect 24436 38054 24438 38106
rect 24276 38052 24300 38054
rect 24356 38052 24380 38054
rect 24436 38052 24460 38054
rect 24220 38032 24516 38052
rect 24220 37020 24516 37040
rect 24276 37018 24300 37020
rect 24356 37018 24380 37020
rect 24436 37018 24460 37020
rect 24298 36966 24300 37018
rect 24362 36966 24374 37018
rect 24436 36966 24438 37018
rect 24276 36964 24300 36966
rect 24356 36964 24380 36966
rect 24436 36964 24460 36966
rect 24220 36944 24516 36964
rect 24124 36168 24176 36174
rect 24124 36110 24176 36116
rect 24136 28218 24164 36110
rect 24220 35932 24516 35952
rect 24276 35930 24300 35932
rect 24356 35930 24380 35932
rect 24436 35930 24460 35932
rect 24298 35878 24300 35930
rect 24362 35878 24374 35930
rect 24436 35878 24438 35930
rect 24276 35876 24300 35878
rect 24356 35876 24380 35878
rect 24436 35876 24460 35878
rect 24220 35856 24516 35876
rect 24220 34844 24516 34864
rect 24276 34842 24300 34844
rect 24356 34842 24380 34844
rect 24436 34842 24460 34844
rect 24298 34790 24300 34842
rect 24362 34790 24374 34842
rect 24436 34790 24438 34842
rect 24276 34788 24300 34790
rect 24356 34788 24380 34790
rect 24436 34788 24460 34790
rect 24220 34768 24516 34788
rect 24220 33756 24516 33776
rect 24276 33754 24300 33756
rect 24356 33754 24380 33756
rect 24436 33754 24460 33756
rect 24298 33702 24300 33754
rect 24362 33702 24374 33754
rect 24436 33702 24438 33754
rect 24276 33700 24300 33702
rect 24356 33700 24380 33702
rect 24436 33700 24460 33702
rect 24220 33680 24516 33700
rect 24220 32668 24516 32688
rect 24276 32666 24300 32668
rect 24356 32666 24380 32668
rect 24436 32666 24460 32668
rect 24298 32614 24300 32666
rect 24362 32614 24374 32666
rect 24436 32614 24438 32666
rect 24276 32612 24300 32614
rect 24356 32612 24380 32614
rect 24436 32612 24460 32614
rect 24220 32592 24516 32612
rect 24688 32570 24716 38830
rect 24780 38826 24808 39238
rect 24768 38820 24820 38826
rect 24768 38762 24820 38768
rect 24676 32564 24728 32570
rect 24676 32506 24728 32512
rect 24220 31580 24516 31600
rect 24276 31578 24300 31580
rect 24356 31578 24380 31580
rect 24436 31578 24460 31580
rect 24298 31526 24300 31578
rect 24362 31526 24374 31578
rect 24436 31526 24438 31578
rect 24276 31524 24300 31526
rect 24356 31524 24380 31526
rect 24436 31524 24460 31526
rect 24220 31504 24516 31524
rect 24220 30492 24516 30512
rect 24276 30490 24300 30492
rect 24356 30490 24380 30492
rect 24436 30490 24460 30492
rect 24298 30438 24300 30490
rect 24362 30438 24374 30490
rect 24436 30438 24438 30490
rect 24276 30436 24300 30438
rect 24356 30436 24380 30438
rect 24436 30436 24460 30438
rect 24220 30416 24516 30436
rect 24220 29404 24516 29424
rect 24276 29402 24300 29404
rect 24356 29402 24380 29404
rect 24436 29402 24460 29404
rect 24298 29350 24300 29402
rect 24362 29350 24374 29402
rect 24436 29350 24438 29402
rect 24276 29348 24300 29350
rect 24356 29348 24380 29350
rect 24436 29348 24460 29350
rect 24220 29328 24516 29348
rect 24688 28370 24716 32506
rect 25688 31340 25740 31346
rect 25688 31282 25740 31288
rect 25044 29028 25096 29034
rect 25044 28970 25096 28976
rect 24596 28342 24716 28370
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24220 28316 24516 28336
rect 24276 28314 24300 28316
rect 24356 28314 24380 28316
rect 24436 28314 24460 28316
rect 24298 28262 24300 28314
rect 24362 28262 24374 28314
rect 24436 28262 24438 28314
rect 24276 28260 24300 28262
rect 24356 28260 24380 28262
rect 24436 28260 24460 28262
rect 24220 28240 24516 28260
rect 24124 28212 24176 28218
rect 24124 28154 24176 28160
rect 24596 28082 24624 28342
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24220 27228 24516 27248
rect 24276 27226 24300 27228
rect 24356 27226 24380 27228
rect 24436 27226 24460 27228
rect 24298 27174 24300 27226
rect 24362 27174 24374 27226
rect 24436 27174 24438 27226
rect 24276 27172 24300 27174
rect 24356 27172 24380 27174
rect 24436 27172 24460 27174
rect 24220 27152 24516 27172
rect 24220 26140 24516 26160
rect 24276 26138 24300 26140
rect 24356 26138 24380 26140
rect 24436 26138 24460 26140
rect 24298 26086 24300 26138
rect 24362 26086 24374 26138
rect 24436 26086 24438 26138
rect 24276 26084 24300 26086
rect 24356 26084 24380 26086
rect 24436 26084 24460 26086
rect 24220 26064 24516 26084
rect 24220 25052 24516 25072
rect 24276 25050 24300 25052
rect 24356 25050 24380 25052
rect 24436 25050 24460 25052
rect 24298 24998 24300 25050
rect 24362 24998 24374 25050
rect 24436 24998 24438 25050
rect 24276 24996 24300 24998
rect 24356 24996 24380 24998
rect 24436 24996 24460 24998
rect 24220 24976 24516 24996
rect 24220 23964 24516 23984
rect 24276 23962 24300 23964
rect 24356 23962 24380 23964
rect 24436 23962 24460 23964
rect 24298 23910 24300 23962
rect 24362 23910 24374 23962
rect 24436 23910 24438 23962
rect 24276 23908 24300 23910
rect 24356 23908 24380 23910
rect 24436 23908 24460 23910
rect 24220 23888 24516 23908
rect 24688 23186 24716 28154
rect 24780 27878 24808 28154
rect 24872 28082 24900 28358
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24768 27872 24820 27878
rect 24768 27814 24820 27820
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24220 22876 24516 22896
rect 24276 22874 24300 22876
rect 24356 22874 24380 22876
rect 24436 22874 24460 22876
rect 24298 22822 24300 22874
rect 24362 22822 24374 22874
rect 24436 22822 24438 22874
rect 24276 22820 24300 22822
rect 24356 22820 24380 22822
rect 24436 22820 24460 22822
rect 24220 22800 24516 22820
rect 24220 21788 24516 21808
rect 24276 21786 24300 21788
rect 24356 21786 24380 21788
rect 24436 21786 24460 21788
rect 24298 21734 24300 21786
rect 24362 21734 24374 21786
rect 24436 21734 24438 21786
rect 24276 21732 24300 21734
rect 24356 21732 24380 21734
rect 24436 21732 24460 21734
rect 24220 21712 24516 21732
rect 24220 20700 24516 20720
rect 24276 20698 24300 20700
rect 24356 20698 24380 20700
rect 24436 20698 24460 20700
rect 24298 20646 24300 20698
rect 24362 20646 24374 20698
rect 24436 20646 24438 20698
rect 24276 20644 24300 20646
rect 24356 20644 24380 20646
rect 24436 20644 24460 20646
rect 24220 20624 24516 20644
rect 24220 19612 24516 19632
rect 24276 19610 24300 19612
rect 24356 19610 24380 19612
rect 24436 19610 24460 19612
rect 24298 19558 24300 19610
rect 24362 19558 24374 19610
rect 24436 19558 24438 19610
rect 24276 19556 24300 19558
rect 24356 19556 24380 19558
rect 24436 19556 24460 19558
rect 24220 19536 24516 19556
rect 25056 16574 25084 28970
rect 25700 23322 25728 31282
rect 25792 29646 25820 45290
rect 29220 45180 29516 45200
rect 29276 45178 29300 45180
rect 29356 45178 29380 45180
rect 29436 45178 29460 45180
rect 29298 45126 29300 45178
rect 29362 45126 29374 45178
rect 29436 45126 29438 45178
rect 29276 45124 29300 45126
rect 29356 45124 29380 45126
rect 29436 45124 29460 45126
rect 29220 45104 29516 45124
rect 39220 45180 39516 45200
rect 39276 45178 39300 45180
rect 39356 45178 39380 45180
rect 39436 45178 39460 45180
rect 39298 45126 39300 45178
rect 39362 45126 39374 45178
rect 39436 45126 39438 45178
rect 39276 45124 39300 45126
rect 39356 45124 39380 45126
rect 39436 45124 39460 45126
rect 39220 45104 39516 45124
rect 34220 44636 34516 44656
rect 34276 44634 34300 44636
rect 34356 44634 34380 44636
rect 34436 44634 34460 44636
rect 34298 44582 34300 44634
rect 34362 44582 34374 44634
rect 34436 44582 34438 44634
rect 34276 44580 34300 44582
rect 34356 44580 34380 44582
rect 34436 44580 34460 44582
rect 34220 44560 34516 44580
rect 44220 44636 44516 44656
rect 44276 44634 44300 44636
rect 44356 44634 44380 44636
rect 44436 44634 44460 44636
rect 44298 44582 44300 44634
rect 44362 44582 44374 44634
rect 44436 44582 44438 44634
rect 44276 44580 44300 44582
rect 44356 44580 44380 44582
rect 44436 44580 44460 44582
rect 44220 44560 44516 44580
rect 29220 44092 29516 44112
rect 29276 44090 29300 44092
rect 29356 44090 29380 44092
rect 29436 44090 29460 44092
rect 29298 44038 29300 44090
rect 29362 44038 29374 44090
rect 29436 44038 29438 44090
rect 29276 44036 29300 44038
rect 29356 44036 29380 44038
rect 29436 44036 29460 44038
rect 29220 44016 29516 44036
rect 39220 44092 39516 44112
rect 39276 44090 39300 44092
rect 39356 44090 39380 44092
rect 39436 44090 39460 44092
rect 39298 44038 39300 44090
rect 39362 44038 39374 44090
rect 39436 44038 39438 44090
rect 39276 44036 39300 44038
rect 39356 44036 39380 44038
rect 39436 44036 39460 44038
rect 39220 44016 39516 44036
rect 34220 43548 34516 43568
rect 34276 43546 34300 43548
rect 34356 43546 34380 43548
rect 34436 43546 34460 43548
rect 34298 43494 34300 43546
rect 34362 43494 34374 43546
rect 34436 43494 34438 43546
rect 34276 43492 34300 43494
rect 34356 43492 34380 43494
rect 34436 43492 34460 43494
rect 34220 43472 34516 43492
rect 44220 43548 44516 43568
rect 44276 43546 44300 43548
rect 44356 43546 44380 43548
rect 44436 43546 44460 43548
rect 44298 43494 44300 43546
rect 44362 43494 44374 43546
rect 44436 43494 44438 43546
rect 44276 43492 44300 43494
rect 44356 43492 44380 43494
rect 44436 43492 44460 43494
rect 44220 43472 44516 43492
rect 29220 43004 29516 43024
rect 29276 43002 29300 43004
rect 29356 43002 29380 43004
rect 29436 43002 29460 43004
rect 29298 42950 29300 43002
rect 29362 42950 29374 43002
rect 29436 42950 29438 43002
rect 29276 42948 29300 42950
rect 29356 42948 29380 42950
rect 29436 42948 29460 42950
rect 29220 42928 29516 42948
rect 39220 43004 39516 43024
rect 39276 43002 39300 43004
rect 39356 43002 39380 43004
rect 39436 43002 39460 43004
rect 39298 42950 39300 43002
rect 39362 42950 39374 43002
rect 39436 42950 39438 43002
rect 39276 42948 39300 42950
rect 39356 42948 39380 42950
rect 39436 42948 39460 42950
rect 39220 42928 39516 42948
rect 39672 42764 39724 42770
rect 39672 42706 39724 42712
rect 42800 42764 42852 42770
rect 42800 42706 42852 42712
rect 35348 42696 35400 42702
rect 35348 42638 35400 42644
rect 34220 42460 34516 42480
rect 34276 42458 34300 42460
rect 34356 42458 34380 42460
rect 34436 42458 34460 42460
rect 34298 42406 34300 42458
rect 34362 42406 34374 42458
rect 34436 42406 34438 42458
rect 34276 42404 34300 42406
rect 34356 42404 34380 42406
rect 34436 42404 34460 42406
rect 34220 42384 34516 42404
rect 29220 41916 29516 41936
rect 29276 41914 29300 41916
rect 29356 41914 29380 41916
rect 29436 41914 29460 41916
rect 29298 41862 29300 41914
rect 29362 41862 29374 41914
rect 29436 41862 29438 41914
rect 29276 41860 29300 41862
rect 29356 41860 29380 41862
rect 29436 41860 29460 41862
rect 29220 41840 29516 41860
rect 34220 41372 34516 41392
rect 34276 41370 34300 41372
rect 34356 41370 34380 41372
rect 34436 41370 34460 41372
rect 34298 41318 34300 41370
rect 34362 41318 34374 41370
rect 34436 41318 34438 41370
rect 34276 41316 34300 41318
rect 34356 41316 34380 41318
rect 34436 41316 34460 41318
rect 34220 41296 34516 41316
rect 29220 40828 29516 40848
rect 29276 40826 29300 40828
rect 29356 40826 29380 40828
rect 29436 40826 29460 40828
rect 29298 40774 29300 40826
rect 29362 40774 29374 40826
rect 29436 40774 29438 40826
rect 29276 40772 29300 40774
rect 29356 40772 29380 40774
rect 29436 40772 29460 40774
rect 29220 40752 29516 40772
rect 34220 40284 34516 40304
rect 34276 40282 34300 40284
rect 34356 40282 34380 40284
rect 34436 40282 34460 40284
rect 34298 40230 34300 40282
rect 34362 40230 34374 40282
rect 34436 40230 34438 40282
rect 34276 40228 34300 40230
rect 34356 40228 34380 40230
rect 34436 40228 34460 40230
rect 34220 40208 34516 40228
rect 29220 39740 29516 39760
rect 29276 39738 29300 39740
rect 29356 39738 29380 39740
rect 29436 39738 29460 39740
rect 29298 39686 29300 39738
rect 29362 39686 29374 39738
rect 29436 39686 29438 39738
rect 29276 39684 29300 39686
rect 29356 39684 29380 39686
rect 29436 39684 29460 39686
rect 29220 39664 29516 39684
rect 35360 39642 35388 42638
rect 38936 42628 38988 42634
rect 38936 42570 38988 42576
rect 35348 39636 35400 39642
rect 35348 39578 35400 39584
rect 34220 39196 34516 39216
rect 34276 39194 34300 39196
rect 34356 39194 34380 39196
rect 34436 39194 34460 39196
rect 34298 39142 34300 39194
rect 34362 39142 34374 39194
rect 34436 39142 34438 39194
rect 34276 39140 34300 39142
rect 34356 39140 34380 39142
rect 34436 39140 34460 39142
rect 34220 39120 34516 39140
rect 32864 39024 32916 39030
rect 32864 38966 32916 38972
rect 32876 38894 32904 38966
rect 32864 38888 32916 38894
rect 32864 38830 32916 38836
rect 33508 38888 33560 38894
rect 33508 38830 33560 38836
rect 29092 38752 29144 38758
rect 29092 38694 29144 38700
rect 29104 38350 29132 38694
rect 29220 38652 29516 38672
rect 29276 38650 29300 38652
rect 29356 38650 29380 38652
rect 29436 38650 29460 38652
rect 29298 38598 29300 38650
rect 29362 38598 29374 38650
rect 29436 38598 29438 38650
rect 29276 38596 29300 38598
rect 29356 38596 29380 38598
rect 29436 38596 29460 38598
rect 29220 38576 29516 38596
rect 32876 38554 32904 38830
rect 33232 38820 33284 38826
rect 33232 38762 33284 38768
rect 32864 38548 32916 38554
rect 32864 38490 32916 38496
rect 29092 38344 29144 38350
rect 29092 38286 29144 38292
rect 27712 38208 27764 38214
rect 27712 38150 27764 38156
rect 28080 38208 28132 38214
rect 28080 38150 28132 38156
rect 29000 38208 29052 38214
rect 29000 38150 29052 38156
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 26056 29640 26108 29646
rect 26056 29582 26108 29588
rect 25792 26994 25820 29582
rect 26068 29034 26096 29582
rect 26056 29028 26108 29034
rect 26056 28970 26108 28976
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25688 23316 25740 23322
rect 25688 23258 25740 23264
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27264 19990 27292 20198
rect 27252 19984 27304 19990
rect 27252 19926 27304 19932
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 27540 19718 27568 19858
rect 27528 19712 27580 19718
rect 27528 19654 27580 19660
rect 27540 18630 27568 19654
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27724 16590 27752 38150
rect 28092 37670 28120 38150
rect 28080 37664 28132 37670
rect 28080 37606 28132 37612
rect 29012 35494 29040 38150
rect 29104 37942 29132 38286
rect 29092 37936 29144 37942
rect 29092 37878 29144 37884
rect 29220 37564 29516 37584
rect 29276 37562 29300 37564
rect 29356 37562 29380 37564
rect 29436 37562 29460 37564
rect 29298 37510 29300 37562
rect 29362 37510 29374 37562
rect 29436 37510 29438 37562
rect 29276 37508 29300 37510
rect 29356 37508 29380 37510
rect 29436 37508 29460 37510
rect 29220 37488 29516 37508
rect 29220 36476 29516 36496
rect 29276 36474 29300 36476
rect 29356 36474 29380 36476
rect 29436 36474 29460 36476
rect 29298 36422 29300 36474
rect 29362 36422 29374 36474
rect 29436 36422 29438 36474
rect 29276 36420 29300 36422
rect 29356 36420 29380 36422
rect 29436 36420 29460 36422
rect 29220 36400 29516 36420
rect 29000 35488 29052 35494
rect 29000 35430 29052 35436
rect 28264 33380 28316 33386
rect 28264 33322 28316 33328
rect 28276 27538 28304 33322
rect 29012 28490 29040 35430
rect 29220 35388 29516 35408
rect 29276 35386 29300 35388
rect 29356 35386 29380 35388
rect 29436 35386 29460 35388
rect 29298 35334 29300 35386
rect 29362 35334 29374 35386
rect 29436 35334 29438 35386
rect 29276 35332 29300 35334
rect 29356 35332 29380 35334
rect 29436 35332 29460 35334
rect 29220 35312 29516 35332
rect 29220 34300 29516 34320
rect 29276 34298 29300 34300
rect 29356 34298 29380 34300
rect 29436 34298 29460 34300
rect 29298 34246 29300 34298
rect 29362 34246 29374 34298
rect 29436 34246 29438 34298
rect 29276 34244 29300 34246
rect 29356 34244 29380 34246
rect 29436 34244 29460 34246
rect 29220 34224 29516 34244
rect 29220 33212 29516 33232
rect 29276 33210 29300 33212
rect 29356 33210 29380 33212
rect 29436 33210 29460 33212
rect 29298 33158 29300 33210
rect 29362 33158 29374 33210
rect 29436 33158 29438 33210
rect 29276 33156 29300 33158
rect 29356 33156 29380 33158
rect 29436 33156 29460 33158
rect 29220 33136 29516 33156
rect 33140 33108 33192 33114
rect 33140 33050 33192 33056
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29220 32124 29516 32144
rect 29276 32122 29300 32124
rect 29356 32122 29380 32124
rect 29436 32122 29460 32124
rect 29298 32070 29300 32122
rect 29362 32070 29374 32122
rect 29436 32070 29438 32122
rect 29276 32068 29300 32070
rect 29356 32068 29380 32070
rect 29436 32068 29460 32070
rect 29220 32048 29516 32068
rect 29220 31036 29516 31056
rect 29276 31034 29300 31036
rect 29356 31034 29380 31036
rect 29436 31034 29460 31036
rect 29298 30982 29300 31034
rect 29362 30982 29374 31034
rect 29436 30982 29438 31034
rect 29276 30980 29300 30982
rect 29356 30980 29380 30982
rect 29436 30980 29460 30982
rect 29220 30960 29516 30980
rect 29220 29948 29516 29968
rect 29276 29946 29300 29948
rect 29356 29946 29380 29948
rect 29436 29946 29460 29948
rect 29298 29894 29300 29946
rect 29362 29894 29374 29946
rect 29436 29894 29438 29946
rect 29276 29892 29300 29894
rect 29356 29892 29380 29894
rect 29436 29892 29460 29894
rect 29220 29872 29516 29892
rect 29220 28860 29516 28880
rect 29276 28858 29300 28860
rect 29356 28858 29380 28860
rect 29436 28858 29460 28860
rect 29298 28806 29300 28858
rect 29362 28806 29374 28858
rect 29436 28806 29438 28858
rect 29276 28804 29300 28806
rect 29356 28804 29380 28806
rect 29436 28804 29460 28806
rect 29220 28784 29516 28804
rect 29000 28484 29052 28490
rect 29000 28426 29052 28432
rect 29220 27772 29516 27792
rect 29276 27770 29300 27772
rect 29356 27770 29380 27772
rect 29436 27770 29460 27772
rect 29298 27718 29300 27770
rect 29362 27718 29374 27770
rect 29436 27718 29438 27770
rect 29276 27716 29300 27718
rect 29356 27716 29380 27718
rect 29436 27716 29460 27718
rect 29220 27696 29516 27716
rect 28264 27532 28316 27538
rect 28264 27474 28316 27480
rect 28276 21962 28304 27474
rect 29220 26684 29516 26704
rect 29276 26682 29300 26684
rect 29356 26682 29380 26684
rect 29436 26682 29460 26684
rect 29298 26630 29300 26682
rect 29362 26630 29374 26682
rect 29436 26630 29438 26682
rect 29276 26628 29300 26630
rect 29356 26628 29380 26630
rect 29436 26628 29460 26630
rect 29220 26608 29516 26628
rect 29220 25596 29516 25616
rect 29276 25594 29300 25596
rect 29356 25594 29380 25596
rect 29436 25594 29460 25596
rect 29298 25542 29300 25594
rect 29362 25542 29374 25594
rect 29436 25542 29438 25594
rect 29276 25540 29300 25542
rect 29356 25540 29380 25542
rect 29436 25540 29460 25542
rect 29220 25520 29516 25540
rect 29748 24614 29776 32914
rect 32404 32768 32456 32774
rect 32404 32710 32456 32716
rect 31852 30864 31904 30870
rect 31852 30806 31904 30812
rect 31864 30054 31892 30806
rect 32416 30734 32444 32710
rect 32404 30728 32456 30734
rect 32404 30670 32456 30676
rect 31852 30048 31904 30054
rect 31852 29990 31904 29996
rect 30840 29504 30892 29510
rect 30840 29446 30892 29452
rect 30852 29034 30880 29446
rect 30840 29028 30892 29034
rect 30840 28970 30892 28976
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 30024 26586 30052 26862
rect 30012 26580 30064 26586
rect 30012 26522 30064 26528
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29220 24508 29516 24528
rect 29276 24506 29300 24508
rect 29356 24506 29380 24508
rect 29436 24506 29460 24508
rect 29298 24454 29300 24506
rect 29362 24454 29374 24506
rect 29436 24454 29438 24506
rect 29276 24452 29300 24454
rect 29356 24452 29380 24454
rect 29436 24452 29460 24454
rect 29220 24432 29516 24452
rect 29220 23420 29516 23440
rect 29276 23418 29300 23420
rect 29356 23418 29380 23420
rect 29436 23418 29460 23420
rect 29298 23366 29300 23418
rect 29362 23366 29374 23418
rect 29436 23366 29438 23418
rect 29276 23364 29300 23366
rect 29356 23364 29380 23366
rect 29436 23364 29460 23366
rect 29220 23344 29516 23364
rect 29220 22332 29516 22352
rect 29276 22330 29300 22332
rect 29356 22330 29380 22332
rect 29436 22330 29460 22332
rect 29298 22278 29300 22330
rect 29362 22278 29374 22330
rect 29436 22278 29438 22330
rect 29276 22276 29300 22278
rect 29356 22276 29380 22278
rect 29436 22276 29460 22278
rect 29220 22256 29516 22276
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29220 21244 29516 21264
rect 29276 21242 29300 21244
rect 29356 21242 29380 21244
rect 29436 21242 29460 21244
rect 29298 21190 29300 21242
rect 29362 21190 29374 21242
rect 29436 21190 29438 21242
rect 29276 21188 29300 21190
rect 29356 21188 29380 21190
rect 29436 21188 29460 21190
rect 29220 21168 29516 21188
rect 29220 20156 29516 20176
rect 29276 20154 29300 20156
rect 29356 20154 29380 20156
rect 29436 20154 29460 20156
rect 29298 20102 29300 20154
rect 29362 20102 29374 20154
rect 29436 20102 29438 20154
rect 29276 20100 29300 20102
rect 29356 20100 29380 20102
rect 29436 20100 29460 20102
rect 29220 20080 29516 20100
rect 29564 19718 29592 21830
rect 29748 19922 29776 24550
rect 30852 19990 30880 28970
rect 31864 28762 31892 29990
rect 31852 28756 31904 28762
rect 31852 28698 31904 28704
rect 31864 28082 31892 28698
rect 31576 28076 31628 28082
rect 31576 28018 31628 28024
rect 31852 28076 31904 28082
rect 31852 28018 31904 28024
rect 31588 27878 31616 28018
rect 31760 28008 31812 28014
rect 31760 27950 31812 27956
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 31484 27872 31536 27878
rect 31484 27814 31536 27820
rect 31576 27872 31628 27878
rect 31576 27814 31628 27820
rect 30944 27674 30972 27814
rect 30932 27668 30984 27674
rect 30932 27610 30984 27616
rect 30840 19984 30892 19990
rect 30840 19926 30892 19932
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29564 17270 29592 19654
rect 29552 17264 29604 17270
rect 29552 17206 29604 17212
rect 29564 16998 29592 17206
rect 31496 17066 31524 27814
rect 31772 27470 31800 27950
rect 31864 27674 31892 28018
rect 31852 27668 31904 27674
rect 31852 27610 31904 27616
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31760 26784 31812 26790
rect 31760 26726 31812 26732
rect 31772 23798 31800 26726
rect 32416 26586 32444 30670
rect 33152 30598 33180 33050
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 32680 28552 32732 28558
rect 32680 28494 32732 28500
rect 32692 28218 32720 28494
rect 32680 28212 32732 28218
rect 32680 28154 32732 28160
rect 32772 27668 32824 27674
rect 32772 27610 32824 27616
rect 32680 26784 32732 26790
rect 32680 26726 32732 26732
rect 32404 26580 32456 26586
rect 32404 26522 32456 26528
rect 31760 23792 31812 23798
rect 31760 23734 31812 23740
rect 31576 19984 31628 19990
rect 31576 19926 31628 19932
rect 31484 17060 31536 17066
rect 31484 17002 31536 17008
rect 29552 16992 29604 16998
rect 29552 16934 29604 16940
rect 24964 16546 25084 16574
rect 27712 16584 27764 16590
rect 24964 14278 24992 16546
rect 31588 16574 31616 19926
rect 31772 19854 31800 23734
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 32692 17610 32720 26726
rect 32312 17604 32364 17610
rect 32312 17546 32364 17552
rect 32680 17604 32732 17610
rect 32680 17546 32732 17552
rect 32324 16658 32352 17546
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32784 16574 32812 27610
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 33060 27062 33088 27406
rect 33152 27130 33180 30534
rect 33244 28218 33272 38762
rect 33520 31754 33548 38830
rect 34220 38108 34516 38128
rect 34276 38106 34300 38108
rect 34356 38106 34380 38108
rect 34436 38106 34460 38108
rect 34298 38054 34300 38106
rect 34362 38054 34374 38106
rect 34436 38054 34438 38106
rect 34276 38052 34300 38054
rect 34356 38052 34380 38054
rect 34436 38052 34460 38054
rect 34220 38032 34516 38052
rect 34220 37020 34516 37040
rect 34276 37018 34300 37020
rect 34356 37018 34380 37020
rect 34436 37018 34460 37020
rect 34298 36966 34300 37018
rect 34362 36966 34374 37018
rect 34436 36966 34438 37018
rect 34276 36964 34300 36966
rect 34356 36964 34380 36966
rect 34436 36964 34460 36966
rect 34220 36944 34516 36964
rect 35072 36372 35124 36378
rect 35072 36314 35124 36320
rect 34220 35932 34516 35952
rect 34276 35930 34300 35932
rect 34356 35930 34380 35932
rect 34436 35930 34460 35932
rect 34298 35878 34300 35930
rect 34362 35878 34374 35930
rect 34436 35878 34438 35930
rect 34276 35876 34300 35878
rect 34356 35876 34380 35878
rect 34436 35876 34460 35878
rect 34220 35856 34516 35876
rect 34220 34844 34516 34864
rect 34276 34842 34300 34844
rect 34356 34842 34380 34844
rect 34436 34842 34460 34844
rect 34298 34790 34300 34842
rect 34362 34790 34374 34842
rect 34436 34790 34438 34842
rect 34276 34788 34300 34790
rect 34356 34788 34380 34790
rect 34436 34788 34460 34790
rect 34220 34768 34516 34788
rect 34220 33756 34516 33776
rect 34276 33754 34300 33756
rect 34356 33754 34380 33756
rect 34436 33754 34460 33756
rect 34298 33702 34300 33754
rect 34362 33702 34374 33754
rect 34436 33702 34438 33754
rect 34276 33700 34300 33702
rect 34356 33700 34380 33702
rect 34436 33700 34460 33702
rect 34220 33680 34516 33700
rect 34220 32668 34516 32688
rect 34276 32666 34300 32668
rect 34356 32666 34380 32668
rect 34436 32666 34460 32668
rect 34298 32614 34300 32666
rect 34362 32614 34374 32666
rect 34436 32614 34438 32666
rect 34276 32612 34300 32614
rect 34356 32612 34380 32614
rect 34436 32612 34460 32614
rect 34220 32592 34516 32612
rect 33520 31726 33824 31754
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33520 29850 33548 30194
rect 33508 29844 33560 29850
rect 33508 29786 33560 29792
rect 33796 29510 33824 31726
rect 34220 31580 34516 31600
rect 34276 31578 34300 31580
rect 34356 31578 34380 31580
rect 34436 31578 34460 31580
rect 34298 31526 34300 31578
rect 34362 31526 34374 31578
rect 34436 31526 34438 31578
rect 34276 31524 34300 31526
rect 34356 31524 34380 31526
rect 34436 31524 34460 31526
rect 34220 31504 34516 31524
rect 34220 30492 34516 30512
rect 34276 30490 34300 30492
rect 34356 30490 34380 30492
rect 34436 30490 34460 30492
rect 34298 30438 34300 30490
rect 34362 30438 34374 30490
rect 34436 30438 34438 30490
rect 34276 30436 34300 30438
rect 34356 30436 34380 30438
rect 34436 30436 34460 30438
rect 34220 30416 34516 30436
rect 35084 30326 35112 36314
rect 35360 30326 35388 39578
rect 38948 37330 38976 42570
rect 39220 41916 39516 41936
rect 39276 41914 39300 41916
rect 39356 41914 39380 41916
rect 39436 41914 39460 41916
rect 39298 41862 39300 41914
rect 39362 41862 39374 41914
rect 39436 41862 39438 41914
rect 39276 41860 39300 41862
rect 39356 41860 39380 41862
rect 39436 41860 39460 41862
rect 39220 41840 39516 41860
rect 39684 41750 39712 42706
rect 42812 42566 42840 42706
rect 43352 42696 43404 42702
rect 43352 42638 43404 42644
rect 43260 42628 43312 42634
rect 43260 42570 43312 42576
rect 42800 42560 42852 42566
rect 42800 42502 42852 42508
rect 40684 42016 40736 42022
rect 40684 41958 40736 41964
rect 39672 41744 39724 41750
rect 39672 41686 39724 41692
rect 39220 40828 39516 40848
rect 39276 40826 39300 40828
rect 39356 40826 39380 40828
rect 39436 40826 39460 40828
rect 39298 40774 39300 40826
rect 39362 40774 39374 40826
rect 39436 40774 39438 40826
rect 39276 40772 39300 40774
rect 39356 40772 39380 40774
rect 39436 40772 39460 40774
rect 39220 40752 39516 40772
rect 39220 39740 39516 39760
rect 39276 39738 39300 39740
rect 39356 39738 39380 39740
rect 39436 39738 39460 39740
rect 39298 39686 39300 39738
rect 39362 39686 39374 39738
rect 39436 39686 39438 39738
rect 39276 39684 39300 39686
rect 39356 39684 39380 39686
rect 39436 39684 39460 39686
rect 39220 39664 39516 39684
rect 39672 39092 39724 39098
rect 39672 39034 39724 39040
rect 39220 38652 39516 38672
rect 39276 38650 39300 38652
rect 39356 38650 39380 38652
rect 39436 38650 39460 38652
rect 39298 38598 39300 38650
rect 39362 38598 39374 38650
rect 39436 38598 39438 38650
rect 39276 38596 39300 38598
rect 39356 38596 39380 38598
rect 39436 38596 39460 38598
rect 39220 38576 39516 38596
rect 39120 37664 39172 37670
rect 39120 37606 39172 37612
rect 38936 37324 38988 37330
rect 38936 37266 38988 37272
rect 38200 33856 38252 33862
rect 38200 33798 38252 33804
rect 38212 33386 38240 33798
rect 38200 33380 38252 33386
rect 38200 33322 38252 33328
rect 38292 33312 38344 33318
rect 38292 33254 38344 33260
rect 38016 32904 38068 32910
rect 38016 32846 38068 32852
rect 38028 32230 38056 32846
rect 37280 32224 37332 32230
rect 37280 32166 37332 32172
rect 38016 32224 38068 32230
rect 38016 32166 38068 32172
rect 37292 31754 37320 32166
rect 38304 31822 38332 33254
rect 38476 32972 38528 32978
rect 38476 32914 38528 32920
rect 38488 32774 38516 32914
rect 38476 32768 38528 32774
rect 38476 32710 38528 32716
rect 38752 32360 38804 32366
rect 38752 32302 38804 32308
rect 38764 32230 38792 32302
rect 38660 32224 38712 32230
rect 38660 32166 38712 32172
rect 38752 32224 38804 32230
rect 38752 32166 38804 32172
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 37292 31726 37596 31754
rect 37464 30932 37516 30938
rect 37464 30874 37516 30880
rect 35072 30320 35124 30326
rect 35072 30262 35124 30268
rect 35348 30320 35400 30326
rect 35348 30262 35400 30268
rect 33784 29504 33836 29510
rect 33784 29446 33836 29452
rect 33232 28212 33284 28218
rect 33232 28154 33284 28160
rect 33244 28082 33272 28154
rect 33232 28076 33284 28082
rect 33232 28018 33284 28024
rect 33140 27124 33192 27130
rect 33140 27066 33192 27072
rect 33048 27056 33100 27062
rect 33048 26998 33100 27004
rect 33796 19922 33824 29446
rect 34220 29404 34516 29424
rect 34276 29402 34300 29404
rect 34356 29402 34380 29404
rect 34436 29402 34460 29404
rect 34298 29350 34300 29402
rect 34362 29350 34374 29402
rect 34436 29350 34438 29402
rect 34276 29348 34300 29350
rect 34356 29348 34380 29350
rect 34436 29348 34460 29350
rect 34220 29328 34516 29348
rect 34220 28316 34516 28336
rect 34276 28314 34300 28316
rect 34356 28314 34380 28316
rect 34436 28314 34460 28316
rect 34298 28262 34300 28314
rect 34362 28262 34374 28314
rect 34436 28262 34438 28314
rect 34276 28260 34300 28262
rect 34356 28260 34380 28262
rect 34436 28260 34460 28262
rect 34220 28240 34516 28260
rect 34220 27228 34516 27248
rect 34276 27226 34300 27228
rect 34356 27226 34380 27228
rect 34436 27226 34460 27228
rect 34298 27174 34300 27226
rect 34362 27174 34374 27226
rect 34436 27174 34438 27226
rect 34276 27172 34300 27174
rect 34356 27172 34380 27174
rect 34436 27172 34460 27174
rect 34220 27152 34516 27172
rect 34220 26140 34516 26160
rect 34276 26138 34300 26140
rect 34356 26138 34380 26140
rect 34436 26138 34460 26140
rect 34298 26086 34300 26138
rect 34362 26086 34374 26138
rect 34436 26086 34438 26138
rect 34276 26084 34300 26086
rect 34356 26084 34380 26086
rect 34436 26084 34460 26086
rect 34220 26064 34516 26084
rect 34220 25052 34516 25072
rect 34276 25050 34300 25052
rect 34356 25050 34380 25052
rect 34436 25050 34460 25052
rect 34298 24998 34300 25050
rect 34362 24998 34374 25050
rect 34436 24998 34438 25050
rect 34276 24996 34300 24998
rect 34356 24996 34380 24998
rect 34436 24996 34460 24998
rect 34220 24976 34516 24996
rect 34220 23964 34516 23984
rect 34276 23962 34300 23964
rect 34356 23962 34380 23964
rect 34436 23962 34460 23964
rect 34298 23910 34300 23962
rect 34362 23910 34374 23962
rect 34436 23910 34438 23962
rect 34276 23908 34300 23910
rect 34356 23908 34380 23910
rect 34436 23908 34460 23910
rect 34220 23888 34516 23908
rect 34220 22876 34516 22896
rect 34276 22874 34300 22876
rect 34356 22874 34380 22876
rect 34436 22874 34460 22876
rect 34298 22822 34300 22874
rect 34362 22822 34374 22874
rect 34436 22822 34438 22874
rect 34276 22820 34300 22822
rect 34356 22820 34380 22822
rect 34436 22820 34460 22822
rect 34220 22800 34516 22820
rect 34220 21788 34516 21808
rect 34276 21786 34300 21788
rect 34356 21786 34380 21788
rect 34436 21786 34460 21788
rect 34298 21734 34300 21786
rect 34362 21734 34374 21786
rect 34436 21734 34438 21786
rect 34276 21732 34300 21734
rect 34356 21732 34380 21734
rect 34436 21732 34460 21734
rect 34220 21712 34516 21732
rect 34220 20700 34516 20720
rect 34276 20698 34300 20700
rect 34356 20698 34380 20700
rect 34436 20698 34460 20700
rect 34298 20646 34300 20698
rect 34362 20646 34374 20698
rect 34436 20646 34438 20698
rect 34276 20644 34300 20646
rect 34356 20644 34380 20646
rect 34436 20644 34460 20646
rect 34220 20624 34516 20644
rect 33784 19916 33836 19922
rect 33784 19858 33836 19864
rect 33796 16574 33824 19858
rect 34220 19612 34516 19632
rect 34276 19610 34300 19612
rect 34356 19610 34380 19612
rect 34436 19610 34460 19612
rect 34298 19558 34300 19610
rect 34362 19558 34374 19610
rect 34436 19558 34438 19610
rect 34276 19556 34300 19558
rect 34356 19556 34380 19558
rect 34436 19556 34460 19558
rect 34220 19536 34516 19556
rect 31588 16546 31708 16574
rect 32784 16546 32996 16574
rect 33796 16546 33916 16574
rect 27712 16526 27764 16532
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 31680 13462 31708 16546
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 31668 13456 31720 13462
rect 31668 13398 31720 13404
rect 32600 13124 32628 15642
rect 32864 9376 32916 9382
rect 32864 9318 32916 9324
rect 32876 9194 32904 9318
rect 32614 9166 32904 9194
rect 32864 6112 32916 6118
rect 24950 6080 25006 6089
rect 32968 6089 32996 16546
rect 32864 6054 32916 6060
rect 32954 6080 33010 6089
rect 24950 6015 25006 6024
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 24964 5710 24992 6015
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 23756 5296 23808 5302
rect 32876 5250 32904 6054
rect 32954 6015 33010 6024
rect 23808 5244 24058 5250
rect 23756 5238 24058 5244
rect 23768 5222 24058 5238
rect 32614 5222 32904 5250
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 9220 2748 9516 2768
rect 9276 2746 9300 2748
rect 9356 2746 9380 2748
rect 9436 2746 9460 2748
rect 9298 2694 9300 2746
rect 9362 2694 9374 2746
rect 9436 2694 9438 2746
rect 9276 2692 9300 2694
rect 9356 2692 9380 2694
rect 9436 2692 9460 2694
rect 9220 2672 9516 2692
rect 10888 2650 10916 2926
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 1398 2544 1454 2553
rect 1398 2479 1400 2488
rect 1452 2479 1454 2488
rect 1400 2450 1452 2456
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 12452 800 12480 3470
rect 14220 3292 14516 3312
rect 14276 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14298 3238 14300 3290
rect 14362 3238 14374 3290
rect 14436 3238 14438 3290
rect 14276 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14220 3216 14516 3236
rect 32968 3126 32996 6015
rect 33888 5778 33916 16546
rect 34612 8084 34664 8090
rect 34612 8026 34664 8032
rect 34624 6361 34652 8026
rect 35360 6914 35388 30262
rect 35624 30184 35676 30190
rect 35624 30126 35676 30132
rect 35636 29510 35664 30126
rect 35624 29504 35676 29510
rect 35624 29446 35676 29452
rect 37280 29504 37332 29510
rect 37280 29446 37332 29452
rect 35636 29102 35664 29446
rect 35624 29096 35676 29102
rect 35624 29038 35676 29044
rect 37292 27130 37320 29446
rect 37372 28552 37424 28558
rect 37372 28494 37424 28500
rect 37280 27124 37332 27130
rect 37280 27066 37332 27072
rect 37384 25430 37412 28494
rect 37372 25424 37424 25430
rect 37372 25366 37424 25372
rect 35716 24268 35768 24274
rect 35716 24210 35768 24216
rect 35728 23798 35756 24210
rect 35716 23792 35768 23798
rect 35716 23734 35768 23740
rect 37280 9104 37332 9110
rect 37280 9046 37332 9052
rect 35268 6886 35388 6914
rect 34610 6352 34666 6361
rect 34610 6287 34666 6296
rect 33876 5772 33928 5778
rect 33876 5714 33928 5720
rect 35268 5030 35296 6886
rect 37292 5953 37320 9046
rect 37476 8022 37504 30874
rect 37568 29646 37596 31726
rect 37556 29640 37608 29646
rect 37556 29582 37608 29588
rect 37568 24342 37596 29582
rect 38108 28552 38160 28558
rect 38108 28494 38160 28500
rect 38120 28422 38148 28494
rect 38016 28416 38068 28422
rect 38016 28358 38068 28364
rect 38108 28416 38160 28422
rect 38108 28358 38160 28364
rect 38028 28234 38056 28358
rect 38028 28206 38148 28234
rect 37740 26784 37792 26790
rect 37740 26726 37792 26732
rect 37556 24336 37608 24342
rect 37556 24278 37608 24284
rect 37648 18624 37700 18630
rect 37648 18566 37700 18572
rect 37464 8016 37516 8022
rect 37464 7958 37516 7964
rect 37278 5944 37334 5953
rect 37660 5914 37688 18566
rect 37752 11286 37780 26726
rect 38016 25424 38068 25430
rect 38016 25366 38068 25372
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 37740 11280 37792 11286
rect 37740 11222 37792 11228
rect 37752 10810 37780 11222
rect 37740 10804 37792 10810
rect 37740 10746 37792 10752
rect 37278 5879 37334 5888
rect 37648 5908 37700 5914
rect 37292 5234 37320 5879
rect 37648 5850 37700 5856
rect 37280 5228 37332 5234
rect 37280 5170 37332 5176
rect 35256 5024 35308 5030
rect 35256 4966 35308 4972
rect 35268 3534 35296 4966
rect 35256 3528 35308 3534
rect 35256 3470 35308 3476
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 37844 2650 37872 16594
rect 37924 11144 37976 11150
rect 37922 11112 37924 11121
rect 37976 11112 37978 11121
rect 37922 11047 37978 11056
rect 38028 6458 38056 25366
rect 38120 8022 38148 28206
rect 38304 13258 38332 31758
rect 38672 31754 38700 32166
rect 38948 31890 38976 37266
rect 39028 34536 39080 34542
rect 39028 34478 39080 34484
rect 38936 31884 38988 31890
rect 38936 31826 38988 31832
rect 38660 31748 38712 31754
rect 38660 31690 38712 31696
rect 38948 31482 38976 31826
rect 38936 31476 38988 31482
rect 38936 31418 38988 31424
rect 38384 31408 38436 31414
rect 38384 31350 38436 31356
rect 38396 30734 38424 31350
rect 38384 30728 38436 30734
rect 38384 30670 38436 30676
rect 38396 28762 38424 30670
rect 38384 28756 38436 28762
rect 38384 28698 38436 28704
rect 38396 28558 38424 28698
rect 38384 28552 38436 28558
rect 38384 28494 38436 28500
rect 38568 28416 38620 28422
rect 38568 28358 38620 28364
rect 38292 13252 38344 13258
rect 38292 13194 38344 13200
rect 38304 8634 38332 13194
rect 38292 8628 38344 8634
rect 38292 8570 38344 8576
rect 38476 8628 38528 8634
rect 38476 8570 38528 8576
rect 38304 8090 38332 8570
rect 38292 8084 38344 8090
rect 38292 8026 38344 8032
rect 38108 8016 38160 8022
rect 38108 7958 38160 7964
rect 38120 7546 38148 7958
rect 38304 7546 38332 8026
rect 38108 7540 38160 7546
rect 38108 7482 38160 7488
rect 38292 7540 38344 7546
rect 38292 7482 38344 7488
rect 38016 6452 38068 6458
rect 38016 6394 38068 6400
rect 38028 5166 38056 6394
rect 38120 5166 38148 7482
rect 38488 6118 38516 8570
rect 38476 6112 38528 6118
rect 38476 6054 38528 6060
rect 38580 5370 38608 28358
rect 39040 27962 39068 34478
rect 39132 31958 39160 37606
rect 39220 37564 39516 37584
rect 39276 37562 39300 37564
rect 39356 37562 39380 37564
rect 39436 37562 39460 37564
rect 39298 37510 39300 37562
rect 39362 37510 39374 37562
rect 39436 37510 39438 37562
rect 39276 37508 39300 37510
rect 39356 37508 39380 37510
rect 39436 37508 39460 37510
rect 39220 37488 39516 37508
rect 39220 36476 39516 36496
rect 39276 36474 39300 36476
rect 39356 36474 39380 36476
rect 39436 36474 39460 36476
rect 39298 36422 39300 36474
rect 39362 36422 39374 36474
rect 39436 36422 39438 36474
rect 39276 36420 39300 36422
rect 39356 36420 39380 36422
rect 39436 36420 39460 36422
rect 39220 36400 39516 36420
rect 39684 35494 39712 39034
rect 39672 35488 39724 35494
rect 39672 35430 39724 35436
rect 39220 35388 39516 35408
rect 39276 35386 39300 35388
rect 39356 35386 39380 35388
rect 39436 35386 39460 35388
rect 39298 35334 39300 35386
rect 39362 35334 39374 35386
rect 39436 35334 39438 35386
rect 39276 35332 39300 35334
rect 39356 35332 39380 35334
rect 39436 35332 39460 35334
rect 39220 35312 39516 35332
rect 39684 34542 39712 35430
rect 39672 34536 39724 34542
rect 39672 34478 39724 34484
rect 39220 34300 39516 34320
rect 39276 34298 39300 34300
rect 39356 34298 39380 34300
rect 39436 34298 39460 34300
rect 39298 34246 39300 34298
rect 39362 34246 39374 34298
rect 39436 34246 39438 34298
rect 39276 34244 39300 34246
rect 39356 34244 39380 34246
rect 39436 34244 39460 34246
rect 39220 34224 39516 34244
rect 39672 33516 39724 33522
rect 39672 33458 39724 33464
rect 39684 33318 39712 33458
rect 39580 33312 39632 33318
rect 39580 33254 39632 33260
rect 39672 33312 39724 33318
rect 39672 33254 39724 33260
rect 39220 33212 39516 33232
rect 39276 33210 39300 33212
rect 39356 33210 39380 33212
rect 39436 33210 39460 33212
rect 39298 33158 39300 33210
rect 39362 33158 39374 33210
rect 39436 33158 39438 33210
rect 39276 33156 39300 33158
rect 39356 33156 39380 33158
rect 39436 33156 39460 33158
rect 39220 33136 39516 33156
rect 39220 32124 39516 32144
rect 39276 32122 39300 32124
rect 39356 32122 39380 32124
rect 39436 32122 39460 32124
rect 39298 32070 39300 32122
rect 39362 32070 39374 32122
rect 39436 32070 39438 32122
rect 39276 32068 39300 32070
rect 39356 32068 39380 32070
rect 39436 32068 39460 32070
rect 39220 32048 39516 32068
rect 39120 31952 39172 31958
rect 39120 31894 39172 31900
rect 39120 31816 39172 31822
rect 39120 31758 39172 31764
rect 39132 31210 39160 31758
rect 39592 31498 39620 33254
rect 39684 31754 39712 33254
rect 39764 32904 39816 32910
rect 39764 32846 39816 32852
rect 39672 31748 39724 31754
rect 39672 31690 39724 31696
rect 39592 31470 39712 31498
rect 39120 31204 39172 31210
rect 39120 31146 39172 31152
rect 38764 27934 39068 27962
rect 38764 11354 38792 27934
rect 38936 27872 38988 27878
rect 38936 27814 38988 27820
rect 38948 26738 38976 27814
rect 38948 26710 39068 26738
rect 38936 24812 38988 24818
rect 38936 24754 38988 24760
rect 38752 11348 38804 11354
rect 38752 11290 38804 11296
rect 38948 6914 38976 24754
rect 39040 7546 39068 26710
rect 39132 12986 39160 31146
rect 39220 31036 39516 31056
rect 39276 31034 39300 31036
rect 39356 31034 39380 31036
rect 39436 31034 39460 31036
rect 39298 30982 39300 31034
rect 39362 30982 39374 31034
rect 39436 30982 39438 31034
rect 39276 30980 39300 30982
rect 39356 30980 39380 30982
rect 39436 30980 39460 30982
rect 39220 30960 39516 30980
rect 39580 30252 39632 30258
rect 39580 30194 39632 30200
rect 39220 29948 39516 29968
rect 39276 29946 39300 29948
rect 39356 29946 39380 29948
rect 39436 29946 39460 29948
rect 39298 29894 39300 29946
rect 39362 29894 39374 29946
rect 39436 29894 39438 29946
rect 39276 29892 39300 29894
rect 39356 29892 39380 29894
rect 39436 29892 39460 29894
rect 39220 29872 39516 29892
rect 39592 29034 39620 30194
rect 39580 29028 39632 29034
rect 39580 28970 39632 28976
rect 39220 28860 39516 28880
rect 39276 28858 39300 28860
rect 39356 28858 39380 28860
rect 39436 28858 39460 28860
rect 39298 28806 39300 28858
rect 39362 28806 39374 28858
rect 39436 28806 39438 28858
rect 39276 28804 39300 28806
rect 39356 28804 39380 28806
rect 39436 28804 39460 28806
rect 39220 28784 39516 28804
rect 39220 27772 39516 27792
rect 39276 27770 39300 27772
rect 39356 27770 39380 27772
rect 39436 27770 39460 27772
rect 39298 27718 39300 27770
rect 39362 27718 39374 27770
rect 39436 27718 39438 27770
rect 39276 27716 39300 27718
rect 39356 27716 39380 27718
rect 39436 27716 39460 27718
rect 39220 27696 39516 27716
rect 39220 26684 39516 26704
rect 39276 26682 39300 26684
rect 39356 26682 39380 26684
rect 39436 26682 39460 26684
rect 39298 26630 39300 26682
rect 39362 26630 39374 26682
rect 39436 26630 39438 26682
rect 39276 26628 39300 26630
rect 39356 26628 39380 26630
rect 39436 26628 39460 26630
rect 39220 26608 39516 26628
rect 39220 25596 39516 25616
rect 39276 25594 39300 25596
rect 39356 25594 39380 25596
rect 39436 25594 39460 25596
rect 39298 25542 39300 25594
rect 39362 25542 39374 25594
rect 39436 25542 39438 25594
rect 39276 25540 39300 25542
rect 39356 25540 39380 25542
rect 39436 25540 39460 25542
rect 39220 25520 39516 25540
rect 39592 25378 39620 28970
rect 39500 25350 39620 25378
rect 39500 24682 39528 25350
rect 39684 24834 39712 31470
rect 39776 30258 39804 32846
rect 40500 32768 40552 32774
rect 40500 32710 40552 32716
rect 39948 32224 40000 32230
rect 39948 32166 40000 32172
rect 39856 31884 39908 31890
rect 39856 31826 39908 31832
rect 39764 30252 39816 30258
rect 39764 30194 39816 30200
rect 39868 30138 39896 31826
rect 39776 30110 39896 30138
rect 39776 24886 39804 30110
rect 39856 30048 39908 30054
rect 39856 29990 39908 29996
rect 39592 24806 39712 24834
rect 39764 24880 39816 24886
rect 39764 24822 39816 24828
rect 39488 24676 39540 24682
rect 39488 24618 39540 24624
rect 39220 24508 39516 24528
rect 39276 24506 39300 24508
rect 39356 24506 39380 24508
rect 39436 24506 39460 24508
rect 39298 24454 39300 24506
rect 39362 24454 39374 24506
rect 39436 24454 39438 24506
rect 39276 24452 39300 24454
rect 39356 24452 39380 24454
rect 39436 24452 39460 24454
rect 39220 24432 39516 24452
rect 39220 23420 39516 23440
rect 39276 23418 39300 23420
rect 39356 23418 39380 23420
rect 39436 23418 39460 23420
rect 39298 23366 39300 23418
rect 39362 23366 39374 23418
rect 39436 23366 39438 23418
rect 39276 23364 39300 23366
rect 39356 23364 39380 23366
rect 39436 23364 39460 23366
rect 39220 23344 39516 23364
rect 39592 22982 39620 24806
rect 39868 24750 39896 29990
rect 39672 24744 39724 24750
rect 39672 24686 39724 24692
rect 39856 24744 39908 24750
rect 39856 24686 39908 24692
rect 39580 22976 39632 22982
rect 39580 22918 39632 22924
rect 39220 22332 39516 22352
rect 39276 22330 39300 22332
rect 39356 22330 39380 22332
rect 39436 22330 39460 22332
rect 39298 22278 39300 22330
rect 39362 22278 39374 22330
rect 39436 22278 39438 22330
rect 39276 22276 39300 22278
rect 39356 22276 39380 22278
rect 39436 22276 39460 22278
rect 39220 22256 39516 22276
rect 39220 21244 39516 21264
rect 39276 21242 39300 21244
rect 39356 21242 39380 21244
rect 39436 21242 39460 21244
rect 39298 21190 39300 21242
rect 39362 21190 39374 21242
rect 39436 21190 39438 21242
rect 39276 21188 39300 21190
rect 39356 21188 39380 21190
rect 39436 21188 39460 21190
rect 39220 21168 39516 21188
rect 39220 20156 39516 20176
rect 39276 20154 39300 20156
rect 39356 20154 39380 20156
rect 39436 20154 39460 20156
rect 39298 20102 39300 20154
rect 39362 20102 39374 20154
rect 39436 20102 39438 20154
rect 39276 20100 39300 20102
rect 39356 20100 39380 20102
rect 39436 20100 39460 20102
rect 39220 20080 39516 20100
rect 39220 19068 39516 19088
rect 39276 19066 39300 19068
rect 39356 19066 39380 19068
rect 39436 19066 39460 19068
rect 39298 19014 39300 19066
rect 39362 19014 39374 19066
rect 39436 19014 39438 19066
rect 39276 19012 39300 19014
rect 39356 19012 39380 19014
rect 39436 19012 39460 19014
rect 39220 18992 39516 19012
rect 39220 17980 39516 18000
rect 39276 17978 39300 17980
rect 39356 17978 39380 17980
rect 39436 17978 39460 17980
rect 39298 17926 39300 17978
rect 39362 17926 39374 17978
rect 39436 17926 39438 17978
rect 39276 17924 39300 17926
rect 39356 17924 39380 17926
rect 39436 17924 39460 17926
rect 39220 17904 39516 17924
rect 39220 16892 39516 16912
rect 39276 16890 39300 16892
rect 39356 16890 39380 16892
rect 39436 16890 39460 16892
rect 39298 16838 39300 16890
rect 39362 16838 39374 16890
rect 39436 16838 39438 16890
rect 39276 16836 39300 16838
rect 39356 16836 39380 16838
rect 39436 16836 39460 16838
rect 39220 16816 39516 16836
rect 39220 15804 39516 15824
rect 39276 15802 39300 15804
rect 39356 15802 39380 15804
rect 39436 15802 39460 15804
rect 39298 15750 39300 15802
rect 39362 15750 39374 15802
rect 39436 15750 39438 15802
rect 39276 15748 39300 15750
rect 39356 15748 39380 15750
rect 39436 15748 39460 15750
rect 39220 15728 39516 15748
rect 39592 15638 39620 22918
rect 39684 17678 39712 24686
rect 39672 17672 39724 17678
rect 39672 17614 39724 17620
rect 39672 17196 39724 17202
rect 39672 17138 39724 17144
rect 39684 16574 39712 17138
rect 39684 16546 39804 16574
rect 39580 15632 39632 15638
rect 39580 15574 39632 15580
rect 39220 14716 39516 14736
rect 39276 14714 39300 14716
rect 39356 14714 39380 14716
rect 39436 14714 39460 14716
rect 39298 14662 39300 14714
rect 39362 14662 39374 14714
rect 39436 14662 39438 14714
rect 39276 14660 39300 14662
rect 39356 14660 39380 14662
rect 39436 14660 39460 14662
rect 39220 14640 39516 14660
rect 39220 13628 39516 13648
rect 39276 13626 39300 13628
rect 39356 13626 39380 13628
rect 39436 13626 39460 13628
rect 39298 13574 39300 13626
rect 39362 13574 39374 13626
rect 39436 13574 39438 13626
rect 39276 13572 39300 13574
rect 39356 13572 39380 13574
rect 39436 13572 39460 13574
rect 39220 13552 39516 13572
rect 39120 12980 39172 12986
rect 39120 12922 39172 12928
rect 39132 8022 39160 12922
rect 39220 12540 39516 12560
rect 39276 12538 39300 12540
rect 39356 12538 39380 12540
rect 39436 12538 39460 12540
rect 39298 12486 39300 12538
rect 39362 12486 39374 12538
rect 39436 12486 39438 12538
rect 39276 12484 39300 12486
rect 39356 12484 39380 12486
rect 39436 12484 39460 12486
rect 39220 12464 39516 12484
rect 39220 11452 39516 11472
rect 39276 11450 39300 11452
rect 39356 11450 39380 11452
rect 39436 11450 39460 11452
rect 39298 11398 39300 11450
rect 39362 11398 39374 11450
rect 39436 11398 39438 11450
rect 39276 11396 39300 11398
rect 39356 11396 39380 11398
rect 39436 11396 39460 11398
rect 39220 11376 39516 11396
rect 39220 10364 39516 10384
rect 39276 10362 39300 10364
rect 39356 10362 39380 10364
rect 39436 10362 39460 10364
rect 39298 10310 39300 10362
rect 39362 10310 39374 10362
rect 39436 10310 39438 10362
rect 39276 10308 39300 10310
rect 39356 10308 39380 10310
rect 39436 10308 39460 10310
rect 39220 10288 39516 10308
rect 39220 9276 39516 9296
rect 39276 9274 39300 9276
rect 39356 9274 39380 9276
rect 39436 9274 39460 9276
rect 39298 9222 39300 9274
rect 39362 9222 39374 9274
rect 39436 9222 39438 9274
rect 39276 9220 39300 9222
rect 39356 9220 39380 9222
rect 39436 9220 39460 9222
rect 39220 9200 39516 9220
rect 39220 8188 39516 8208
rect 39276 8186 39300 8188
rect 39356 8186 39380 8188
rect 39436 8186 39460 8188
rect 39298 8134 39300 8186
rect 39362 8134 39374 8186
rect 39436 8134 39438 8186
rect 39276 8132 39300 8134
rect 39356 8132 39380 8134
rect 39436 8132 39460 8134
rect 39220 8112 39516 8132
rect 39120 8016 39172 8022
rect 39120 7958 39172 7964
rect 39028 7540 39080 7546
rect 39028 7482 39080 7488
rect 39132 7206 39160 7958
rect 39776 7478 39804 16546
rect 39960 8090 39988 32166
rect 40512 17338 40540 32710
rect 40696 32434 40724 41958
rect 42064 37936 42116 37942
rect 42064 37878 42116 37884
rect 40776 36032 40828 36038
rect 40776 35974 40828 35980
rect 40684 32428 40736 32434
rect 40684 32370 40736 32376
rect 40696 31414 40724 32370
rect 40684 31408 40736 31414
rect 40684 31350 40736 31356
rect 40500 17332 40552 17338
rect 40500 17274 40552 17280
rect 40788 15502 40816 35974
rect 41052 32020 41104 32026
rect 41052 31962 41104 31968
rect 40776 15496 40828 15502
rect 40776 15438 40828 15444
rect 40788 15162 40816 15438
rect 40776 15156 40828 15162
rect 40776 15098 40828 15104
rect 39948 8084 40000 8090
rect 39948 8026 40000 8032
rect 39764 7472 39816 7478
rect 39684 7420 39764 7426
rect 39684 7414 39816 7420
rect 39684 7398 39804 7414
rect 39120 7200 39172 7206
rect 39120 7142 39172 7148
rect 39132 7002 39160 7142
rect 39220 7100 39516 7120
rect 39276 7098 39300 7100
rect 39356 7098 39380 7100
rect 39436 7098 39460 7100
rect 39298 7046 39300 7098
rect 39362 7046 39374 7098
rect 39436 7046 39438 7098
rect 39276 7044 39300 7046
rect 39356 7044 39380 7046
rect 39436 7044 39460 7046
rect 39220 7024 39516 7044
rect 39684 7002 39712 7398
rect 39764 7336 39816 7342
rect 39764 7278 39816 7284
rect 39776 7206 39804 7278
rect 39764 7200 39816 7206
rect 39764 7142 39816 7148
rect 39120 6996 39172 7002
rect 39120 6938 39172 6944
rect 39672 6996 39724 7002
rect 39672 6938 39724 6944
rect 38856 6886 38976 6914
rect 38568 5364 38620 5370
rect 38568 5306 38620 5312
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 38108 5160 38160 5166
rect 38108 5102 38160 5108
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 38120 4826 38148 5102
rect 38108 4820 38160 4826
rect 38108 4762 38160 4768
rect 38304 4282 38332 5102
rect 38856 5098 38884 6886
rect 39220 6012 39516 6032
rect 39276 6010 39300 6012
rect 39356 6010 39380 6012
rect 39436 6010 39460 6012
rect 39298 5958 39300 6010
rect 39362 5958 39374 6010
rect 39436 5958 39438 6010
rect 39276 5956 39300 5958
rect 39356 5956 39380 5958
rect 39436 5956 39460 5958
rect 39220 5936 39516 5956
rect 38844 5092 38896 5098
rect 38844 5034 38896 5040
rect 39028 5024 39080 5030
rect 39028 4966 39080 4972
rect 38292 4276 38344 4282
rect 38292 4218 38344 4224
rect 39040 3058 39068 4966
rect 39220 4924 39516 4944
rect 39276 4922 39300 4924
rect 39356 4922 39380 4924
rect 39436 4922 39460 4924
rect 39298 4870 39300 4922
rect 39362 4870 39374 4922
rect 39436 4870 39438 4922
rect 39276 4868 39300 4870
rect 39356 4868 39380 4870
rect 39436 4868 39460 4870
rect 39220 4848 39516 4868
rect 39220 3836 39516 3856
rect 39276 3834 39300 3836
rect 39356 3834 39380 3836
rect 39436 3834 39460 3836
rect 39298 3782 39300 3834
rect 39362 3782 39374 3834
rect 39436 3782 39438 3834
rect 39276 3780 39300 3782
rect 39356 3780 39380 3782
rect 39436 3780 39460 3782
rect 39220 3760 39516 3780
rect 41064 3738 41092 31962
rect 41236 31816 41288 31822
rect 41236 31758 41288 31764
rect 41052 3732 41104 3738
rect 41052 3674 41104 3680
rect 41248 3602 41276 31758
rect 41696 28960 41748 28966
rect 41696 28902 41748 28908
rect 41604 27056 41656 27062
rect 41604 26998 41656 27004
rect 41616 3738 41644 26998
rect 41708 17066 41736 28902
rect 42076 25702 42104 37878
rect 42708 32836 42760 32842
rect 42708 32778 42760 32784
rect 42720 29578 42748 32778
rect 42708 29572 42760 29578
rect 42708 29514 42760 29520
rect 42064 25696 42116 25702
rect 42064 25638 42116 25644
rect 42076 24886 42104 25638
rect 42064 24880 42116 24886
rect 42064 24822 42116 24828
rect 42616 24880 42668 24886
rect 42616 24822 42668 24828
rect 41696 17060 41748 17066
rect 41696 17002 41748 17008
rect 42432 15904 42484 15910
rect 42432 15846 42484 15852
rect 42444 15502 42472 15846
rect 42432 15496 42484 15502
rect 42432 15438 42484 15444
rect 42156 13932 42208 13938
rect 42156 13874 42208 13880
rect 42168 8090 42196 13874
rect 42444 11694 42472 15438
rect 42432 11688 42484 11694
rect 42432 11630 42484 11636
rect 42156 8084 42208 8090
rect 42156 8026 42208 8032
rect 42444 7886 42472 11630
rect 42628 8090 42656 24822
rect 42708 17128 42760 17134
rect 42708 17070 42760 17076
rect 42720 15910 42748 17070
rect 42708 15904 42760 15910
rect 42708 15846 42760 15852
rect 42616 8084 42668 8090
rect 42616 8026 42668 8032
rect 42432 7880 42484 7886
rect 42432 7822 42484 7828
rect 42444 7478 42472 7822
rect 42628 7546 42656 8026
rect 42616 7540 42668 7546
rect 42616 7482 42668 7488
rect 42432 7472 42484 7478
rect 42432 7414 42484 7420
rect 42340 4004 42392 4010
rect 42340 3946 42392 3952
rect 41604 3732 41656 3738
rect 41604 3674 41656 3680
rect 42352 3602 42380 3946
rect 42812 3738 42840 42502
rect 43272 30258 43300 42570
rect 43364 42022 43392 42638
rect 44220 42460 44516 42480
rect 44276 42458 44300 42460
rect 44356 42458 44380 42460
rect 44436 42458 44460 42460
rect 44298 42406 44300 42458
rect 44362 42406 44374 42458
rect 44436 42406 44438 42458
rect 44276 42404 44300 42406
rect 44356 42404 44380 42406
rect 44436 42404 44460 42406
rect 44220 42384 44516 42404
rect 43352 42016 43404 42022
rect 43352 41958 43404 41964
rect 48134 41712 48190 41721
rect 48134 41647 48136 41656
rect 48188 41647 48190 41656
rect 48136 41618 48188 41624
rect 44548 41472 44600 41478
rect 44548 41414 44600 41420
rect 44220 41372 44516 41392
rect 44276 41370 44300 41372
rect 44356 41370 44380 41372
rect 44436 41370 44460 41372
rect 44298 41318 44300 41370
rect 44362 41318 44374 41370
rect 44436 41318 44438 41370
rect 44276 41316 44300 41318
rect 44356 41316 44380 41318
rect 44436 41316 44460 41318
rect 44220 41296 44516 41316
rect 44220 40284 44516 40304
rect 44276 40282 44300 40284
rect 44356 40282 44380 40284
rect 44436 40282 44460 40284
rect 44298 40230 44300 40282
rect 44362 40230 44374 40282
rect 44436 40230 44438 40282
rect 44276 40228 44300 40230
rect 44356 40228 44380 40230
rect 44436 40228 44460 40230
rect 44220 40208 44516 40228
rect 44560 39302 44588 41414
rect 43996 39296 44048 39302
rect 43996 39238 44048 39244
rect 44548 39296 44600 39302
rect 44548 39238 44600 39244
rect 43260 30252 43312 30258
rect 43260 30194 43312 30200
rect 44008 29850 44036 39238
rect 44220 39196 44516 39216
rect 44276 39194 44300 39196
rect 44356 39194 44380 39196
rect 44436 39194 44460 39196
rect 44298 39142 44300 39194
rect 44362 39142 44374 39194
rect 44436 39142 44438 39194
rect 44276 39140 44300 39142
rect 44356 39140 44380 39142
rect 44436 39140 44460 39142
rect 44220 39120 44516 39140
rect 44220 38108 44516 38128
rect 44276 38106 44300 38108
rect 44356 38106 44380 38108
rect 44436 38106 44460 38108
rect 44298 38054 44300 38106
rect 44362 38054 44374 38106
rect 44436 38054 44438 38106
rect 44276 38052 44300 38054
rect 44356 38052 44380 38054
rect 44436 38052 44460 38054
rect 44220 38032 44516 38052
rect 44220 37020 44516 37040
rect 44276 37018 44300 37020
rect 44356 37018 44380 37020
rect 44436 37018 44460 37020
rect 44298 36966 44300 37018
rect 44362 36966 44374 37018
rect 44436 36966 44438 37018
rect 44276 36964 44300 36966
rect 44356 36964 44380 36966
rect 44436 36964 44460 36966
rect 44220 36944 44516 36964
rect 44220 35932 44516 35952
rect 44276 35930 44300 35932
rect 44356 35930 44380 35932
rect 44436 35930 44460 35932
rect 44298 35878 44300 35930
rect 44362 35878 44374 35930
rect 44436 35878 44438 35930
rect 44276 35876 44300 35878
rect 44356 35876 44380 35878
rect 44436 35876 44460 35878
rect 44220 35856 44516 35876
rect 47676 35624 47728 35630
rect 47676 35566 47728 35572
rect 44220 34844 44516 34864
rect 44276 34842 44300 34844
rect 44356 34842 44380 34844
rect 44436 34842 44460 34844
rect 44298 34790 44300 34842
rect 44362 34790 44374 34842
rect 44436 34790 44438 34842
rect 44276 34788 44300 34790
rect 44356 34788 44380 34790
rect 44436 34788 44460 34790
rect 44220 34768 44516 34788
rect 44220 33756 44516 33776
rect 44276 33754 44300 33756
rect 44356 33754 44380 33756
rect 44436 33754 44460 33756
rect 44298 33702 44300 33754
rect 44362 33702 44374 33754
rect 44436 33702 44438 33754
rect 44276 33700 44300 33702
rect 44356 33700 44380 33702
rect 44436 33700 44460 33702
rect 44220 33680 44516 33700
rect 47032 33312 47084 33318
rect 47032 33254 47084 33260
rect 47044 32910 47072 33254
rect 47032 32904 47084 32910
rect 47032 32846 47084 32852
rect 46756 32768 46808 32774
rect 46756 32710 46808 32716
rect 44220 32668 44516 32688
rect 44276 32666 44300 32668
rect 44356 32666 44380 32668
rect 44436 32666 44460 32668
rect 44298 32614 44300 32666
rect 44362 32614 44374 32666
rect 44436 32614 44438 32666
rect 44276 32612 44300 32614
rect 44356 32612 44380 32614
rect 44436 32612 44460 32614
rect 44220 32592 44516 32612
rect 45560 32564 45612 32570
rect 45560 32506 45612 32512
rect 44220 31580 44516 31600
rect 44276 31578 44300 31580
rect 44356 31578 44380 31580
rect 44436 31578 44460 31580
rect 44298 31526 44300 31578
rect 44362 31526 44374 31578
rect 44436 31526 44438 31578
rect 44276 31524 44300 31526
rect 44356 31524 44380 31526
rect 44436 31524 44460 31526
rect 44220 31504 44516 31524
rect 44220 30492 44516 30512
rect 44276 30490 44300 30492
rect 44356 30490 44380 30492
rect 44436 30490 44460 30492
rect 44298 30438 44300 30490
rect 44362 30438 44374 30490
rect 44436 30438 44438 30490
rect 44276 30436 44300 30438
rect 44356 30436 44380 30438
rect 44436 30436 44460 30438
rect 44220 30416 44516 30436
rect 44088 30320 44140 30326
rect 44088 30262 44140 30268
rect 43996 29844 44048 29850
rect 43996 29786 44048 29792
rect 44008 29238 44036 29786
rect 44100 29306 44128 30262
rect 45008 30184 45060 30190
rect 45008 30126 45060 30132
rect 45020 29646 45048 30126
rect 45008 29640 45060 29646
rect 45008 29582 45060 29588
rect 45192 29572 45244 29578
rect 45192 29514 45244 29520
rect 44548 29504 44600 29510
rect 44548 29446 44600 29452
rect 44220 29404 44516 29424
rect 44276 29402 44300 29404
rect 44356 29402 44380 29404
rect 44436 29402 44460 29404
rect 44298 29350 44300 29402
rect 44362 29350 44374 29402
rect 44436 29350 44438 29402
rect 44276 29348 44300 29350
rect 44356 29348 44380 29350
rect 44436 29348 44460 29350
rect 44220 29328 44516 29348
rect 44088 29300 44140 29306
rect 44088 29242 44140 29248
rect 43996 29232 44048 29238
rect 43996 29174 44048 29180
rect 43444 28144 43496 28150
rect 43444 28086 43496 28092
rect 43352 16040 43404 16046
rect 43352 15982 43404 15988
rect 43364 15706 43392 15982
rect 43352 15700 43404 15706
rect 43352 15642 43404 15648
rect 43260 7472 43312 7478
rect 43260 7414 43312 7420
rect 42524 3732 42576 3738
rect 42524 3674 42576 3680
rect 42800 3732 42852 3738
rect 42800 3674 42852 3680
rect 42536 3602 42564 3674
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 42340 3596 42392 3602
rect 42340 3538 42392 3544
rect 42524 3596 42576 3602
rect 42524 3538 42576 3544
rect 41248 3194 41276 3538
rect 42432 3460 42484 3466
rect 42432 3402 42484 3408
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 42444 3126 42472 3402
rect 42432 3120 42484 3126
rect 42432 3062 42484 3068
rect 39028 3052 39080 3058
rect 39028 2994 39080 3000
rect 43272 2990 43300 7414
rect 43364 3738 43392 15642
rect 43456 11898 43484 28086
rect 43536 23860 43588 23866
rect 43536 23802 43588 23808
rect 43444 11892 43496 11898
rect 43444 11834 43496 11840
rect 43548 4146 43576 23802
rect 44008 16046 44036 29174
rect 44100 29170 44128 29242
rect 44088 29164 44140 29170
rect 44088 29106 44140 29112
rect 44560 29102 44588 29446
rect 45204 29102 45232 29514
rect 44180 29096 44232 29102
rect 44180 29038 44232 29044
rect 44548 29096 44600 29102
rect 44548 29038 44600 29044
rect 45192 29096 45244 29102
rect 45192 29038 45244 29044
rect 44192 28762 44220 29038
rect 44180 28756 44232 28762
rect 44180 28698 44232 28704
rect 44220 28316 44516 28336
rect 44276 28314 44300 28316
rect 44356 28314 44380 28316
rect 44436 28314 44460 28316
rect 44298 28262 44300 28314
rect 44362 28262 44374 28314
rect 44436 28262 44438 28314
rect 44276 28260 44300 28262
rect 44356 28260 44380 28262
rect 44436 28260 44460 28262
rect 44220 28240 44516 28260
rect 44220 27228 44516 27248
rect 44276 27226 44300 27228
rect 44356 27226 44380 27228
rect 44436 27226 44460 27228
rect 44298 27174 44300 27226
rect 44362 27174 44374 27226
rect 44436 27174 44438 27226
rect 44276 27172 44300 27174
rect 44356 27172 44380 27174
rect 44436 27172 44460 27174
rect 44220 27152 44516 27172
rect 44220 26140 44516 26160
rect 44276 26138 44300 26140
rect 44356 26138 44380 26140
rect 44436 26138 44460 26140
rect 44298 26086 44300 26138
rect 44362 26086 44374 26138
rect 44436 26086 44438 26138
rect 44276 26084 44300 26086
rect 44356 26084 44380 26086
rect 44436 26084 44460 26086
rect 44220 26064 44516 26084
rect 45192 25356 45244 25362
rect 45192 25298 45244 25304
rect 45204 25158 45232 25298
rect 45192 25152 45244 25158
rect 45192 25094 45244 25100
rect 44220 25052 44516 25072
rect 44276 25050 44300 25052
rect 44356 25050 44380 25052
rect 44436 25050 44460 25052
rect 44298 24998 44300 25050
rect 44362 24998 44374 25050
rect 44436 24998 44438 25050
rect 44276 24996 44300 24998
rect 44356 24996 44380 24998
rect 44436 24996 44460 24998
rect 44220 24976 44516 24996
rect 44220 23964 44516 23984
rect 44276 23962 44300 23964
rect 44356 23962 44380 23964
rect 44436 23962 44460 23964
rect 44298 23910 44300 23962
rect 44362 23910 44374 23962
rect 44436 23910 44438 23962
rect 44276 23908 44300 23910
rect 44356 23908 44380 23910
rect 44436 23908 44460 23910
rect 44220 23888 44516 23908
rect 44220 22876 44516 22896
rect 44276 22874 44300 22876
rect 44356 22874 44380 22876
rect 44436 22874 44460 22876
rect 44298 22822 44300 22874
rect 44362 22822 44374 22874
rect 44436 22822 44438 22874
rect 44276 22820 44300 22822
rect 44356 22820 44380 22822
rect 44436 22820 44460 22822
rect 44220 22800 44516 22820
rect 44220 21788 44516 21808
rect 44276 21786 44300 21788
rect 44356 21786 44380 21788
rect 44436 21786 44460 21788
rect 44298 21734 44300 21786
rect 44362 21734 44374 21786
rect 44436 21734 44438 21786
rect 44276 21732 44300 21734
rect 44356 21732 44380 21734
rect 44436 21732 44460 21734
rect 44220 21712 44516 21732
rect 44220 20700 44516 20720
rect 44276 20698 44300 20700
rect 44356 20698 44380 20700
rect 44436 20698 44460 20700
rect 44298 20646 44300 20698
rect 44362 20646 44374 20698
rect 44436 20646 44438 20698
rect 44276 20644 44300 20646
rect 44356 20644 44380 20646
rect 44436 20644 44460 20646
rect 44220 20624 44516 20644
rect 44548 20256 44600 20262
rect 44548 20198 44600 20204
rect 44220 19612 44516 19632
rect 44276 19610 44300 19612
rect 44356 19610 44380 19612
rect 44436 19610 44460 19612
rect 44298 19558 44300 19610
rect 44362 19558 44374 19610
rect 44436 19558 44438 19610
rect 44276 19556 44300 19558
rect 44356 19556 44380 19558
rect 44436 19556 44460 19558
rect 44220 19536 44516 19556
rect 44220 18524 44516 18544
rect 44276 18522 44300 18524
rect 44356 18522 44380 18524
rect 44436 18522 44460 18524
rect 44298 18470 44300 18522
rect 44362 18470 44374 18522
rect 44436 18470 44438 18522
rect 44276 18468 44300 18470
rect 44356 18468 44380 18470
rect 44436 18468 44460 18470
rect 44220 18448 44516 18468
rect 44220 17436 44516 17456
rect 44276 17434 44300 17436
rect 44356 17434 44380 17436
rect 44436 17434 44460 17436
rect 44298 17382 44300 17434
rect 44362 17382 44374 17434
rect 44436 17382 44438 17434
rect 44276 17380 44300 17382
rect 44356 17380 44380 17382
rect 44436 17380 44460 17382
rect 44220 17360 44516 17380
rect 44220 16348 44516 16368
rect 44276 16346 44300 16348
rect 44356 16346 44380 16348
rect 44436 16346 44460 16348
rect 44298 16294 44300 16346
rect 44362 16294 44374 16346
rect 44436 16294 44438 16346
rect 44276 16292 44300 16294
rect 44356 16292 44380 16294
rect 44436 16292 44460 16294
rect 44220 16272 44516 16292
rect 43996 16040 44048 16046
rect 43996 15982 44048 15988
rect 44220 15260 44516 15280
rect 44276 15258 44300 15260
rect 44356 15258 44380 15260
rect 44436 15258 44460 15260
rect 44298 15206 44300 15258
rect 44362 15206 44374 15258
rect 44436 15206 44438 15258
rect 44276 15204 44300 15206
rect 44356 15204 44380 15206
rect 44436 15204 44460 15206
rect 44220 15184 44516 15204
rect 44220 14172 44516 14192
rect 44276 14170 44300 14172
rect 44356 14170 44380 14172
rect 44436 14170 44460 14172
rect 44298 14118 44300 14170
rect 44362 14118 44374 14170
rect 44436 14118 44438 14170
rect 44276 14116 44300 14118
rect 44356 14116 44380 14118
rect 44436 14116 44460 14118
rect 44220 14096 44516 14116
rect 44220 13084 44516 13104
rect 44276 13082 44300 13084
rect 44356 13082 44380 13084
rect 44436 13082 44460 13084
rect 44298 13030 44300 13082
rect 44362 13030 44374 13082
rect 44436 13030 44438 13082
rect 44276 13028 44300 13030
rect 44356 13028 44380 13030
rect 44436 13028 44460 13030
rect 44220 13008 44516 13028
rect 44220 11996 44516 12016
rect 44276 11994 44300 11996
rect 44356 11994 44380 11996
rect 44436 11994 44460 11996
rect 44298 11942 44300 11994
rect 44362 11942 44374 11994
rect 44436 11942 44438 11994
rect 44276 11940 44300 11942
rect 44356 11940 44380 11942
rect 44436 11940 44460 11942
rect 44220 11920 44516 11940
rect 43720 11688 43772 11694
rect 43720 11630 43772 11636
rect 43732 11354 43760 11630
rect 43720 11348 43772 11354
rect 43720 11290 43772 11296
rect 44220 10908 44516 10928
rect 44276 10906 44300 10908
rect 44356 10906 44380 10908
rect 44436 10906 44460 10908
rect 44298 10854 44300 10906
rect 44362 10854 44374 10906
rect 44436 10854 44438 10906
rect 44276 10852 44300 10854
rect 44356 10852 44380 10854
rect 44436 10852 44460 10854
rect 44220 10832 44516 10852
rect 44220 9820 44516 9840
rect 44276 9818 44300 9820
rect 44356 9818 44380 9820
rect 44436 9818 44460 9820
rect 44298 9766 44300 9818
rect 44362 9766 44374 9818
rect 44436 9766 44438 9818
rect 44276 9764 44300 9766
rect 44356 9764 44380 9766
rect 44436 9764 44460 9766
rect 44220 9744 44516 9764
rect 44220 8732 44516 8752
rect 44276 8730 44300 8732
rect 44356 8730 44380 8732
rect 44436 8730 44460 8732
rect 44298 8678 44300 8730
rect 44362 8678 44374 8730
rect 44436 8678 44438 8730
rect 44276 8676 44300 8678
rect 44356 8676 44380 8678
rect 44436 8676 44460 8678
rect 44220 8656 44516 8676
rect 44220 7644 44516 7664
rect 44276 7642 44300 7644
rect 44356 7642 44380 7644
rect 44436 7642 44460 7644
rect 44298 7590 44300 7642
rect 44362 7590 44374 7642
rect 44436 7590 44438 7642
rect 44276 7588 44300 7590
rect 44356 7588 44380 7590
rect 44436 7588 44460 7590
rect 44220 7568 44516 7588
rect 44220 6556 44516 6576
rect 44276 6554 44300 6556
rect 44356 6554 44380 6556
rect 44436 6554 44460 6556
rect 44298 6502 44300 6554
rect 44362 6502 44374 6554
rect 44436 6502 44438 6554
rect 44276 6500 44300 6502
rect 44356 6500 44380 6502
rect 44436 6500 44460 6502
rect 44220 6480 44516 6500
rect 44220 5468 44516 5488
rect 44276 5466 44300 5468
rect 44356 5466 44380 5468
rect 44436 5466 44460 5468
rect 44298 5414 44300 5466
rect 44362 5414 44374 5466
rect 44436 5414 44438 5466
rect 44276 5412 44300 5414
rect 44356 5412 44380 5414
rect 44436 5412 44460 5414
rect 44220 5392 44516 5412
rect 44220 4380 44516 4400
rect 44276 4378 44300 4380
rect 44356 4378 44380 4380
rect 44436 4378 44460 4380
rect 44298 4326 44300 4378
rect 44362 4326 44374 4378
rect 44436 4326 44438 4378
rect 44276 4324 44300 4326
rect 44356 4324 44380 4326
rect 44436 4324 44460 4326
rect 44220 4304 44516 4324
rect 43536 4140 43588 4146
rect 43536 4082 43588 4088
rect 43352 3732 43404 3738
rect 43352 3674 43404 3680
rect 43364 3466 43392 3674
rect 43548 3670 43576 4082
rect 44560 3738 44588 20198
rect 44640 14612 44692 14618
rect 44640 14554 44692 14560
rect 44652 4146 44680 14554
rect 45204 9110 45232 25094
rect 45572 11898 45600 32506
rect 45928 25696 45980 25702
rect 45928 25638 45980 25644
rect 45652 25492 45704 25498
rect 45652 25434 45704 25440
rect 45664 24750 45692 25434
rect 45940 25430 45968 25638
rect 46768 25498 46796 32710
rect 47044 28626 47072 32846
rect 47584 32768 47636 32774
rect 47584 32710 47636 32716
rect 47596 30802 47624 32710
rect 47584 30796 47636 30802
rect 47584 30738 47636 30744
rect 47032 28620 47084 28626
rect 47032 28562 47084 28568
rect 46756 25492 46808 25498
rect 46756 25434 46808 25440
rect 45928 25424 45980 25430
rect 45928 25366 45980 25372
rect 46768 25362 46796 25434
rect 46572 25356 46624 25362
rect 46572 25298 46624 25304
rect 46756 25356 46808 25362
rect 46756 25298 46808 25304
rect 46204 25152 46256 25158
rect 46204 25094 46256 25100
rect 45652 24744 45704 24750
rect 45652 24686 45704 24692
rect 45560 11892 45612 11898
rect 45560 11834 45612 11840
rect 45192 9104 45244 9110
rect 45192 9046 45244 9052
rect 44640 4140 44692 4146
rect 44640 4082 44692 4088
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 43536 3664 43588 3670
rect 43536 3606 43588 3612
rect 44652 3602 44680 4082
rect 44640 3596 44692 3602
rect 44640 3538 44692 3544
rect 43352 3460 43404 3466
rect 43352 3402 43404 3408
rect 44220 3292 44516 3312
rect 44276 3290 44300 3292
rect 44356 3290 44380 3292
rect 44436 3290 44460 3292
rect 44298 3238 44300 3290
rect 44362 3238 44374 3290
rect 44436 3238 44438 3290
rect 44276 3236 44300 3238
rect 44356 3236 44380 3238
rect 44436 3236 44460 3238
rect 44220 3216 44516 3236
rect 46216 3058 46244 25094
rect 46584 24954 46612 25298
rect 46572 24948 46624 24954
rect 46572 24890 46624 24896
rect 47688 15570 47716 35566
rect 47860 32972 47912 32978
rect 47860 32914 47912 32920
rect 47872 32570 47900 32914
rect 47860 32564 47912 32570
rect 47860 32506 47912 32512
rect 48136 25356 48188 25362
rect 48136 25298 48188 25304
rect 47952 25152 48004 25158
rect 47952 25094 48004 25100
rect 47676 15564 47728 15570
rect 47676 15506 47728 15512
rect 47964 9382 47992 25094
rect 48148 24993 48176 25298
rect 48134 24984 48190 24993
rect 48134 24919 48190 24928
rect 47952 9376 48004 9382
rect 47952 9318 48004 9324
rect 48136 9036 48188 9042
rect 48136 8978 48188 8984
rect 47952 8832 48004 8838
rect 47952 8774 48004 8780
rect 47964 8634 47992 8774
rect 47952 8628 48004 8634
rect 47952 8570 48004 8576
rect 48148 8401 48176 8978
rect 48134 8392 48190 8401
rect 48134 8327 48190 8336
rect 46204 3052 46256 3058
rect 46204 2994 46256 3000
rect 43260 2984 43312 2990
rect 43260 2926 43312 2932
rect 37924 2848 37976 2854
rect 37924 2790 37976 2796
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 37936 2514 37964 2790
rect 39220 2748 39516 2768
rect 39276 2746 39300 2748
rect 39356 2746 39380 2748
rect 39436 2746 39460 2748
rect 39298 2694 39300 2746
rect 39362 2694 39374 2746
rect 39436 2694 39438 2746
rect 39276 2692 39300 2694
rect 39356 2692 39380 2694
rect 39436 2692 39460 2694
rect 39220 2672 39516 2692
rect 43272 2650 43300 2926
rect 43260 2644 43312 2650
rect 43260 2586 43312 2592
rect 37372 2508 37424 2514
rect 37372 2450 37424 2456
rect 37924 2508 37976 2514
rect 37924 2450 37976 2456
rect 14220 2204 14516 2224
rect 14276 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14298 2150 14300 2202
rect 14362 2150 14374 2202
rect 14436 2150 14438 2202
rect 14276 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14220 2128 14516 2148
rect 37384 800 37412 2450
rect 44220 2204 44516 2224
rect 44276 2202 44300 2204
rect 44356 2202 44380 2204
rect 44436 2202 44460 2204
rect 44298 2150 44300 2202
rect 44362 2150 44374 2202
rect 44436 2150 44438 2202
rect 44276 2148 44300 2150
rect 44356 2148 44380 2150
rect 44436 2148 44460 2150
rect 44220 2128 44516 2148
rect 12438 0 12494 800
rect 37370 0 37426 800
<< via2 >>
rect 1858 47504 1914 47560
rect 9220 47354 9276 47356
rect 9300 47354 9356 47356
rect 9380 47354 9436 47356
rect 9460 47354 9516 47356
rect 9220 47302 9246 47354
rect 9246 47302 9276 47354
rect 9300 47302 9310 47354
rect 9310 47302 9356 47354
rect 9380 47302 9426 47354
rect 9426 47302 9436 47354
rect 9460 47302 9490 47354
rect 9490 47302 9516 47354
rect 9220 47300 9276 47302
rect 9300 47300 9356 47302
rect 9380 47300 9436 47302
rect 9460 47300 9516 47302
rect 19220 47354 19276 47356
rect 19300 47354 19356 47356
rect 19380 47354 19436 47356
rect 19460 47354 19516 47356
rect 19220 47302 19246 47354
rect 19246 47302 19276 47354
rect 19300 47302 19310 47354
rect 19310 47302 19356 47354
rect 19380 47302 19426 47354
rect 19426 47302 19436 47354
rect 19460 47302 19490 47354
rect 19490 47302 19516 47354
rect 19220 47300 19276 47302
rect 19300 47300 19356 47302
rect 19380 47300 19436 47302
rect 19460 47300 19516 47302
rect 29220 47354 29276 47356
rect 29300 47354 29356 47356
rect 29380 47354 29436 47356
rect 29460 47354 29516 47356
rect 29220 47302 29246 47354
rect 29246 47302 29276 47354
rect 29300 47302 29310 47354
rect 29310 47302 29356 47354
rect 29380 47302 29426 47354
rect 29426 47302 29436 47354
rect 29460 47302 29490 47354
rect 29490 47302 29516 47354
rect 29220 47300 29276 47302
rect 29300 47300 29356 47302
rect 29380 47300 29436 47302
rect 29460 47300 29516 47302
rect 39220 47354 39276 47356
rect 39300 47354 39356 47356
rect 39380 47354 39436 47356
rect 39460 47354 39516 47356
rect 39220 47302 39246 47354
rect 39246 47302 39276 47354
rect 39300 47302 39310 47354
rect 39310 47302 39356 47354
rect 39380 47302 39426 47354
rect 39426 47302 39436 47354
rect 39460 47302 39490 47354
rect 39490 47302 39516 47354
rect 39220 47300 39276 47302
rect 39300 47300 39356 47302
rect 39380 47300 39436 47302
rect 39460 47300 39516 47302
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 14220 46810 14276 46812
rect 14300 46810 14356 46812
rect 14380 46810 14436 46812
rect 14460 46810 14516 46812
rect 14220 46758 14246 46810
rect 14246 46758 14276 46810
rect 14300 46758 14310 46810
rect 14310 46758 14356 46810
rect 14380 46758 14426 46810
rect 14426 46758 14436 46810
rect 14460 46758 14490 46810
rect 14490 46758 14516 46810
rect 14220 46756 14276 46758
rect 14300 46756 14356 46758
rect 14380 46756 14436 46758
rect 14460 46756 14516 46758
rect 9220 46266 9276 46268
rect 9300 46266 9356 46268
rect 9380 46266 9436 46268
rect 9460 46266 9516 46268
rect 9220 46214 9246 46266
rect 9246 46214 9276 46266
rect 9300 46214 9310 46266
rect 9310 46214 9356 46266
rect 9380 46214 9426 46266
rect 9426 46214 9436 46266
rect 9460 46214 9490 46266
rect 9490 46214 9516 46266
rect 9220 46212 9276 46214
rect 9300 46212 9356 46214
rect 9380 46212 9436 46214
rect 9460 46212 9516 46214
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 14220 45722 14276 45724
rect 14300 45722 14356 45724
rect 14380 45722 14436 45724
rect 14460 45722 14516 45724
rect 14220 45670 14246 45722
rect 14246 45670 14276 45722
rect 14300 45670 14310 45722
rect 14310 45670 14356 45722
rect 14380 45670 14426 45722
rect 14426 45670 14436 45722
rect 14460 45670 14490 45722
rect 14490 45670 14516 45722
rect 14220 45668 14276 45670
rect 14300 45668 14356 45670
rect 14380 45668 14436 45670
rect 14460 45668 14516 45670
rect 1858 42508 1860 42528
rect 1860 42508 1912 42528
rect 1912 42508 1914 42528
rect 1858 42472 1914 42508
rect 1858 37460 1914 37496
rect 1858 37440 1860 37460
rect 1860 37440 1912 37460
rect 1912 37440 1914 37460
rect 1766 32428 1822 32464
rect 1766 32408 1768 32428
rect 1768 32408 1820 32428
rect 1820 32408 1822 32428
rect 1766 27548 1768 27568
rect 1768 27548 1820 27568
rect 1820 27548 1822 27568
rect 1766 27512 1822 27548
rect 9220 45178 9276 45180
rect 9300 45178 9356 45180
rect 9380 45178 9436 45180
rect 9460 45178 9516 45180
rect 9220 45126 9246 45178
rect 9246 45126 9276 45178
rect 9300 45126 9310 45178
rect 9310 45126 9356 45178
rect 9380 45126 9426 45178
rect 9426 45126 9436 45178
rect 9460 45126 9490 45178
rect 9490 45126 9516 45178
rect 9220 45124 9276 45126
rect 9300 45124 9356 45126
rect 9380 45124 9436 45126
rect 9460 45124 9516 45126
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 14220 44634 14276 44636
rect 14300 44634 14356 44636
rect 14380 44634 14436 44636
rect 14460 44634 14516 44636
rect 14220 44582 14246 44634
rect 14246 44582 14276 44634
rect 14300 44582 14310 44634
rect 14310 44582 14356 44634
rect 14380 44582 14426 44634
rect 14426 44582 14436 44634
rect 14460 44582 14490 44634
rect 14490 44582 14516 44634
rect 14220 44580 14276 44582
rect 14300 44580 14356 44582
rect 14380 44580 14436 44582
rect 14460 44580 14516 44582
rect 9220 44090 9276 44092
rect 9300 44090 9356 44092
rect 9380 44090 9436 44092
rect 9460 44090 9516 44092
rect 9220 44038 9246 44090
rect 9246 44038 9276 44090
rect 9300 44038 9310 44090
rect 9310 44038 9356 44090
rect 9380 44038 9426 44090
rect 9426 44038 9436 44090
rect 9460 44038 9490 44090
rect 9490 44038 9516 44090
rect 9220 44036 9276 44038
rect 9300 44036 9356 44038
rect 9380 44036 9436 44038
rect 9460 44036 9516 44038
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 14220 43546 14276 43548
rect 14300 43546 14356 43548
rect 14380 43546 14436 43548
rect 14460 43546 14516 43548
rect 14220 43494 14246 43546
rect 14246 43494 14276 43546
rect 14300 43494 14310 43546
rect 14310 43494 14356 43546
rect 14380 43494 14426 43546
rect 14426 43494 14436 43546
rect 14460 43494 14490 43546
rect 14490 43494 14516 43546
rect 14220 43492 14276 43494
rect 14300 43492 14356 43494
rect 14380 43492 14436 43494
rect 14460 43492 14516 43494
rect 9220 43002 9276 43004
rect 9300 43002 9356 43004
rect 9380 43002 9436 43004
rect 9460 43002 9516 43004
rect 9220 42950 9246 43002
rect 9246 42950 9276 43002
rect 9300 42950 9310 43002
rect 9310 42950 9356 43002
rect 9380 42950 9426 43002
rect 9426 42950 9436 43002
rect 9460 42950 9490 43002
rect 9490 42950 9516 43002
rect 9220 42948 9276 42950
rect 9300 42948 9356 42950
rect 9380 42948 9436 42950
rect 9460 42948 9516 42950
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 9220 41914 9276 41916
rect 9300 41914 9356 41916
rect 9380 41914 9436 41916
rect 9460 41914 9516 41916
rect 9220 41862 9246 41914
rect 9246 41862 9276 41914
rect 9300 41862 9310 41914
rect 9310 41862 9356 41914
rect 9380 41862 9426 41914
rect 9426 41862 9436 41914
rect 9460 41862 9490 41914
rect 9490 41862 9516 41914
rect 9220 41860 9276 41862
rect 9300 41860 9356 41862
rect 9380 41860 9436 41862
rect 9460 41860 9516 41862
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 9220 40826 9276 40828
rect 9300 40826 9356 40828
rect 9380 40826 9436 40828
rect 9460 40826 9516 40828
rect 9220 40774 9246 40826
rect 9246 40774 9276 40826
rect 9300 40774 9310 40826
rect 9310 40774 9356 40826
rect 9380 40774 9426 40826
rect 9426 40774 9436 40826
rect 9460 40774 9490 40826
rect 9490 40774 9516 40826
rect 9220 40772 9276 40774
rect 9300 40772 9356 40774
rect 9380 40772 9436 40774
rect 9460 40772 9516 40774
rect 9220 39738 9276 39740
rect 9300 39738 9356 39740
rect 9380 39738 9436 39740
rect 9460 39738 9516 39740
rect 9220 39686 9246 39738
rect 9246 39686 9276 39738
rect 9300 39686 9310 39738
rect 9310 39686 9356 39738
rect 9380 39686 9426 39738
rect 9426 39686 9436 39738
rect 9460 39686 9490 39738
rect 9490 39686 9516 39738
rect 9220 39684 9276 39686
rect 9300 39684 9356 39686
rect 9380 39684 9436 39686
rect 9460 39684 9516 39686
rect 9220 38650 9276 38652
rect 9300 38650 9356 38652
rect 9380 38650 9436 38652
rect 9460 38650 9516 38652
rect 9220 38598 9246 38650
rect 9246 38598 9276 38650
rect 9300 38598 9310 38650
rect 9310 38598 9356 38650
rect 9380 38598 9426 38650
rect 9426 38598 9436 38650
rect 9460 38598 9490 38650
rect 9490 38598 9516 38650
rect 9220 38596 9276 38598
rect 9300 38596 9356 38598
rect 9380 38596 9436 38598
rect 9460 38596 9516 38598
rect 9220 37562 9276 37564
rect 9300 37562 9356 37564
rect 9380 37562 9436 37564
rect 9460 37562 9516 37564
rect 9220 37510 9246 37562
rect 9246 37510 9276 37562
rect 9300 37510 9310 37562
rect 9310 37510 9356 37562
rect 9380 37510 9426 37562
rect 9426 37510 9436 37562
rect 9460 37510 9490 37562
rect 9490 37510 9516 37562
rect 9220 37508 9276 37510
rect 9300 37508 9356 37510
rect 9380 37508 9436 37510
rect 9460 37508 9516 37510
rect 9220 36474 9276 36476
rect 9300 36474 9356 36476
rect 9380 36474 9436 36476
rect 9460 36474 9516 36476
rect 9220 36422 9246 36474
rect 9246 36422 9276 36474
rect 9300 36422 9310 36474
rect 9310 36422 9356 36474
rect 9380 36422 9426 36474
rect 9426 36422 9436 36474
rect 9460 36422 9490 36474
rect 9490 36422 9516 36474
rect 9220 36420 9276 36422
rect 9300 36420 9356 36422
rect 9380 36420 9436 36422
rect 9460 36420 9516 36422
rect 9220 35386 9276 35388
rect 9300 35386 9356 35388
rect 9380 35386 9436 35388
rect 9460 35386 9516 35388
rect 9220 35334 9246 35386
rect 9246 35334 9276 35386
rect 9300 35334 9310 35386
rect 9310 35334 9356 35386
rect 9380 35334 9426 35386
rect 9426 35334 9436 35386
rect 9460 35334 9490 35386
rect 9490 35334 9516 35386
rect 9220 35332 9276 35334
rect 9300 35332 9356 35334
rect 9380 35332 9436 35334
rect 9460 35332 9516 35334
rect 9220 34298 9276 34300
rect 9300 34298 9356 34300
rect 9380 34298 9436 34300
rect 9460 34298 9516 34300
rect 9220 34246 9246 34298
rect 9246 34246 9276 34298
rect 9300 34246 9310 34298
rect 9310 34246 9356 34298
rect 9380 34246 9426 34298
rect 9426 34246 9436 34298
rect 9460 34246 9490 34298
rect 9490 34246 9516 34298
rect 9220 34244 9276 34246
rect 9300 34244 9356 34246
rect 9380 34244 9436 34246
rect 9460 34244 9516 34246
rect 9220 33210 9276 33212
rect 9300 33210 9356 33212
rect 9380 33210 9436 33212
rect 9460 33210 9516 33212
rect 9220 33158 9246 33210
rect 9246 33158 9276 33210
rect 9300 33158 9310 33210
rect 9310 33158 9356 33210
rect 9380 33158 9426 33210
rect 9426 33158 9436 33210
rect 9460 33158 9490 33210
rect 9490 33158 9516 33210
rect 9220 33156 9276 33158
rect 9300 33156 9356 33158
rect 9380 33156 9436 33158
rect 9460 33156 9516 33158
rect 9220 32122 9276 32124
rect 9300 32122 9356 32124
rect 9380 32122 9436 32124
rect 9460 32122 9516 32124
rect 9220 32070 9246 32122
rect 9246 32070 9276 32122
rect 9300 32070 9310 32122
rect 9310 32070 9356 32122
rect 9380 32070 9426 32122
rect 9426 32070 9436 32122
rect 9460 32070 9490 32122
rect 9490 32070 9516 32122
rect 9220 32068 9276 32070
rect 9300 32068 9356 32070
rect 9380 32068 9436 32070
rect 9460 32068 9516 32070
rect 9220 31034 9276 31036
rect 9300 31034 9356 31036
rect 9380 31034 9436 31036
rect 9460 31034 9516 31036
rect 9220 30982 9246 31034
rect 9246 30982 9276 31034
rect 9300 30982 9310 31034
rect 9310 30982 9356 31034
rect 9380 30982 9426 31034
rect 9426 30982 9436 31034
rect 9460 30982 9490 31034
rect 9490 30982 9516 31034
rect 9220 30980 9276 30982
rect 9300 30980 9356 30982
rect 9380 30980 9436 30982
rect 9460 30980 9516 30982
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 1766 22500 1822 22536
rect 1766 22480 1768 22500
rect 1768 22480 1820 22500
rect 1820 22480 1822 22500
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 1858 17484 1860 17504
rect 1860 17484 1912 17504
rect 1912 17484 1914 17504
rect 1858 17448 1914 17484
rect 1858 12436 1914 12472
rect 1858 12416 1860 12436
rect 1860 12416 1912 12436
rect 1912 12416 1914 12436
rect 1766 7420 1768 7440
rect 1768 7420 1820 7440
rect 1820 7420 1822 7440
rect 1766 7384 1822 7420
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 9220 29946 9276 29948
rect 9300 29946 9356 29948
rect 9380 29946 9436 29948
rect 9460 29946 9516 29948
rect 9220 29894 9246 29946
rect 9246 29894 9276 29946
rect 9300 29894 9310 29946
rect 9310 29894 9356 29946
rect 9380 29894 9426 29946
rect 9426 29894 9436 29946
rect 9460 29894 9490 29946
rect 9490 29894 9516 29946
rect 9220 29892 9276 29894
rect 9300 29892 9356 29894
rect 9380 29892 9436 29894
rect 9460 29892 9516 29894
rect 9220 28858 9276 28860
rect 9300 28858 9356 28860
rect 9380 28858 9436 28860
rect 9460 28858 9516 28860
rect 9220 28806 9246 28858
rect 9246 28806 9276 28858
rect 9300 28806 9310 28858
rect 9310 28806 9356 28858
rect 9380 28806 9426 28858
rect 9426 28806 9436 28858
rect 9460 28806 9490 28858
rect 9490 28806 9516 28858
rect 9220 28804 9276 28806
rect 9300 28804 9356 28806
rect 9380 28804 9436 28806
rect 9460 28804 9516 28806
rect 9220 27770 9276 27772
rect 9300 27770 9356 27772
rect 9380 27770 9436 27772
rect 9460 27770 9516 27772
rect 9220 27718 9246 27770
rect 9246 27718 9276 27770
rect 9300 27718 9310 27770
rect 9310 27718 9356 27770
rect 9380 27718 9426 27770
rect 9426 27718 9436 27770
rect 9460 27718 9490 27770
rect 9490 27718 9516 27770
rect 9220 27716 9276 27718
rect 9300 27716 9356 27718
rect 9380 27716 9436 27718
rect 9460 27716 9516 27718
rect 9220 26682 9276 26684
rect 9300 26682 9356 26684
rect 9380 26682 9436 26684
rect 9460 26682 9516 26684
rect 9220 26630 9246 26682
rect 9246 26630 9276 26682
rect 9300 26630 9310 26682
rect 9310 26630 9356 26682
rect 9380 26630 9426 26682
rect 9426 26630 9436 26682
rect 9460 26630 9490 26682
rect 9490 26630 9516 26682
rect 9220 26628 9276 26630
rect 9300 26628 9356 26630
rect 9380 26628 9436 26630
rect 9460 26628 9516 26630
rect 9220 25594 9276 25596
rect 9300 25594 9356 25596
rect 9380 25594 9436 25596
rect 9460 25594 9516 25596
rect 9220 25542 9246 25594
rect 9246 25542 9276 25594
rect 9300 25542 9310 25594
rect 9310 25542 9356 25594
rect 9380 25542 9426 25594
rect 9426 25542 9436 25594
rect 9460 25542 9490 25594
rect 9490 25542 9516 25594
rect 9220 25540 9276 25542
rect 9300 25540 9356 25542
rect 9380 25540 9436 25542
rect 9460 25540 9516 25542
rect 9220 24506 9276 24508
rect 9300 24506 9356 24508
rect 9380 24506 9436 24508
rect 9460 24506 9516 24508
rect 9220 24454 9246 24506
rect 9246 24454 9276 24506
rect 9300 24454 9310 24506
rect 9310 24454 9356 24506
rect 9380 24454 9426 24506
rect 9426 24454 9436 24506
rect 9460 24454 9490 24506
rect 9490 24454 9516 24506
rect 9220 24452 9276 24454
rect 9300 24452 9356 24454
rect 9380 24452 9436 24454
rect 9460 24452 9516 24454
rect 9220 23418 9276 23420
rect 9300 23418 9356 23420
rect 9380 23418 9436 23420
rect 9460 23418 9516 23420
rect 9220 23366 9246 23418
rect 9246 23366 9276 23418
rect 9300 23366 9310 23418
rect 9310 23366 9356 23418
rect 9380 23366 9426 23418
rect 9426 23366 9436 23418
rect 9460 23366 9490 23418
rect 9490 23366 9516 23418
rect 9220 23364 9276 23366
rect 9300 23364 9356 23366
rect 9380 23364 9436 23366
rect 9460 23364 9516 23366
rect 9220 22330 9276 22332
rect 9300 22330 9356 22332
rect 9380 22330 9436 22332
rect 9460 22330 9516 22332
rect 9220 22278 9246 22330
rect 9246 22278 9276 22330
rect 9300 22278 9310 22330
rect 9310 22278 9356 22330
rect 9380 22278 9426 22330
rect 9426 22278 9436 22330
rect 9460 22278 9490 22330
rect 9490 22278 9516 22330
rect 9220 22276 9276 22278
rect 9300 22276 9356 22278
rect 9380 22276 9436 22278
rect 9460 22276 9516 22278
rect 9220 21242 9276 21244
rect 9300 21242 9356 21244
rect 9380 21242 9436 21244
rect 9460 21242 9516 21244
rect 9220 21190 9246 21242
rect 9246 21190 9276 21242
rect 9300 21190 9310 21242
rect 9310 21190 9356 21242
rect 9380 21190 9426 21242
rect 9426 21190 9436 21242
rect 9460 21190 9490 21242
rect 9490 21190 9516 21242
rect 9220 21188 9276 21190
rect 9300 21188 9356 21190
rect 9380 21188 9436 21190
rect 9460 21188 9516 21190
rect 9220 20154 9276 20156
rect 9300 20154 9356 20156
rect 9380 20154 9436 20156
rect 9460 20154 9516 20156
rect 9220 20102 9246 20154
rect 9246 20102 9276 20154
rect 9300 20102 9310 20154
rect 9310 20102 9356 20154
rect 9380 20102 9426 20154
rect 9426 20102 9436 20154
rect 9460 20102 9490 20154
rect 9490 20102 9516 20154
rect 9220 20100 9276 20102
rect 9300 20100 9356 20102
rect 9380 20100 9436 20102
rect 9460 20100 9516 20102
rect 9220 19066 9276 19068
rect 9300 19066 9356 19068
rect 9380 19066 9436 19068
rect 9460 19066 9516 19068
rect 9220 19014 9246 19066
rect 9246 19014 9276 19066
rect 9300 19014 9310 19066
rect 9310 19014 9356 19066
rect 9380 19014 9426 19066
rect 9426 19014 9436 19066
rect 9460 19014 9490 19066
rect 9490 19014 9516 19066
rect 9220 19012 9276 19014
rect 9300 19012 9356 19014
rect 9380 19012 9436 19014
rect 9460 19012 9516 19014
rect 9220 17978 9276 17980
rect 9300 17978 9356 17980
rect 9380 17978 9436 17980
rect 9460 17978 9516 17980
rect 9220 17926 9246 17978
rect 9246 17926 9276 17978
rect 9300 17926 9310 17978
rect 9310 17926 9356 17978
rect 9380 17926 9426 17978
rect 9426 17926 9436 17978
rect 9460 17926 9490 17978
rect 9490 17926 9516 17978
rect 9220 17924 9276 17926
rect 9300 17924 9356 17926
rect 9380 17924 9436 17926
rect 9460 17924 9516 17926
rect 9220 16890 9276 16892
rect 9300 16890 9356 16892
rect 9380 16890 9436 16892
rect 9460 16890 9516 16892
rect 9220 16838 9246 16890
rect 9246 16838 9276 16890
rect 9300 16838 9310 16890
rect 9310 16838 9356 16890
rect 9380 16838 9426 16890
rect 9426 16838 9436 16890
rect 9460 16838 9490 16890
rect 9490 16838 9516 16890
rect 9220 16836 9276 16838
rect 9300 16836 9356 16838
rect 9380 16836 9436 16838
rect 9460 16836 9516 16838
rect 9220 15802 9276 15804
rect 9300 15802 9356 15804
rect 9380 15802 9436 15804
rect 9460 15802 9516 15804
rect 9220 15750 9246 15802
rect 9246 15750 9276 15802
rect 9300 15750 9310 15802
rect 9310 15750 9356 15802
rect 9380 15750 9426 15802
rect 9426 15750 9436 15802
rect 9460 15750 9490 15802
rect 9490 15750 9516 15802
rect 9220 15748 9276 15750
rect 9300 15748 9356 15750
rect 9380 15748 9436 15750
rect 9460 15748 9516 15750
rect 9220 14714 9276 14716
rect 9300 14714 9356 14716
rect 9380 14714 9436 14716
rect 9460 14714 9516 14716
rect 9220 14662 9246 14714
rect 9246 14662 9276 14714
rect 9300 14662 9310 14714
rect 9310 14662 9356 14714
rect 9380 14662 9426 14714
rect 9426 14662 9436 14714
rect 9460 14662 9490 14714
rect 9490 14662 9516 14714
rect 9220 14660 9276 14662
rect 9300 14660 9356 14662
rect 9380 14660 9436 14662
rect 9460 14660 9516 14662
rect 9220 13626 9276 13628
rect 9300 13626 9356 13628
rect 9380 13626 9436 13628
rect 9460 13626 9516 13628
rect 9220 13574 9246 13626
rect 9246 13574 9276 13626
rect 9300 13574 9310 13626
rect 9310 13574 9356 13626
rect 9380 13574 9426 13626
rect 9426 13574 9436 13626
rect 9460 13574 9490 13626
rect 9490 13574 9516 13626
rect 9220 13572 9276 13574
rect 9300 13572 9356 13574
rect 9380 13572 9436 13574
rect 9460 13572 9516 13574
rect 9220 12538 9276 12540
rect 9300 12538 9356 12540
rect 9380 12538 9436 12540
rect 9460 12538 9516 12540
rect 9220 12486 9246 12538
rect 9246 12486 9276 12538
rect 9300 12486 9310 12538
rect 9310 12486 9356 12538
rect 9380 12486 9426 12538
rect 9426 12486 9436 12538
rect 9460 12486 9490 12538
rect 9490 12486 9516 12538
rect 9220 12484 9276 12486
rect 9300 12484 9356 12486
rect 9380 12484 9436 12486
rect 9460 12484 9516 12486
rect 9220 11450 9276 11452
rect 9300 11450 9356 11452
rect 9380 11450 9436 11452
rect 9460 11450 9516 11452
rect 9220 11398 9246 11450
rect 9246 11398 9276 11450
rect 9300 11398 9310 11450
rect 9310 11398 9356 11450
rect 9380 11398 9426 11450
rect 9426 11398 9436 11450
rect 9460 11398 9490 11450
rect 9490 11398 9516 11450
rect 9220 11396 9276 11398
rect 9300 11396 9356 11398
rect 9380 11396 9436 11398
rect 9460 11396 9516 11398
rect 9220 10362 9276 10364
rect 9300 10362 9356 10364
rect 9380 10362 9436 10364
rect 9460 10362 9516 10364
rect 9220 10310 9246 10362
rect 9246 10310 9276 10362
rect 9300 10310 9310 10362
rect 9310 10310 9356 10362
rect 9380 10310 9426 10362
rect 9426 10310 9436 10362
rect 9460 10310 9490 10362
rect 9490 10310 9516 10362
rect 9220 10308 9276 10310
rect 9300 10308 9356 10310
rect 9380 10308 9436 10310
rect 9460 10308 9516 10310
rect 9220 9274 9276 9276
rect 9300 9274 9356 9276
rect 9380 9274 9436 9276
rect 9460 9274 9516 9276
rect 9220 9222 9246 9274
rect 9246 9222 9276 9274
rect 9300 9222 9310 9274
rect 9310 9222 9356 9274
rect 9380 9222 9426 9274
rect 9426 9222 9436 9274
rect 9460 9222 9490 9274
rect 9490 9222 9516 9274
rect 9220 9220 9276 9222
rect 9300 9220 9356 9222
rect 9380 9220 9436 9222
rect 9460 9220 9516 9222
rect 9220 8186 9276 8188
rect 9300 8186 9356 8188
rect 9380 8186 9436 8188
rect 9460 8186 9516 8188
rect 9220 8134 9246 8186
rect 9246 8134 9276 8186
rect 9300 8134 9310 8186
rect 9310 8134 9356 8186
rect 9380 8134 9426 8186
rect 9426 8134 9436 8186
rect 9460 8134 9490 8186
rect 9490 8134 9516 8186
rect 9220 8132 9276 8134
rect 9300 8132 9356 8134
rect 9380 8132 9436 8134
rect 9460 8132 9516 8134
rect 9220 7098 9276 7100
rect 9300 7098 9356 7100
rect 9380 7098 9436 7100
rect 9460 7098 9516 7100
rect 9220 7046 9246 7098
rect 9246 7046 9276 7098
rect 9300 7046 9310 7098
rect 9310 7046 9356 7098
rect 9380 7046 9426 7098
rect 9426 7046 9436 7098
rect 9460 7046 9490 7098
rect 9490 7046 9516 7098
rect 9220 7044 9276 7046
rect 9300 7044 9356 7046
rect 9380 7044 9436 7046
rect 9460 7044 9516 7046
rect 9220 6010 9276 6012
rect 9300 6010 9356 6012
rect 9380 6010 9436 6012
rect 9460 6010 9516 6012
rect 9220 5958 9246 6010
rect 9246 5958 9276 6010
rect 9300 5958 9310 6010
rect 9310 5958 9356 6010
rect 9380 5958 9426 6010
rect 9426 5958 9436 6010
rect 9460 5958 9490 6010
rect 9490 5958 9516 6010
rect 9220 5956 9276 5958
rect 9300 5956 9356 5958
rect 9380 5956 9436 5958
rect 9460 5956 9516 5958
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 9220 4922 9276 4924
rect 9300 4922 9356 4924
rect 9380 4922 9436 4924
rect 9460 4922 9516 4924
rect 9220 4870 9246 4922
rect 9246 4870 9276 4922
rect 9300 4870 9310 4922
rect 9310 4870 9356 4922
rect 9380 4870 9426 4922
rect 9426 4870 9436 4922
rect 9460 4870 9490 4922
rect 9490 4870 9516 4922
rect 9220 4868 9276 4870
rect 9300 4868 9356 4870
rect 9380 4868 9436 4870
rect 9460 4868 9516 4870
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 9220 3834 9276 3836
rect 9300 3834 9356 3836
rect 9380 3834 9436 3836
rect 9460 3834 9516 3836
rect 9220 3782 9246 3834
rect 9246 3782 9276 3834
rect 9300 3782 9310 3834
rect 9310 3782 9356 3834
rect 9380 3782 9426 3834
rect 9426 3782 9436 3834
rect 9460 3782 9490 3834
rect 9490 3782 9516 3834
rect 9220 3780 9276 3782
rect 9300 3780 9356 3782
rect 9380 3780 9436 3782
rect 9460 3780 9516 3782
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 14220 42458 14276 42460
rect 14300 42458 14356 42460
rect 14380 42458 14436 42460
rect 14460 42458 14516 42460
rect 14220 42406 14246 42458
rect 14246 42406 14276 42458
rect 14300 42406 14310 42458
rect 14310 42406 14356 42458
rect 14380 42406 14426 42458
rect 14426 42406 14436 42458
rect 14460 42406 14490 42458
rect 14490 42406 14516 42458
rect 14220 42404 14276 42406
rect 14300 42404 14356 42406
rect 14380 42404 14436 42406
rect 14460 42404 14516 42406
rect 14220 41370 14276 41372
rect 14300 41370 14356 41372
rect 14380 41370 14436 41372
rect 14460 41370 14516 41372
rect 14220 41318 14246 41370
rect 14246 41318 14276 41370
rect 14300 41318 14310 41370
rect 14310 41318 14356 41370
rect 14380 41318 14426 41370
rect 14426 41318 14436 41370
rect 14460 41318 14490 41370
rect 14490 41318 14516 41370
rect 14220 41316 14276 41318
rect 14300 41316 14356 41318
rect 14380 41316 14436 41318
rect 14460 41316 14516 41318
rect 14220 40282 14276 40284
rect 14300 40282 14356 40284
rect 14380 40282 14436 40284
rect 14460 40282 14516 40284
rect 14220 40230 14246 40282
rect 14246 40230 14276 40282
rect 14300 40230 14310 40282
rect 14310 40230 14356 40282
rect 14380 40230 14426 40282
rect 14426 40230 14436 40282
rect 14460 40230 14490 40282
rect 14490 40230 14516 40282
rect 14220 40228 14276 40230
rect 14300 40228 14356 40230
rect 14380 40228 14436 40230
rect 14460 40228 14516 40230
rect 14220 39194 14276 39196
rect 14300 39194 14356 39196
rect 14380 39194 14436 39196
rect 14460 39194 14516 39196
rect 14220 39142 14246 39194
rect 14246 39142 14276 39194
rect 14300 39142 14310 39194
rect 14310 39142 14356 39194
rect 14380 39142 14426 39194
rect 14426 39142 14436 39194
rect 14460 39142 14490 39194
rect 14490 39142 14516 39194
rect 14220 39140 14276 39142
rect 14300 39140 14356 39142
rect 14380 39140 14436 39142
rect 14460 39140 14516 39142
rect 14220 38106 14276 38108
rect 14300 38106 14356 38108
rect 14380 38106 14436 38108
rect 14460 38106 14516 38108
rect 14220 38054 14246 38106
rect 14246 38054 14276 38106
rect 14300 38054 14310 38106
rect 14310 38054 14356 38106
rect 14380 38054 14426 38106
rect 14426 38054 14436 38106
rect 14460 38054 14490 38106
rect 14490 38054 14516 38106
rect 14220 38052 14276 38054
rect 14300 38052 14356 38054
rect 14380 38052 14436 38054
rect 14460 38052 14516 38054
rect 14220 37018 14276 37020
rect 14300 37018 14356 37020
rect 14380 37018 14436 37020
rect 14460 37018 14516 37020
rect 14220 36966 14246 37018
rect 14246 36966 14276 37018
rect 14300 36966 14310 37018
rect 14310 36966 14356 37018
rect 14380 36966 14426 37018
rect 14426 36966 14436 37018
rect 14460 36966 14490 37018
rect 14490 36966 14516 37018
rect 14220 36964 14276 36966
rect 14300 36964 14356 36966
rect 14380 36964 14436 36966
rect 14460 36964 14516 36966
rect 14220 35930 14276 35932
rect 14300 35930 14356 35932
rect 14380 35930 14436 35932
rect 14460 35930 14516 35932
rect 14220 35878 14246 35930
rect 14246 35878 14276 35930
rect 14300 35878 14310 35930
rect 14310 35878 14356 35930
rect 14380 35878 14426 35930
rect 14426 35878 14436 35930
rect 14460 35878 14490 35930
rect 14490 35878 14516 35930
rect 14220 35876 14276 35878
rect 14300 35876 14356 35878
rect 14380 35876 14436 35878
rect 14460 35876 14516 35878
rect 14220 34842 14276 34844
rect 14300 34842 14356 34844
rect 14380 34842 14436 34844
rect 14460 34842 14516 34844
rect 14220 34790 14246 34842
rect 14246 34790 14276 34842
rect 14300 34790 14310 34842
rect 14310 34790 14356 34842
rect 14380 34790 14426 34842
rect 14426 34790 14436 34842
rect 14460 34790 14490 34842
rect 14490 34790 14516 34842
rect 14220 34788 14276 34790
rect 14300 34788 14356 34790
rect 14380 34788 14436 34790
rect 14460 34788 14516 34790
rect 14220 33754 14276 33756
rect 14300 33754 14356 33756
rect 14380 33754 14436 33756
rect 14460 33754 14516 33756
rect 14220 33702 14246 33754
rect 14246 33702 14276 33754
rect 14300 33702 14310 33754
rect 14310 33702 14356 33754
rect 14380 33702 14426 33754
rect 14426 33702 14436 33754
rect 14460 33702 14490 33754
rect 14490 33702 14516 33754
rect 14220 33700 14276 33702
rect 14300 33700 14356 33702
rect 14380 33700 14436 33702
rect 14460 33700 14516 33702
rect 14220 32666 14276 32668
rect 14300 32666 14356 32668
rect 14380 32666 14436 32668
rect 14460 32666 14516 32668
rect 14220 32614 14246 32666
rect 14246 32614 14276 32666
rect 14300 32614 14310 32666
rect 14310 32614 14356 32666
rect 14380 32614 14426 32666
rect 14426 32614 14436 32666
rect 14460 32614 14490 32666
rect 14490 32614 14516 32666
rect 14220 32612 14276 32614
rect 14300 32612 14356 32614
rect 14380 32612 14436 32614
rect 14460 32612 14516 32614
rect 14220 31578 14276 31580
rect 14300 31578 14356 31580
rect 14380 31578 14436 31580
rect 14460 31578 14516 31580
rect 14220 31526 14246 31578
rect 14246 31526 14276 31578
rect 14300 31526 14310 31578
rect 14310 31526 14356 31578
rect 14380 31526 14426 31578
rect 14426 31526 14436 31578
rect 14460 31526 14490 31578
rect 14490 31526 14516 31578
rect 14220 31524 14276 31526
rect 14300 31524 14356 31526
rect 14380 31524 14436 31526
rect 14460 31524 14516 31526
rect 14220 30490 14276 30492
rect 14300 30490 14356 30492
rect 14380 30490 14436 30492
rect 14460 30490 14516 30492
rect 14220 30438 14246 30490
rect 14246 30438 14276 30490
rect 14300 30438 14310 30490
rect 14310 30438 14356 30490
rect 14380 30438 14426 30490
rect 14426 30438 14436 30490
rect 14460 30438 14490 30490
rect 14490 30438 14516 30490
rect 14220 30436 14276 30438
rect 14300 30436 14356 30438
rect 14380 30436 14436 30438
rect 14460 30436 14516 30438
rect 14220 29402 14276 29404
rect 14300 29402 14356 29404
rect 14380 29402 14436 29404
rect 14460 29402 14516 29404
rect 14220 29350 14246 29402
rect 14246 29350 14276 29402
rect 14300 29350 14310 29402
rect 14310 29350 14356 29402
rect 14380 29350 14426 29402
rect 14426 29350 14436 29402
rect 14460 29350 14490 29402
rect 14490 29350 14516 29402
rect 14220 29348 14276 29350
rect 14300 29348 14356 29350
rect 14380 29348 14436 29350
rect 14460 29348 14516 29350
rect 14220 28314 14276 28316
rect 14300 28314 14356 28316
rect 14380 28314 14436 28316
rect 14460 28314 14516 28316
rect 14220 28262 14246 28314
rect 14246 28262 14276 28314
rect 14300 28262 14310 28314
rect 14310 28262 14356 28314
rect 14380 28262 14426 28314
rect 14426 28262 14436 28314
rect 14460 28262 14490 28314
rect 14490 28262 14516 28314
rect 14220 28260 14276 28262
rect 14300 28260 14356 28262
rect 14380 28260 14436 28262
rect 14460 28260 14516 28262
rect 14220 27226 14276 27228
rect 14300 27226 14356 27228
rect 14380 27226 14436 27228
rect 14460 27226 14516 27228
rect 14220 27174 14246 27226
rect 14246 27174 14276 27226
rect 14300 27174 14310 27226
rect 14310 27174 14356 27226
rect 14380 27174 14426 27226
rect 14426 27174 14436 27226
rect 14460 27174 14490 27226
rect 14490 27174 14516 27226
rect 14220 27172 14276 27174
rect 14300 27172 14356 27174
rect 14380 27172 14436 27174
rect 14460 27172 14516 27174
rect 14220 26138 14276 26140
rect 14300 26138 14356 26140
rect 14380 26138 14436 26140
rect 14460 26138 14516 26140
rect 14220 26086 14246 26138
rect 14246 26086 14276 26138
rect 14300 26086 14310 26138
rect 14310 26086 14356 26138
rect 14380 26086 14426 26138
rect 14426 26086 14436 26138
rect 14460 26086 14490 26138
rect 14490 26086 14516 26138
rect 14220 26084 14276 26086
rect 14300 26084 14356 26086
rect 14380 26084 14436 26086
rect 14460 26084 14516 26086
rect 14220 25050 14276 25052
rect 14300 25050 14356 25052
rect 14380 25050 14436 25052
rect 14460 25050 14516 25052
rect 14220 24998 14246 25050
rect 14246 24998 14276 25050
rect 14300 24998 14310 25050
rect 14310 24998 14356 25050
rect 14380 24998 14426 25050
rect 14426 24998 14436 25050
rect 14460 24998 14490 25050
rect 14490 24998 14516 25050
rect 14220 24996 14276 24998
rect 14300 24996 14356 24998
rect 14380 24996 14436 24998
rect 14460 24996 14516 24998
rect 14220 23962 14276 23964
rect 14300 23962 14356 23964
rect 14380 23962 14436 23964
rect 14460 23962 14516 23964
rect 14220 23910 14246 23962
rect 14246 23910 14276 23962
rect 14300 23910 14310 23962
rect 14310 23910 14356 23962
rect 14380 23910 14426 23962
rect 14426 23910 14436 23962
rect 14460 23910 14490 23962
rect 14490 23910 14516 23962
rect 14220 23908 14276 23910
rect 14300 23908 14356 23910
rect 14380 23908 14436 23910
rect 14460 23908 14516 23910
rect 14220 22874 14276 22876
rect 14300 22874 14356 22876
rect 14380 22874 14436 22876
rect 14460 22874 14516 22876
rect 14220 22822 14246 22874
rect 14246 22822 14276 22874
rect 14300 22822 14310 22874
rect 14310 22822 14356 22874
rect 14380 22822 14426 22874
rect 14426 22822 14436 22874
rect 14460 22822 14490 22874
rect 14490 22822 14516 22874
rect 14220 22820 14276 22822
rect 14300 22820 14356 22822
rect 14380 22820 14436 22822
rect 14460 22820 14516 22822
rect 14220 21786 14276 21788
rect 14300 21786 14356 21788
rect 14380 21786 14436 21788
rect 14460 21786 14516 21788
rect 14220 21734 14246 21786
rect 14246 21734 14276 21786
rect 14300 21734 14310 21786
rect 14310 21734 14356 21786
rect 14380 21734 14426 21786
rect 14426 21734 14436 21786
rect 14460 21734 14490 21786
rect 14490 21734 14516 21786
rect 14220 21732 14276 21734
rect 14300 21732 14356 21734
rect 14380 21732 14436 21734
rect 14460 21732 14516 21734
rect 14220 20698 14276 20700
rect 14300 20698 14356 20700
rect 14380 20698 14436 20700
rect 14460 20698 14516 20700
rect 14220 20646 14246 20698
rect 14246 20646 14276 20698
rect 14300 20646 14310 20698
rect 14310 20646 14356 20698
rect 14380 20646 14426 20698
rect 14426 20646 14436 20698
rect 14460 20646 14490 20698
rect 14490 20646 14516 20698
rect 14220 20644 14276 20646
rect 14300 20644 14356 20646
rect 14380 20644 14436 20646
rect 14460 20644 14516 20646
rect 14220 19610 14276 19612
rect 14300 19610 14356 19612
rect 14380 19610 14436 19612
rect 14460 19610 14516 19612
rect 14220 19558 14246 19610
rect 14246 19558 14276 19610
rect 14300 19558 14310 19610
rect 14310 19558 14356 19610
rect 14380 19558 14426 19610
rect 14426 19558 14436 19610
rect 14460 19558 14490 19610
rect 14490 19558 14516 19610
rect 14220 19556 14276 19558
rect 14300 19556 14356 19558
rect 14380 19556 14436 19558
rect 14460 19556 14516 19558
rect 14220 18522 14276 18524
rect 14300 18522 14356 18524
rect 14380 18522 14436 18524
rect 14460 18522 14516 18524
rect 14220 18470 14246 18522
rect 14246 18470 14276 18522
rect 14300 18470 14310 18522
rect 14310 18470 14356 18522
rect 14380 18470 14426 18522
rect 14426 18470 14436 18522
rect 14460 18470 14490 18522
rect 14490 18470 14516 18522
rect 14220 18468 14276 18470
rect 14300 18468 14356 18470
rect 14380 18468 14436 18470
rect 14460 18468 14516 18470
rect 14220 17434 14276 17436
rect 14300 17434 14356 17436
rect 14380 17434 14436 17436
rect 14460 17434 14516 17436
rect 14220 17382 14246 17434
rect 14246 17382 14276 17434
rect 14300 17382 14310 17434
rect 14310 17382 14356 17434
rect 14380 17382 14426 17434
rect 14426 17382 14436 17434
rect 14460 17382 14490 17434
rect 14490 17382 14516 17434
rect 14220 17380 14276 17382
rect 14300 17380 14356 17382
rect 14380 17380 14436 17382
rect 14460 17380 14516 17382
rect 14220 16346 14276 16348
rect 14300 16346 14356 16348
rect 14380 16346 14436 16348
rect 14460 16346 14516 16348
rect 14220 16294 14246 16346
rect 14246 16294 14276 16346
rect 14300 16294 14310 16346
rect 14310 16294 14356 16346
rect 14380 16294 14426 16346
rect 14426 16294 14436 16346
rect 14460 16294 14490 16346
rect 14490 16294 14516 16346
rect 14220 16292 14276 16294
rect 14300 16292 14356 16294
rect 14380 16292 14436 16294
rect 14460 16292 14516 16294
rect 14220 15258 14276 15260
rect 14300 15258 14356 15260
rect 14380 15258 14436 15260
rect 14460 15258 14516 15260
rect 14220 15206 14246 15258
rect 14246 15206 14276 15258
rect 14300 15206 14310 15258
rect 14310 15206 14356 15258
rect 14380 15206 14426 15258
rect 14426 15206 14436 15258
rect 14460 15206 14490 15258
rect 14490 15206 14516 15258
rect 14220 15204 14276 15206
rect 14300 15204 14356 15206
rect 14380 15204 14436 15206
rect 14460 15204 14516 15206
rect 14220 14170 14276 14172
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14220 14118 14246 14170
rect 14246 14118 14276 14170
rect 14300 14118 14310 14170
rect 14310 14118 14356 14170
rect 14380 14118 14426 14170
rect 14426 14118 14436 14170
rect 14460 14118 14490 14170
rect 14490 14118 14516 14170
rect 14220 14116 14276 14118
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 24220 46810 24276 46812
rect 24300 46810 24356 46812
rect 24380 46810 24436 46812
rect 24460 46810 24516 46812
rect 24220 46758 24246 46810
rect 24246 46758 24276 46810
rect 24300 46758 24310 46810
rect 24310 46758 24356 46810
rect 24380 46758 24426 46810
rect 24426 46758 24436 46810
rect 24460 46758 24490 46810
rect 24490 46758 24516 46810
rect 24220 46756 24276 46758
rect 24300 46756 24356 46758
rect 24380 46756 24436 46758
rect 24460 46756 24516 46758
rect 34220 46810 34276 46812
rect 34300 46810 34356 46812
rect 34380 46810 34436 46812
rect 34460 46810 34516 46812
rect 34220 46758 34246 46810
rect 34246 46758 34276 46810
rect 34300 46758 34310 46810
rect 34310 46758 34356 46810
rect 34380 46758 34426 46810
rect 34426 46758 34436 46810
rect 34460 46758 34490 46810
rect 34490 46758 34516 46810
rect 34220 46756 34276 46758
rect 34300 46756 34356 46758
rect 34380 46756 34436 46758
rect 34460 46756 34516 46758
rect 44220 46810 44276 46812
rect 44300 46810 44356 46812
rect 44380 46810 44436 46812
rect 44460 46810 44516 46812
rect 44220 46758 44246 46810
rect 44246 46758 44276 46810
rect 44300 46758 44310 46810
rect 44310 46758 44356 46810
rect 44380 46758 44426 46810
rect 44426 46758 44436 46810
rect 44460 46758 44490 46810
rect 44490 46758 44516 46810
rect 44220 46756 44276 46758
rect 44300 46756 44356 46758
rect 44380 46756 44436 46758
rect 44460 46756 44516 46758
rect 19220 46266 19276 46268
rect 19300 46266 19356 46268
rect 19380 46266 19436 46268
rect 19460 46266 19516 46268
rect 19220 46214 19246 46266
rect 19246 46214 19276 46266
rect 19300 46214 19310 46266
rect 19310 46214 19356 46266
rect 19380 46214 19426 46266
rect 19426 46214 19436 46266
rect 19460 46214 19490 46266
rect 19490 46214 19516 46266
rect 19220 46212 19276 46214
rect 19300 46212 19356 46214
rect 19380 46212 19436 46214
rect 19460 46212 19516 46214
rect 29220 46266 29276 46268
rect 29300 46266 29356 46268
rect 29380 46266 29436 46268
rect 29460 46266 29516 46268
rect 29220 46214 29246 46266
rect 29246 46214 29276 46266
rect 29300 46214 29310 46266
rect 29310 46214 29356 46266
rect 29380 46214 29426 46266
rect 29426 46214 29436 46266
rect 29460 46214 29490 46266
rect 29490 46214 29516 46266
rect 29220 46212 29276 46214
rect 29300 46212 29356 46214
rect 29380 46212 29436 46214
rect 29460 46212 29516 46214
rect 39220 46266 39276 46268
rect 39300 46266 39356 46268
rect 39380 46266 39436 46268
rect 39460 46266 39516 46268
rect 39220 46214 39246 46266
rect 39246 46214 39276 46266
rect 39300 46214 39310 46266
rect 39310 46214 39356 46266
rect 39380 46214 39426 46266
rect 39426 46214 39436 46266
rect 39460 46214 39490 46266
rect 39490 46214 39516 46266
rect 39220 46212 39276 46214
rect 39300 46212 39356 46214
rect 39380 46212 39436 46214
rect 39460 46212 39516 46214
rect 24220 45722 24276 45724
rect 24300 45722 24356 45724
rect 24380 45722 24436 45724
rect 24460 45722 24516 45724
rect 24220 45670 24246 45722
rect 24246 45670 24276 45722
rect 24300 45670 24310 45722
rect 24310 45670 24356 45722
rect 24380 45670 24426 45722
rect 24426 45670 24436 45722
rect 24460 45670 24490 45722
rect 24490 45670 24516 45722
rect 24220 45668 24276 45670
rect 24300 45668 24356 45670
rect 24380 45668 24436 45670
rect 24460 45668 24516 45670
rect 34220 45722 34276 45724
rect 34300 45722 34356 45724
rect 34380 45722 34436 45724
rect 34460 45722 34516 45724
rect 34220 45670 34246 45722
rect 34246 45670 34276 45722
rect 34300 45670 34310 45722
rect 34310 45670 34356 45722
rect 34380 45670 34426 45722
rect 34426 45670 34436 45722
rect 34460 45670 34490 45722
rect 34490 45670 34516 45722
rect 34220 45668 34276 45670
rect 34300 45668 34356 45670
rect 34380 45668 34436 45670
rect 34460 45668 34516 45670
rect 44220 45722 44276 45724
rect 44300 45722 44356 45724
rect 44380 45722 44436 45724
rect 44460 45722 44516 45724
rect 44220 45670 44246 45722
rect 44246 45670 44276 45722
rect 44300 45670 44310 45722
rect 44310 45670 44356 45722
rect 44380 45670 44426 45722
rect 44426 45670 44436 45722
rect 44460 45670 44490 45722
rect 44490 45670 44516 45722
rect 44220 45668 44276 45670
rect 44300 45668 44356 45670
rect 44380 45668 44436 45670
rect 44460 45668 44516 45670
rect 19220 45178 19276 45180
rect 19300 45178 19356 45180
rect 19380 45178 19436 45180
rect 19460 45178 19516 45180
rect 19220 45126 19246 45178
rect 19246 45126 19276 45178
rect 19300 45126 19310 45178
rect 19310 45126 19356 45178
rect 19380 45126 19426 45178
rect 19426 45126 19436 45178
rect 19460 45126 19490 45178
rect 19490 45126 19516 45178
rect 19220 45124 19276 45126
rect 19300 45124 19356 45126
rect 19380 45124 19436 45126
rect 19460 45124 19516 45126
rect 19220 44090 19276 44092
rect 19300 44090 19356 44092
rect 19380 44090 19436 44092
rect 19460 44090 19516 44092
rect 19220 44038 19246 44090
rect 19246 44038 19276 44090
rect 19300 44038 19310 44090
rect 19310 44038 19356 44090
rect 19380 44038 19426 44090
rect 19426 44038 19436 44090
rect 19460 44038 19490 44090
rect 19490 44038 19516 44090
rect 19220 44036 19276 44038
rect 19300 44036 19356 44038
rect 19380 44036 19436 44038
rect 19460 44036 19516 44038
rect 19220 43002 19276 43004
rect 19300 43002 19356 43004
rect 19380 43002 19436 43004
rect 19460 43002 19516 43004
rect 19220 42950 19246 43002
rect 19246 42950 19276 43002
rect 19300 42950 19310 43002
rect 19310 42950 19356 43002
rect 19380 42950 19426 43002
rect 19426 42950 19436 43002
rect 19460 42950 19490 43002
rect 19490 42950 19516 43002
rect 19220 42948 19276 42950
rect 19300 42948 19356 42950
rect 19380 42948 19436 42950
rect 19460 42948 19516 42950
rect 19220 41914 19276 41916
rect 19300 41914 19356 41916
rect 19380 41914 19436 41916
rect 19460 41914 19516 41916
rect 19220 41862 19246 41914
rect 19246 41862 19276 41914
rect 19300 41862 19310 41914
rect 19310 41862 19356 41914
rect 19380 41862 19426 41914
rect 19426 41862 19436 41914
rect 19460 41862 19490 41914
rect 19490 41862 19516 41914
rect 19220 41860 19276 41862
rect 19300 41860 19356 41862
rect 19380 41860 19436 41862
rect 19460 41860 19516 41862
rect 19220 40826 19276 40828
rect 19300 40826 19356 40828
rect 19380 40826 19436 40828
rect 19460 40826 19516 40828
rect 19220 40774 19246 40826
rect 19246 40774 19276 40826
rect 19300 40774 19310 40826
rect 19310 40774 19356 40826
rect 19380 40774 19426 40826
rect 19426 40774 19436 40826
rect 19460 40774 19490 40826
rect 19490 40774 19516 40826
rect 19220 40772 19276 40774
rect 19300 40772 19356 40774
rect 19380 40772 19436 40774
rect 19460 40772 19516 40774
rect 19220 39738 19276 39740
rect 19300 39738 19356 39740
rect 19380 39738 19436 39740
rect 19460 39738 19516 39740
rect 19220 39686 19246 39738
rect 19246 39686 19276 39738
rect 19300 39686 19310 39738
rect 19310 39686 19356 39738
rect 19380 39686 19426 39738
rect 19426 39686 19436 39738
rect 19460 39686 19490 39738
rect 19490 39686 19516 39738
rect 19220 39684 19276 39686
rect 19300 39684 19356 39686
rect 19380 39684 19436 39686
rect 19460 39684 19516 39686
rect 19220 38650 19276 38652
rect 19300 38650 19356 38652
rect 19380 38650 19436 38652
rect 19460 38650 19516 38652
rect 19220 38598 19246 38650
rect 19246 38598 19276 38650
rect 19300 38598 19310 38650
rect 19310 38598 19356 38650
rect 19380 38598 19426 38650
rect 19426 38598 19436 38650
rect 19460 38598 19490 38650
rect 19490 38598 19516 38650
rect 19220 38596 19276 38598
rect 19300 38596 19356 38598
rect 19380 38596 19436 38598
rect 19460 38596 19516 38598
rect 19220 37562 19276 37564
rect 19300 37562 19356 37564
rect 19380 37562 19436 37564
rect 19460 37562 19516 37564
rect 19220 37510 19246 37562
rect 19246 37510 19276 37562
rect 19300 37510 19310 37562
rect 19310 37510 19356 37562
rect 19380 37510 19426 37562
rect 19426 37510 19436 37562
rect 19460 37510 19490 37562
rect 19490 37510 19516 37562
rect 19220 37508 19276 37510
rect 19300 37508 19356 37510
rect 19380 37508 19436 37510
rect 19460 37508 19516 37510
rect 24220 44634 24276 44636
rect 24300 44634 24356 44636
rect 24380 44634 24436 44636
rect 24460 44634 24516 44636
rect 24220 44582 24246 44634
rect 24246 44582 24276 44634
rect 24300 44582 24310 44634
rect 24310 44582 24356 44634
rect 24380 44582 24426 44634
rect 24426 44582 24436 44634
rect 24460 44582 24490 44634
rect 24490 44582 24516 44634
rect 24220 44580 24276 44582
rect 24300 44580 24356 44582
rect 24380 44580 24436 44582
rect 24460 44580 24516 44582
rect 24220 43546 24276 43548
rect 24300 43546 24356 43548
rect 24380 43546 24436 43548
rect 24460 43546 24516 43548
rect 24220 43494 24246 43546
rect 24246 43494 24276 43546
rect 24300 43494 24310 43546
rect 24310 43494 24356 43546
rect 24380 43494 24426 43546
rect 24426 43494 24436 43546
rect 24460 43494 24490 43546
rect 24490 43494 24516 43546
rect 24220 43492 24276 43494
rect 24300 43492 24356 43494
rect 24380 43492 24436 43494
rect 24460 43492 24516 43494
rect 24220 42458 24276 42460
rect 24300 42458 24356 42460
rect 24380 42458 24436 42460
rect 24460 42458 24516 42460
rect 24220 42406 24246 42458
rect 24246 42406 24276 42458
rect 24300 42406 24310 42458
rect 24310 42406 24356 42458
rect 24380 42406 24426 42458
rect 24426 42406 24436 42458
rect 24460 42406 24490 42458
rect 24490 42406 24516 42458
rect 24220 42404 24276 42406
rect 24300 42404 24356 42406
rect 24380 42404 24436 42406
rect 24460 42404 24516 42406
rect 24220 41370 24276 41372
rect 24300 41370 24356 41372
rect 24380 41370 24436 41372
rect 24460 41370 24516 41372
rect 24220 41318 24246 41370
rect 24246 41318 24276 41370
rect 24300 41318 24310 41370
rect 24310 41318 24356 41370
rect 24380 41318 24426 41370
rect 24426 41318 24436 41370
rect 24460 41318 24490 41370
rect 24490 41318 24516 41370
rect 24220 41316 24276 41318
rect 24300 41316 24356 41318
rect 24380 41316 24436 41318
rect 24460 41316 24516 41318
rect 24220 40282 24276 40284
rect 24300 40282 24356 40284
rect 24380 40282 24436 40284
rect 24460 40282 24516 40284
rect 24220 40230 24246 40282
rect 24246 40230 24276 40282
rect 24300 40230 24310 40282
rect 24310 40230 24356 40282
rect 24380 40230 24426 40282
rect 24426 40230 24436 40282
rect 24460 40230 24490 40282
rect 24490 40230 24516 40282
rect 24220 40228 24276 40230
rect 24300 40228 24356 40230
rect 24380 40228 24436 40230
rect 24460 40228 24516 40230
rect 19220 36474 19276 36476
rect 19300 36474 19356 36476
rect 19380 36474 19436 36476
rect 19460 36474 19516 36476
rect 19220 36422 19246 36474
rect 19246 36422 19276 36474
rect 19300 36422 19310 36474
rect 19310 36422 19356 36474
rect 19380 36422 19426 36474
rect 19426 36422 19436 36474
rect 19460 36422 19490 36474
rect 19490 36422 19516 36474
rect 19220 36420 19276 36422
rect 19300 36420 19356 36422
rect 19380 36420 19436 36422
rect 19460 36420 19516 36422
rect 19220 35386 19276 35388
rect 19300 35386 19356 35388
rect 19380 35386 19436 35388
rect 19460 35386 19516 35388
rect 19220 35334 19246 35386
rect 19246 35334 19276 35386
rect 19300 35334 19310 35386
rect 19310 35334 19356 35386
rect 19380 35334 19426 35386
rect 19426 35334 19436 35386
rect 19460 35334 19490 35386
rect 19490 35334 19516 35386
rect 19220 35332 19276 35334
rect 19300 35332 19356 35334
rect 19380 35332 19436 35334
rect 19460 35332 19516 35334
rect 19220 34298 19276 34300
rect 19300 34298 19356 34300
rect 19380 34298 19436 34300
rect 19460 34298 19516 34300
rect 19220 34246 19246 34298
rect 19246 34246 19276 34298
rect 19300 34246 19310 34298
rect 19310 34246 19356 34298
rect 19380 34246 19426 34298
rect 19426 34246 19436 34298
rect 19460 34246 19490 34298
rect 19490 34246 19516 34298
rect 19220 34244 19276 34246
rect 19300 34244 19356 34246
rect 19380 34244 19436 34246
rect 19460 34244 19516 34246
rect 14220 13082 14276 13084
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14220 13030 14246 13082
rect 14246 13030 14276 13082
rect 14300 13030 14310 13082
rect 14310 13030 14356 13082
rect 14380 13030 14426 13082
rect 14426 13030 14436 13082
rect 14460 13030 14490 13082
rect 14490 13030 14516 13082
rect 14220 13028 14276 13030
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14220 11994 14276 11996
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14220 11942 14246 11994
rect 14246 11942 14276 11994
rect 14300 11942 14310 11994
rect 14310 11942 14356 11994
rect 14380 11942 14426 11994
rect 14426 11942 14436 11994
rect 14460 11942 14490 11994
rect 14490 11942 14516 11994
rect 14220 11940 14276 11942
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14220 10906 14276 10908
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14220 10854 14246 10906
rect 14246 10854 14276 10906
rect 14300 10854 14310 10906
rect 14310 10854 14356 10906
rect 14380 10854 14426 10906
rect 14426 10854 14436 10906
rect 14460 10854 14490 10906
rect 14490 10854 14516 10906
rect 14220 10852 14276 10854
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14220 9818 14276 9820
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14220 9766 14246 9818
rect 14246 9766 14276 9818
rect 14300 9766 14310 9818
rect 14310 9766 14356 9818
rect 14380 9766 14426 9818
rect 14426 9766 14436 9818
rect 14460 9766 14490 9818
rect 14490 9766 14516 9818
rect 14220 9764 14276 9766
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14220 8730 14276 8732
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14220 8678 14246 8730
rect 14246 8678 14276 8730
rect 14300 8678 14310 8730
rect 14310 8678 14356 8730
rect 14380 8678 14426 8730
rect 14426 8678 14436 8730
rect 14460 8678 14490 8730
rect 14490 8678 14516 8730
rect 14220 8676 14276 8678
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14220 7642 14276 7644
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14220 7590 14246 7642
rect 14246 7590 14276 7642
rect 14300 7590 14310 7642
rect 14310 7590 14356 7642
rect 14380 7590 14426 7642
rect 14426 7590 14436 7642
rect 14460 7590 14490 7642
rect 14490 7590 14516 7642
rect 14220 7588 14276 7590
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14220 6554 14276 6556
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14220 6502 14246 6554
rect 14246 6502 14276 6554
rect 14300 6502 14310 6554
rect 14310 6502 14356 6554
rect 14380 6502 14426 6554
rect 14426 6502 14436 6554
rect 14460 6502 14490 6554
rect 14490 6502 14516 6554
rect 14220 6500 14276 6502
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 16026 11056 16082 11112
rect 18050 6976 18106 7032
rect 14220 5466 14276 5468
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14220 5414 14246 5466
rect 14246 5414 14276 5466
rect 14300 5414 14310 5466
rect 14310 5414 14356 5466
rect 14380 5414 14426 5466
rect 14426 5414 14436 5466
rect 14460 5414 14490 5466
rect 14490 5414 14516 5466
rect 14220 5412 14276 5414
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 19220 33210 19276 33212
rect 19300 33210 19356 33212
rect 19380 33210 19436 33212
rect 19460 33210 19516 33212
rect 19220 33158 19246 33210
rect 19246 33158 19276 33210
rect 19300 33158 19310 33210
rect 19310 33158 19356 33210
rect 19380 33158 19426 33210
rect 19426 33158 19436 33210
rect 19460 33158 19490 33210
rect 19490 33158 19516 33210
rect 19220 33156 19276 33158
rect 19300 33156 19356 33158
rect 19380 33156 19436 33158
rect 19460 33156 19516 33158
rect 19220 32122 19276 32124
rect 19300 32122 19356 32124
rect 19380 32122 19436 32124
rect 19460 32122 19516 32124
rect 19220 32070 19246 32122
rect 19246 32070 19276 32122
rect 19300 32070 19310 32122
rect 19310 32070 19356 32122
rect 19380 32070 19426 32122
rect 19426 32070 19436 32122
rect 19460 32070 19490 32122
rect 19490 32070 19516 32122
rect 19220 32068 19276 32070
rect 19300 32068 19356 32070
rect 19380 32068 19436 32070
rect 19460 32068 19516 32070
rect 19220 31034 19276 31036
rect 19300 31034 19356 31036
rect 19380 31034 19436 31036
rect 19460 31034 19516 31036
rect 19220 30982 19246 31034
rect 19246 30982 19276 31034
rect 19300 30982 19310 31034
rect 19310 30982 19356 31034
rect 19380 30982 19426 31034
rect 19426 30982 19436 31034
rect 19460 30982 19490 31034
rect 19490 30982 19516 31034
rect 19220 30980 19276 30982
rect 19300 30980 19356 30982
rect 19380 30980 19436 30982
rect 19460 30980 19516 30982
rect 19220 29946 19276 29948
rect 19300 29946 19356 29948
rect 19380 29946 19436 29948
rect 19460 29946 19516 29948
rect 19220 29894 19246 29946
rect 19246 29894 19276 29946
rect 19300 29894 19310 29946
rect 19310 29894 19356 29946
rect 19380 29894 19426 29946
rect 19426 29894 19436 29946
rect 19460 29894 19490 29946
rect 19490 29894 19516 29946
rect 19220 29892 19276 29894
rect 19300 29892 19356 29894
rect 19380 29892 19436 29894
rect 19460 29892 19516 29894
rect 19220 28858 19276 28860
rect 19300 28858 19356 28860
rect 19380 28858 19436 28860
rect 19460 28858 19516 28860
rect 19220 28806 19246 28858
rect 19246 28806 19276 28858
rect 19300 28806 19310 28858
rect 19310 28806 19356 28858
rect 19380 28806 19426 28858
rect 19426 28806 19436 28858
rect 19460 28806 19490 28858
rect 19490 28806 19516 28858
rect 19220 28804 19276 28806
rect 19300 28804 19356 28806
rect 19380 28804 19436 28806
rect 19460 28804 19516 28806
rect 19220 27770 19276 27772
rect 19300 27770 19356 27772
rect 19380 27770 19436 27772
rect 19460 27770 19516 27772
rect 19220 27718 19246 27770
rect 19246 27718 19276 27770
rect 19300 27718 19310 27770
rect 19310 27718 19356 27770
rect 19380 27718 19426 27770
rect 19426 27718 19436 27770
rect 19460 27718 19490 27770
rect 19490 27718 19516 27770
rect 19220 27716 19276 27718
rect 19300 27716 19356 27718
rect 19380 27716 19436 27718
rect 19460 27716 19516 27718
rect 19220 26682 19276 26684
rect 19300 26682 19356 26684
rect 19380 26682 19436 26684
rect 19460 26682 19516 26684
rect 19220 26630 19246 26682
rect 19246 26630 19276 26682
rect 19300 26630 19310 26682
rect 19310 26630 19356 26682
rect 19380 26630 19426 26682
rect 19426 26630 19436 26682
rect 19460 26630 19490 26682
rect 19490 26630 19516 26682
rect 19220 26628 19276 26630
rect 19300 26628 19356 26630
rect 19380 26628 19436 26630
rect 19460 26628 19516 26630
rect 19220 25594 19276 25596
rect 19300 25594 19356 25596
rect 19380 25594 19436 25596
rect 19460 25594 19516 25596
rect 19220 25542 19246 25594
rect 19246 25542 19276 25594
rect 19300 25542 19310 25594
rect 19310 25542 19356 25594
rect 19380 25542 19426 25594
rect 19426 25542 19436 25594
rect 19460 25542 19490 25594
rect 19490 25542 19516 25594
rect 19220 25540 19276 25542
rect 19300 25540 19356 25542
rect 19380 25540 19436 25542
rect 19460 25540 19516 25542
rect 19220 24506 19276 24508
rect 19300 24506 19356 24508
rect 19380 24506 19436 24508
rect 19460 24506 19516 24508
rect 19220 24454 19246 24506
rect 19246 24454 19276 24506
rect 19300 24454 19310 24506
rect 19310 24454 19356 24506
rect 19380 24454 19426 24506
rect 19426 24454 19436 24506
rect 19460 24454 19490 24506
rect 19490 24454 19516 24506
rect 19220 24452 19276 24454
rect 19300 24452 19356 24454
rect 19380 24452 19436 24454
rect 19460 24452 19516 24454
rect 19220 23418 19276 23420
rect 19300 23418 19356 23420
rect 19380 23418 19436 23420
rect 19460 23418 19516 23420
rect 19220 23366 19246 23418
rect 19246 23366 19276 23418
rect 19300 23366 19310 23418
rect 19310 23366 19356 23418
rect 19380 23366 19426 23418
rect 19426 23366 19436 23418
rect 19460 23366 19490 23418
rect 19490 23366 19516 23418
rect 19220 23364 19276 23366
rect 19300 23364 19356 23366
rect 19380 23364 19436 23366
rect 19460 23364 19516 23366
rect 19220 22330 19276 22332
rect 19300 22330 19356 22332
rect 19380 22330 19436 22332
rect 19460 22330 19516 22332
rect 19220 22278 19246 22330
rect 19246 22278 19276 22330
rect 19300 22278 19310 22330
rect 19310 22278 19356 22330
rect 19380 22278 19426 22330
rect 19426 22278 19436 22330
rect 19460 22278 19490 22330
rect 19490 22278 19516 22330
rect 19220 22276 19276 22278
rect 19300 22276 19356 22278
rect 19380 22276 19436 22278
rect 19460 22276 19516 22278
rect 14220 4378 14276 4380
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14220 4326 14246 4378
rect 14246 4326 14276 4378
rect 14300 4326 14310 4378
rect 14310 4326 14356 4378
rect 14380 4326 14426 4378
rect 14426 4326 14436 4378
rect 14460 4326 14490 4378
rect 14490 4326 14516 4378
rect 14220 4324 14276 4326
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 19220 21242 19276 21244
rect 19300 21242 19356 21244
rect 19380 21242 19436 21244
rect 19460 21242 19516 21244
rect 19220 21190 19246 21242
rect 19246 21190 19276 21242
rect 19300 21190 19310 21242
rect 19310 21190 19356 21242
rect 19380 21190 19426 21242
rect 19426 21190 19436 21242
rect 19460 21190 19490 21242
rect 19490 21190 19516 21242
rect 19220 21188 19276 21190
rect 19300 21188 19356 21190
rect 19380 21188 19436 21190
rect 19460 21188 19516 21190
rect 19220 20154 19276 20156
rect 19300 20154 19356 20156
rect 19380 20154 19436 20156
rect 19460 20154 19516 20156
rect 19220 20102 19246 20154
rect 19246 20102 19276 20154
rect 19300 20102 19310 20154
rect 19310 20102 19356 20154
rect 19380 20102 19426 20154
rect 19426 20102 19436 20154
rect 19460 20102 19490 20154
rect 19490 20102 19516 20154
rect 19220 20100 19276 20102
rect 19300 20100 19356 20102
rect 19380 20100 19436 20102
rect 19460 20100 19516 20102
rect 24220 39194 24276 39196
rect 24300 39194 24356 39196
rect 24380 39194 24436 39196
rect 24460 39194 24516 39196
rect 24220 39142 24246 39194
rect 24246 39142 24276 39194
rect 24300 39142 24310 39194
rect 24310 39142 24356 39194
rect 24380 39142 24426 39194
rect 24426 39142 24436 39194
rect 24460 39142 24490 39194
rect 24490 39142 24516 39194
rect 24220 39140 24276 39142
rect 24300 39140 24356 39142
rect 24380 39140 24436 39142
rect 24460 39140 24516 39142
rect 22842 15578 22898 15634
rect 22842 15498 22898 15554
rect 22840 13088 23216 13224
rect 22841 13068 23216 13088
rect 22841 12932 23217 13068
rect 22842 12846 23218 12902
rect 22843 12826 23218 12846
rect 22843 12690 23219 12826
rect 21822 6976 21878 7032
rect 21822 6296 21878 6352
rect 21730 6160 21786 6216
rect 24220 38106 24276 38108
rect 24300 38106 24356 38108
rect 24380 38106 24436 38108
rect 24460 38106 24516 38108
rect 24220 38054 24246 38106
rect 24246 38054 24276 38106
rect 24300 38054 24310 38106
rect 24310 38054 24356 38106
rect 24380 38054 24426 38106
rect 24426 38054 24436 38106
rect 24460 38054 24490 38106
rect 24490 38054 24516 38106
rect 24220 38052 24276 38054
rect 24300 38052 24356 38054
rect 24380 38052 24436 38054
rect 24460 38052 24516 38054
rect 24220 37018 24276 37020
rect 24300 37018 24356 37020
rect 24380 37018 24436 37020
rect 24460 37018 24516 37020
rect 24220 36966 24246 37018
rect 24246 36966 24276 37018
rect 24300 36966 24310 37018
rect 24310 36966 24356 37018
rect 24380 36966 24426 37018
rect 24426 36966 24436 37018
rect 24460 36966 24490 37018
rect 24490 36966 24516 37018
rect 24220 36964 24276 36966
rect 24300 36964 24356 36966
rect 24380 36964 24436 36966
rect 24460 36964 24516 36966
rect 24220 35930 24276 35932
rect 24300 35930 24356 35932
rect 24380 35930 24436 35932
rect 24460 35930 24516 35932
rect 24220 35878 24246 35930
rect 24246 35878 24276 35930
rect 24300 35878 24310 35930
rect 24310 35878 24356 35930
rect 24380 35878 24426 35930
rect 24426 35878 24436 35930
rect 24460 35878 24490 35930
rect 24490 35878 24516 35930
rect 24220 35876 24276 35878
rect 24300 35876 24356 35878
rect 24380 35876 24436 35878
rect 24460 35876 24516 35878
rect 24220 34842 24276 34844
rect 24300 34842 24356 34844
rect 24380 34842 24436 34844
rect 24460 34842 24516 34844
rect 24220 34790 24246 34842
rect 24246 34790 24276 34842
rect 24300 34790 24310 34842
rect 24310 34790 24356 34842
rect 24380 34790 24426 34842
rect 24426 34790 24436 34842
rect 24460 34790 24490 34842
rect 24490 34790 24516 34842
rect 24220 34788 24276 34790
rect 24300 34788 24356 34790
rect 24380 34788 24436 34790
rect 24460 34788 24516 34790
rect 24220 33754 24276 33756
rect 24300 33754 24356 33756
rect 24380 33754 24436 33756
rect 24460 33754 24516 33756
rect 24220 33702 24246 33754
rect 24246 33702 24276 33754
rect 24300 33702 24310 33754
rect 24310 33702 24356 33754
rect 24380 33702 24426 33754
rect 24426 33702 24436 33754
rect 24460 33702 24490 33754
rect 24490 33702 24516 33754
rect 24220 33700 24276 33702
rect 24300 33700 24356 33702
rect 24380 33700 24436 33702
rect 24460 33700 24516 33702
rect 24220 32666 24276 32668
rect 24300 32666 24356 32668
rect 24380 32666 24436 32668
rect 24460 32666 24516 32668
rect 24220 32614 24246 32666
rect 24246 32614 24276 32666
rect 24300 32614 24310 32666
rect 24310 32614 24356 32666
rect 24380 32614 24426 32666
rect 24426 32614 24436 32666
rect 24460 32614 24490 32666
rect 24490 32614 24516 32666
rect 24220 32612 24276 32614
rect 24300 32612 24356 32614
rect 24380 32612 24436 32614
rect 24460 32612 24516 32614
rect 24220 31578 24276 31580
rect 24300 31578 24356 31580
rect 24380 31578 24436 31580
rect 24460 31578 24516 31580
rect 24220 31526 24246 31578
rect 24246 31526 24276 31578
rect 24300 31526 24310 31578
rect 24310 31526 24356 31578
rect 24380 31526 24426 31578
rect 24426 31526 24436 31578
rect 24460 31526 24490 31578
rect 24490 31526 24516 31578
rect 24220 31524 24276 31526
rect 24300 31524 24356 31526
rect 24380 31524 24436 31526
rect 24460 31524 24516 31526
rect 24220 30490 24276 30492
rect 24300 30490 24356 30492
rect 24380 30490 24436 30492
rect 24460 30490 24516 30492
rect 24220 30438 24246 30490
rect 24246 30438 24276 30490
rect 24300 30438 24310 30490
rect 24310 30438 24356 30490
rect 24380 30438 24426 30490
rect 24426 30438 24436 30490
rect 24460 30438 24490 30490
rect 24490 30438 24516 30490
rect 24220 30436 24276 30438
rect 24300 30436 24356 30438
rect 24380 30436 24436 30438
rect 24460 30436 24516 30438
rect 24220 29402 24276 29404
rect 24300 29402 24356 29404
rect 24380 29402 24436 29404
rect 24460 29402 24516 29404
rect 24220 29350 24246 29402
rect 24246 29350 24276 29402
rect 24300 29350 24310 29402
rect 24310 29350 24356 29402
rect 24380 29350 24426 29402
rect 24426 29350 24436 29402
rect 24460 29350 24490 29402
rect 24490 29350 24516 29402
rect 24220 29348 24276 29350
rect 24300 29348 24356 29350
rect 24380 29348 24436 29350
rect 24460 29348 24516 29350
rect 24220 28314 24276 28316
rect 24300 28314 24356 28316
rect 24380 28314 24436 28316
rect 24460 28314 24516 28316
rect 24220 28262 24246 28314
rect 24246 28262 24276 28314
rect 24300 28262 24310 28314
rect 24310 28262 24356 28314
rect 24380 28262 24426 28314
rect 24426 28262 24436 28314
rect 24460 28262 24490 28314
rect 24490 28262 24516 28314
rect 24220 28260 24276 28262
rect 24300 28260 24356 28262
rect 24380 28260 24436 28262
rect 24460 28260 24516 28262
rect 24220 27226 24276 27228
rect 24300 27226 24356 27228
rect 24380 27226 24436 27228
rect 24460 27226 24516 27228
rect 24220 27174 24246 27226
rect 24246 27174 24276 27226
rect 24300 27174 24310 27226
rect 24310 27174 24356 27226
rect 24380 27174 24426 27226
rect 24426 27174 24436 27226
rect 24460 27174 24490 27226
rect 24490 27174 24516 27226
rect 24220 27172 24276 27174
rect 24300 27172 24356 27174
rect 24380 27172 24436 27174
rect 24460 27172 24516 27174
rect 24220 26138 24276 26140
rect 24300 26138 24356 26140
rect 24380 26138 24436 26140
rect 24460 26138 24516 26140
rect 24220 26086 24246 26138
rect 24246 26086 24276 26138
rect 24300 26086 24310 26138
rect 24310 26086 24356 26138
rect 24380 26086 24426 26138
rect 24426 26086 24436 26138
rect 24460 26086 24490 26138
rect 24490 26086 24516 26138
rect 24220 26084 24276 26086
rect 24300 26084 24356 26086
rect 24380 26084 24436 26086
rect 24460 26084 24516 26086
rect 24220 25050 24276 25052
rect 24300 25050 24356 25052
rect 24380 25050 24436 25052
rect 24460 25050 24516 25052
rect 24220 24998 24246 25050
rect 24246 24998 24276 25050
rect 24300 24998 24310 25050
rect 24310 24998 24356 25050
rect 24380 24998 24426 25050
rect 24426 24998 24436 25050
rect 24460 24998 24490 25050
rect 24490 24998 24516 25050
rect 24220 24996 24276 24998
rect 24300 24996 24356 24998
rect 24380 24996 24436 24998
rect 24460 24996 24516 24998
rect 24220 23962 24276 23964
rect 24300 23962 24356 23964
rect 24380 23962 24436 23964
rect 24460 23962 24516 23964
rect 24220 23910 24246 23962
rect 24246 23910 24276 23962
rect 24300 23910 24310 23962
rect 24310 23910 24356 23962
rect 24380 23910 24426 23962
rect 24426 23910 24436 23962
rect 24460 23910 24490 23962
rect 24490 23910 24516 23962
rect 24220 23908 24276 23910
rect 24300 23908 24356 23910
rect 24380 23908 24436 23910
rect 24460 23908 24516 23910
rect 24220 22874 24276 22876
rect 24300 22874 24356 22876
rect 24380 22874 24436 22876
rect 24460 22874 24516 22876
rect 24220 22822 24246 22874
rect 24246 22822 24276 22874
rect 24300 22822 24310 22874
rect 24310 22822 24356 22874
rect 24380 22822 24426 22874
rect 24426 22822 24436 22874
rect 24460 22822 24490 22874
rect 24490 22822 24516 22874
rect 24220 22820 24276 22822
rect 24300 22820 24356 22822
rect 24380 22820 24436 22822
rect 24460 22820 24516 22822
rect 24220 21786 24276 21788
rect 24300 21786 24356 21788
rect 24380 21786 24436 21788
rect 24460 21786 24516 21788
rect 24220 21734 24246 21786
rect 24246 21734 24276 21786
rect 24300 21734 24310 21786
rect 24310 21734 24356 21786
rect 24380 21734 24426 21786
rect 24426 21734 24436 21786
rect 24460 21734 24490 21786
rect 24490 21734 24516 21786
rect 24220 21732 24276 21734
rect 24300 21732 24356 21734
rect 24380 21732 24436 21734
rect 24460 21732 24516 21734
rect 24220 20698 24276 20700
rect 24300 20698 24356 20700
rect 24380 20698 24436 20700
rect 24460 20698 24516 20700
rect 24220 20646 24246 20698
rect 24246 20646 24276 20698
rect 24300 20646 24310 20698
rect 24310 20646 24356 20698
rect 24380 20646 24426 20698
rect 24426 20646 24436 20698
rect 24460 20646 24490 20698
rect 24490 20646 24516 20698
rect 24220 20644 24276 20646
rect 24300 20644 24356 20646
rect 24380 20644 24436 20646
rect 24460 20644 24516 20646
rect 24220 19610 24276 19612
rect 24300 19610 24356 19612
rect 24380 19610 24436 19612
rect 24460 19610 24516 19612
rect 24220 19558 24246 19610
rect 24246 19558 24276 19610
rect 24300 19558 24310 19610
rect 24310 19558 24356 19610
rect 24380 19558 24426 19610
rect 24426 19558 24436 19610
rect 24460 19558 24490 19610
rect 24490 19558 24516 19610
rect 24220 19556 24276 19558
rect 24300 19556 24356 19558
rect 24380 19556 24436 19558
rect 24460 19556 24516 19558
rect 29220 45178 29276 45180
rect 29300 45178 29356 45180
rect 29380 45178 29436 45180
rect 29460 45178 29516 45180
rect 29220 45126 29246 45178
rect 29246 45126 29276 45178
rect 29300 45126 29310 45178
rect 29310 45126 29356 45178
rect 29380 45126 29426 45178
rect 29426 45126 29436 45178
rect 29460 45126 29490 45178
rect 29490 45126 29516 45178
rect 29220 45124 29276 45126
rect 29300 45124 29356 45126
rect 29380 45124 29436 45126
rect 29460 45124 29516 45126
rect 39220 45178 39276 45180
rect 39300 45178 39356 45180
rect 39380 45178 39436 45180
rect 39460 45178 39516 45180
rect 39220 45126 39246 45178
rect 39246 45126 39276 45178
rect 39300 45126 39310 45178
rect 39310 45126 39356 45178
rect 39380 45126 39426 45178
rect 39426 45126 39436 45178
rect 39460 45126 39490 45178
rect 39490 45126 39516 45178
rect 39220 45124 39276 45126
rect 39300 45124 39356 45126
rect 39380 45124 39436 45126
rect 39460 45124 39516 45126
rect 34220 44634 34276 44636
rect 34300 44634 34356 44636
rect 34380 44634 34436 44636
rect 34460 44634 34516 44636
rect 34220 44582 34246 44634
rect 34246 44582 34276 44634
rect 34300 44582 34310 44634
rect 34310 44582 34356 44634
rect 34380 44582 34426 44634
rect 34426 44582 34436 44634
rect 34460 44582 34490 44634
rect 34490 44582 34516 44634
rect 34220 44580 34276 44582
rect 34300 44580 34356 44582
rect 34380 44580 34436 44582
rect 34460 44580 34516 44582
rect 44220 44634 44276 44636
rect 44300 44634 44356 44636
rect 44380 44634 44436 44636
rect 44460 44634 44516 44636
rect 44220 44582 44246 44634
rect 44246 44582 44276 44634
rect 44300 44582 44310 44634
rect 44310 44582 44356 44634
rect 44380 44582 44426 44634
rect 44426 44582 44436 44634
rect 44460 44582 44490 44634
rect 44490 44582 44516 44634
rect 44220 44580 44276 44582
rect 44300 44580 44356 44582
rect 44380 44580 44436 44582
rect 44460 44580 44516 44582
rect 29220 44090 29276 44092
rect 29300 44090 29356 44092
rect 29380 44090 29436 44092
rect 29460 44090 29516 44092
rect 29220 44038 29246 44090
rect 29246 44038 29276 44090
rect 29300 44038 29310 44090
rect 29310 44038 29356 44090
rect 29380 44038 29426 44090
rect 29426 44038 29436 44090
rect 29460 44038 29490 44090
rect 29490 44038 29516 44090
rect 29220 44036 29276 44038
rect 29300 44036 29356 44038
rect 29380 44036 29436 44038
rect 29460 44036 29516 44038
rect 39220 44090 39276 44092
rect 39300 44090 39356 44092
rect 39380 44090 39436 44092
rect 39460 44090 39516 44092
rect 39220 44038 39246 44090
rect 39246 44038 39276 44090
rect 39300 44038 39310 44090
rect 39310 44038 39356 44090
rect 39380 44038 39426 44090
rect 39426 44038 39436 44090
rect 39460 44038 39490 44090
rect 39490 44038 39516 44090
rect 39220 44036 39276 44038
rect 39300 44036 39356 44038
rect 39380 44036 39436 44038
rect 39460 44036 39516 44038
rect 34220 43546 34276 43548
rect 34300 43546 34356 43548
rect 34380 43546 34436 43548
rect 34460 43546 34516 43548
rect 34220 43494 34246 43546
rect 34246 43494 34276 43546
rect 34300 43494 34310 43546
rect 34310 43494 34356 43546
rect 34380 43494 34426 43546
rect 34426 43494 34436 43546
rect 34460 43494 34490 43546
rect 34490 43494 34516 43546
rect 34220 43492 34276 43494
rect 34300 43492 34356 43494
rect 34380 43492 34436 43494
rect 34460 43492 34516 43494
rect 44220 43546 44276 43548
rect 44300 43546 44356 43548
rect 44380 43546 44436 43548
rect 44460 43546 44516 43548
rect 44220 43494 44246 43546
rect 44246 43494 44276 43546
rect 44300 43494 44310 43546
rect 44310 43494 44356 43546
rect 44380 43494 44426 43546
rect 44426 43494 44436 43546
rect 44460 43494 44490 43546
rect 44490 43494 44516 43546
rect 44220 43492 44276 43494
rect 44300 43492 44356 43494
rect 44380 43492 44436 43494
rect 44460 43492 44516 43494
rect 29220 43002 29276 43004
rect 29300 43002 29356 43004
rect 29380 43002 29436 43004
rect 29460 43002 29516 43004
rect 29220 42950 29246 43002
rect 29246 42950 29276 43002
rect 29300 42950 29310 43002
rect 29310 42950 29356 43002
rect 29380 42950 29426 43002
rect 29426 42950 29436 43002
rect 29460 42950 29490 43002
rect 29490 42950 29516 43002
rect 29220 42948 29276 42950
rect 29300 42948 29356 42950
rect 29380 42948 29436 42950
rect 29460 42948 29516 42950
rect 39220 43002 39276 43004
rect 39300 43002 39356 43004
rect 39380 43002 39436 43004
rect 39460 43002 39516 43004
rect 39220 42950 39246 43002
rect 39246 42950 39276 43002
rect 39300 42950 39310 43002
rect 39310 42950 39356 43002
rect 39380 42950 39426 43002
rect 39426 42950 39436 43002
rect 39460 42950 39490 43002
rect 39490 42950 39516 43002
rect 39220 42948 39276 42950
rect 39300 42948 39356 42950
rect 39380 42948 39436 42950
rect 39460 42948 39516 42950
rect 34220 42458 34276 42460
rect 34300 42458 34356 42460
rect 34380 42458 34436 42460
rect 34460 42458 34516 42460
rect 34220 42406 34246 42458
rect 34246 42406 34276 42458
rect 34300 42406 34310 42458
rect 34310 42406 34356 42458
rect 34380 42406 34426 42458
rect 34426 42406 34436 42458
rect 34460 42406 34490 42458
rect 34490 42406 34516 42458
rect 34220 42404 34276 42406
rect 34300 42404 34356 42406
rect 34380 42404 34436 42406
rect 34460 42404 34516 42406
rect 29220 41914 29276 41916
rect 29300 41914 29356 41916
rect 29380 41914 29436 41916
rect 29460 41914 29516 41916
rect 29220 41862 29246 41914
rect 29246 41862 29276 41914
rect 29300 41862 29310 41914
rect 29310 41862 29356 41914
rect 29380 41862 29426 41914
rect 29426 41862 29436 41914
rect 29460 41862 29490 41914
rect 29490 41862 29516 41914
rect 29220 41860 29276 41862
rect 29300 41860 29356 41862
rect 29380 41860 29436 41862
rect 29460 41860 29516 41862
rect 34220 41370 34276 41372
rect 34300 41370 34356 41372
rect 34380 41370 34436 41372
rect 34460 41370 34516 41372
rect 34220 41318 34246 41370
rect 34246 41318 34276 41370
rect 34300 41318 34310 41370
rect 34310 41318 34356 41370
rect 34380 41318 34426 41370
rect 34426 41318 34436 41370
rect 34460 41318 34490 41370
rect 34490 41318 34516 41370
rect 34220 41316 34276 41318
rect 34300 41316 34356 41318
rect 34380 41316 34436 41318
rect 34460 41316 34516 41318
rect 29220 40826 29276 40828
rect 29300 40826 29356 40828
rect 29380 40826 29436 40828
rect 29460 40826 29516 40828
rect 29220 40774 29246 40826
rect 29246 40774 29276 40826
rect 29300 40774 29310 40826
rect 29310 40774 29356 40826
rect 29380 40774 29426 40826
rect 29426 40774 29436 40826
rect 29460 40774 29490 40826
rect 29490 40774 29516 40826
rect 29220 40772 29276 40774
rect 29300 40772 29356 40774
rect 29380 40772 29436 40774
rect 29460 40772 29516 40774
rect 34220 40282 34276 40284
rect 34300 40282 34356 40284
rect 34380 40282 34436 40284
rect 34460 40282 34516 40284
rect 34220 40230 34246 40282
rect 34246 40230 34276 40282
rect 34300 40230 34310 40282
rect 34310 40230 34356 40282
rect 34380 40230 34426 40282
rect 34426 40230 34436 40282
rect 34460 40230 34490 40282
rect 34490 40230 34516 40282
rect 34220 40228 34276 40230
rect 34300 40228 34356 40230
rect 34380 40228 34436 40230
rect 34460 40228 34516 40230
rect 29220 39738 29276 39740
rect 29300 39738 29356 39740
rect 29380 39738 29436 39740
rect 29460 39738 29516 39740
rect 29220 39686 29246 39738
rect 29246 39686 29276 39738
rect 29300 39686 29310 39738
rect 29310 39686 29356 39738
rect 29380 39686 29426 39738
rect 29426 39686 29436 39738
rect 29460 39686 29490 39738
rect 29490 39686 29516 39738
rect 29220 39684 29276 39686
rect 29300 39684 29356 39686
rect 29380 39684 29436 39686
rect 29460 39684 29516 39686
rect 34220 39194 34276 39196
rect 34300 39194 34356 39196
rect 34380 39194 34436 39196
rect 34460 39194 34516 39196
rect 34220 39142 34246 39194
rect 34246 39142 34276 39194
rect 34300 39142 34310 39194
rect 34310 39142 34356 39194
rect 34380 39142 34426 39194
rect 34426 39142 34436 39194
rect 34460 39142 34490 39194
rect 34490 39142 34516 39194
rect 34220 39140 34276 39142
rect 34300 39140 34356 39142
rect 34380 39140 34436 39142
rect 34460 39140 34516 39142
rect 29220 38650 29276 38652
rect 29300 38650 29356 38652
rect 29380 38650 29436 38652
rect 29460 38650 29516 38652
rect 29220 38598 29246 38650
rect 29246 38598 29276 38650
rect 29300 38598 29310 38650
rect 29310 38598 29356 38650
rect 29380 38598 29426 38650
rect 29426 38598 29436 38650
rect 29460 38598 29490 38650
rect 29490 38598 29516 38650
rect 29220 38596 29276 38598
rect 29300 38596 29356 38598
rect 29380 38596 29436 38598
rect 29460 38596 29516 38598
rect 29220 37562 29276 37564
rect 29300 37562 29356 37564
rect 29380 37562 29436 37564
rect 29460 37562 29516 37564
rect 29220 37510 29246 37562
rect 29246 37510 29276 37562
rect 29300 37510 29310 37562
rect 29310 37510 29356 37562
rect 29380 37510 29426 37562
rect 29426 37510 29436 37562
rect 29460 37510 29490 37562
rect 29490 37510 29516 37562
rect 29220 37508 29276 37510
rect 29300 37508 29356 37510
rect 29380 37508 29436 37510
rect 29460 37508 29516 37510
rect 29220 36474 29276 36476
rect 29300 36474 29356 36476
rect 29380 36474 29436 36476
rect 29460 36474 29516 36476
rect 29220 36422 29246 36474
rect 29246 36422 29276 36474
rect 29300 36422 29310 36474
rect 29310 36422 29356 36474
rect 29380 36422 29426 36474
rect 29426 36422 29436 36474
rect 29460 36422 29490 36474
rect 29490 36422 29516 36474
rect 29220 36420 29276 36422
rect 29300 36420 29356 36422
rect 29380 36420 29436 36422
rect 29460 36420 29516 36422
rect 29220 35386 29276 35388
rect 29300 35386 29356 35388
rect 29380 35386 29436 35388
rect 29460 35386 29516 35388
rect 29220 35334 29246 35386
rect 29246 35334 29276 35386
rect 29300 35334 29310 35386
rect 29310 35334 29356 35386
rect 29380 35334 29426 35386
rect 29426 35334 29436 35386
rect 29460 35334 29490 35386
rect 29490 35334 29516 35386
rect 29220 35332 29276 35334
rect 29300 35332 29356 35334
rect 29380 35332 29436 35334
rect 29460 35332 29516 35334
rect 29220 34298 29276 34300
rect 29300 34298 29356 34300
rect 29380 34298 29436 34300
rect 29460 34298 29516 34300
rect 29220 34246 29246 34298
rect 29246 34246 29276 34298
rect 29300 34246 29310 34298
rect 29310 34246 29356 34298
rect 29380 34246 29426 34298
rect 29426 34246 29436 34298
rect 29460 34246 29490 34298
rect 29490 34246 29516 34298
rect 29220 34244 29276 34246
rect 29300 34244 29356 34246
rect 29380 34244 29436 34246
rect 29460 34244 29516 34246
rect 29220 33210 29276 33212
rect 29300 33210 29356 33212
rect 29380 33210 29436 33212
rect 29460 33210 29516 33212
rect 29220 33158 29246 33210
rect 29246 33158 29276 33210
rect 29300 33158 29310 33210
rect 29310 33158 29356 33210
rect 29380 33158 29426 33210
rect 29426 33158 29436 33210
rect 29460 33158 29490 33210
rect 29490 33158 29516 33210
rect 29220 33156 29276 33158
rect 29300 33156 29356 33158
rect 29380 33156 29436 33158
rect 29460 33156 29516 33158
rect 29220 32122 29276 32124
rect 29300 32122 29356 32124
rect 29380 32122 29436 32124
rect 29460 32122 29516 32124
rect 29220 32070 29246 32122
rect 29246 32070 29276 32122
rect 29300 32070 29310 32122
rect 29310 32070 29356 32122
rect 29380 32070 29426 32122
rect 29426 32070 29436 32122
rect 29460 32070 29490 32122
rect 29490 32070 29516 32122
rect 29220 32068 29276 32070
rect 29300 32068 29356 32070
rect 29380 32068 29436 32070
rect 29460 32068 29516 32070
rect 29220 31034 29276 31036
rect 29300 31034 29356 31036
rect 29380 31034 29436 31036
rect 29460 31034 29516 31036
rect 29220 30982 29246 31034
rect 29246 30982 29276 31034
rect 29300 30982 29310 31034
rect 29310 30982 29356 31034
rect 29380 30982 29426 31034
rect 29426 30982 29436 31034
rect 29460 30982 29490 31034
rect 29490 30982 29516 31034
rect 29220 30980 29276 30982
rect 29300 30980 29356 30982
rect 29380 30980 29436 30982
rect 29460 30980 29516 30982
rect 29220 29946 29276 29948
rect 29300 29946 29356 29948
rect 29380 29946 29436 29948
rect 29460 29946 29516 29948
rect 29220 29894 29246 29946
rect 29246 29894 29276 29946
rect 29300 29894 29310 29946
rect 29310 29894 29356 29946
rect 29380 29894 29426 29946
rect 29426 29894 29436 29946
rect 29460 29894 29490 29946
rect 29490 29894 29516 29946
rect 29220 29892 29276 29894
rect 29300 29892 29356 29894
rect 29380 29892 29436 29894
rect 29460 29892 29516 29894
rect 29220 28858 29276 28860
rect 29300 28858 29356 28860
rect 29380 28858 29436 28860
rect 29460 28858 29516 28860
rect 29220 28806 29246 28858
rect 29246 28806 29276 28858
rect 29300 28806 29310 28858
rect 29310 28806 29356 28858
rect 29380 28806 29426 28858
rect 29426 28806 29436 28858
rect 29460 28806 29490 28858
rect 29490 28806 29516 28858
rect 29220 28804 29276 28806
rect 29300 28804 29356 28806
rect 29380 28804 29436 28806
rect 29460 28804 29516 28806
rect 29220 27770 29276 27772
rect 29300 27770 29356 27772
rect 29380 27770 29436 27772
rect 29460 27770 29516 27772
rect 29220 27718 29246 27770
rect 29246 27718 29276 27770
rect 29300 27718 29310 27770
rect 29310 27718 29356 27770
rect 29380 27718 29426 27770
rect 29426 27718 29436 27770
rect 29460 27718 29490 27770
rect 29490 27718 29516 27770
rect 29220 27716 29276 27718
rect 29300 27716 29356 27718
rect 29380 27716 29436 27718
rect 29460 27716 29516 27718
rect 29220 26682 29276 26684
rect 29300 26682 29356 26684
rect 29380 26682 29436 26684
rect 29460 26682 29516 26684
rect 29220 26630 29246 26682
rect 29246 26630 29276 26682
rect 29300 26630 29310 26682
rect 29310 26630 29356 26682
rect 29380 26630 29426 26682
rect 29426 26630 29436 26682
rect 29460 26630 29490 26682
rect 29490 26630 29516 26682
rect 29220 26628 29276 26630
rect 29300 26628 29356 26630
rect 29380 26628 29436 26630
rect 29460 26628 29516 26630
rect 29220 25594 29276 25596
rect 29300 25594 29356 25596
rect 29380 25594 29436 25596
rect 29460 25594 29516 25596
rect 29220 25542 29246 25594
rect 29246 25542 29276 25594
rect 29300 25542 29310 25594
rect 29310 25542 29356 25594
rect 29380 25542 29426 25594
rect 29426 25542 29436 25594
rect 29460 25542 29490 25594
rect 29490 25542 29516 25594
rect 29220 25540 29276 25542
rect 29300 25540 29356 25542
rect 29380 25540 29436 25542
rect 29460 25540 29516 25542
rect 29220 24506 29276 24508
rect 29300 24506 29356 24508
rect 29380 24506 29436 24508
rect 29460 24506 29516 24508
rect 29220 24454 29246 24506
rect 29246 24454 29276 24506
rect 29300 24454 29310 24506
rect 29310 24454 29356 24506
rect 29380 24454 29426 24506
rect 29426 24454 29436 24506
rect 29460 24454 29490 24506
rect 29490 24454 29516 24506
rect 29220 24452 29276 24454
rect 29300 24452 29356 24454
rect 29380 24452 29436 24454
rect 29460 24452 29516 24454
rect 29220 23418 29276 23420
rect 29300 23418 29356 23420
rect 29380 23418 29436 23420
rect 29460 23418 29516 23420
rect 29220 23366 29246 23418
rect 29246 23366 29276 23418
rect 29300 23366 29310 23418
rect 29310 23366 29356 23418
rect 29380 23366 29426 23418
rect 29426 23366 29436 23418
rect 29460 23366 29490 23418
rect 29490 23366 29516 23418
rect 29220 23364 29276 23366
rect 29300 23364 29356 23366
rect 29380 23364 29436 23366
rect 29460 23364 29516 23366
rect 29220 22330 29276 22332
rect 29300 22330 29356 22332
rect 29380 22330 29436 22332
rect 29460 22330 29516 22332
rect 29220 22278 29246 22330
rect 29246 22278 29276 22330
rect 29300 22278 29310 22330
rect 29310 22278 29356 22330
rect 29380 22278 29426 22330
rect 29426 22278 29436 22330
rect 29460 22278 29490 22330
rect 29490 22278 29516 22330
rect 29220 22276 29276 22278
rect 29300 22276 29356 22278
rect 29380 22276 29436 22278
rect 29460 22276 29516 22278
rect 29220 21242 29276 21244
rect 29300 21242 29356 21244
rect 29380 21242 29436 21244
rect 29460 21242 29516 21244
rect 29220 21190 29246 21242
rect 29246 21190 29276 21242
rect 29300 21190 29310 21242
rect 29310 21190 29356 21242
rect 29380 21190 29426 21242
rect 29426 21190 29436 21242
rect 29460 21190 29490 21242
rect 29490 21190 29516 21242
rect 29220 21188 29276 21190
rect 29300 21188 29356 21190
rect 29380 21188 29436 21190
rect 29460 21188 29516 21190
rect 29220 20154 29276 20156
rect 29300 20154 29356 20156
rect 29380 20154 29436 20156
rect 29460 20154 29516 20156
rect 29220 20102 29246 20154
rect 29246 20102 29276 20154
rect 29300 20102 29310 20154
rect 29310 20102 29356 20154
rect 29380 20102 29426 20154
rect 29426 20102 29436 20154
rect 29460 20102 29490 20154
rect 29490 20102 29516 20154
rect 29220 20100 29276 20102
rect 29300 20100 29356 20102
rect 29380 20100 29436 20102
rect 29460 20100 29516 20102
rect 34220 38106 34276 38108
rect 34300 38106 34356 38108
rect 34380 38106 34436 38108
rect 34460 38106 34516 38108
rect 34220 38054 34246 38106
rect 34246 38054 34276 38106
rect 34300 38054 34310 38106
rect 34310 38054 34356 38106
rect 34380 38054 34426 38106
rect 34426 38054 34436 38106
rect 34460 38054 34490 38106
rect 34490 38054 34516 38106
rect 34220 38052 34276 38054
rect 34300 38052 34356 38054
rect 34380 38052 34436 38054
rect 34460 38052 34516 38054
rect 34220 37018 34276 37020
rect 34300 37018 34356 37020
rect 34380 37018 34436 37020
rect 34460 37018 34516 37020
rect 34220 36966 34246 37018
rect 34246 36966 34276 37018
rect 34300 36966 34310 37018
rect 34310 36966 34356 37018
rect 34380 36966 34426 37018
rect 34426 36966 34436 37018
rect 34460 36966 34490 37018
rect 34490 36966 34516 37018
rect 34220 36964 34276 36966
rect 34300 36964 34356 36966
rect 34380 36964 34436 36966
rect 34460 36964 34516 36966
rect 34220 35930 34276 35932
rect 34300 35930 34356 35932
rect 34380 35930 34436 35932
rect 34460 35930 34516 35932
rect 34220 35878 34246 35930
rect 34246 35878 34276 35930
rect 34300 35878 34310 35930
rect 34310 35878 34356 35930
rect 34380 35878 34426 35930
rect 34426 35878 34436 35930
rect 34460 35878 34490 35930
rect 34490 35878 34516 35930
rect 34220 35876 34276 35878
rect 34300 35876 34356 35878
rect 34380 35876 34436 35878
rect 34460 35876 34516 35878
rect 34220 34842 34276 34844
rect 34300 34842 34356 34844
rect 34380 34842 34436 34844
rect 34460 34842 34516 34844
rect 34220 34790 34246 34842
rect 34246 34790 34276 34842
rect 34300 34790 34310 34842
rect 34310 34790 34356 34842
rect 34380 34790 34426 34842
rect 34426 34790 34436 34842
rect 34460 34790 34490 34842
rect 34490 34790 34516 34842
rect 34220 34788 34276 34790
rect 34300 34788 34356 34790
rect 34380 34788 34436 34790
rect 34460 34788 34516 34790
rect 34220 33754 34276 33756
rect 34300 33754 34356 33756
rect 34380 33754 34436 33756
rect 34460 33754 34516 33756
rect 34220 33702 34246 33754
rect 34246 33702 34276 33754
rect 34300 33702 34310 33754
rect 34310 33702 34356 33754
rect 34380 33702 34426 33754
rect 34426 33702 34436 33754
rect 34460 33702 34490 33754
rect 34490 33702 34516 33754
rect 34220 33700 34276 33702
rect 34300 33700 34356 33702
rect 34380 33700 34436 33702
rect 34460 33700 34516 33702
rect 34220 32666 34276 32668
rect 34300 32666 34356 32668
rect 34380 32666 34436 32668
rect 34460 32666 34516 32668
rect 34220 32614 34246 32666
rect 34246 32614 34276 32666
rect 34300 32614 34310 32666
rect 34310 32614 34356 32666
rect 34380 32614 34426 32666
rect 34426 32614 34436 32666
rect 34460 32614 34490 32666
rect 34490 32614 34516 32666
rect 34220 32612 34276 32614
rect 34300 32612 34356 32614
rect 34380 32612 34436 32614
rect 34460 32612 34516 32614
rect 34220 31578 34276 31580
rect 34300 31578 34356 31580
rect 34380 31578 34436 31580
rect 34460 31578 34516 31580
rect 34220 31526 34246 31578
rect 34246 31526 34276 31578
rect 34300 31526 34310 31578
rect 34310 31526 34356 31578
rect 34380 31526 34426 31578
rect 34426 31526 34436 31578
rect 34460 31526 34490 31578
rect 34490 31526 34516 31578
rect 34220 31524 34276 31526
rect 34300 31524 34356 31526
rect 34380 31524 34436 31526
rect 34460 31524 34516 31526
rect 34220 30490 34276 30492
rect 34300 30490 34356 30492
rect 34380 30490 34436 30492
rect 34460 30490 34516 30492
rect 34220 30438 34246 30490
rect 34246 30438 34276 30490
rect 34300 30438 34310 30490
rect 34310 30438 34356 30490
rect 34380 30438 34426 30490
rect 34426 30438 34436 30490
rect 34460 30438 34490 30490
rect 34490 30438 34516 30490
rect 34220 30436 34276 30438
rect 34300 30436 34356 30438
rect 34380 30436 34436 30438
rect 34460 30436 34516 30438
rect 39220 41914 39276 41916
rect 39300 41914 39356 41916
rect 39380 41914 39436 41916
rect 39460 41914 39516 41916
rect 39220 41862 39246 41914
rect 39246 41862 39276 41914
rect 39300 41862 39310 41914
rect 39310 41862 39356 41914
rect 39380 41862 39426 41914
rect 39426 41862 39436 41914
rect 39460 41862 39490 41914
rect 39490 41862 39516 41914
rect 39220 41860 39276 41862
rect 39300 41860 39356 41862
rect 39380 41860 39436 41862
rect 39460 41860 39516 41862
rect 39220 40826 39276 40828
rect 39300 40826 39356 40828
rect 39380 40826 39436 40828
rect 39460 40826 39516 40828
rect 39220 40774 39246 40826
rect 39246 40774 39276 40826
rect 39300 40774 39310 40826
rect 39310 40774 39356 40826
rect 39380 40774 39426 40826
rect 39426 40774 39436 40826
rect 39460 40774 39490 40826
rect 39490 40774 39516 40826
rect 39220 40772 39276 40774
rect 39300 40772 39356 40774
rect 39380 40772 39436 40774
rect 39460 40772 39516 40774
rect 39220 39738 39276 39740
rect 39300 39738 39356 39740
rect 39380 39738 39436 39740
rect 39460 39738 39516 39740
rect 39220 39686 39246 39738
rect 39246 39686 39276 39738
rect 39300 39686 39310 39738
rect 39310 39686 39356 39738
rect 39380 39686 39426 39738
rect 39426 39686 39436 39738
rect 39460 39686 39490 39738
rect 39490 39686 39516 39738
rect 39220 39684 39276 39686
rect 39300 39684 39356 39686
rect 39380 39684 39436 39686
rect 39460 39684 39516 39686
rect 39220 38650 39276 38652
rect 39300 38650 39356 38652
rect 39380 38650 39436 38652
rect 39460 38650 39516 38652
rect 39220 38598 39246 38650
rect 39246 38598 39276 38650
rect 39300 38598 39310 38650
rect 39310 38598 39356 38650
rect 39380 38598 39426 38650
rect 39426 38598 39436 38650
rect 39460 38598 39490 38650
rect 39490 38598 39516 38650
rect 39220 38596 39276 38598
rect 39300 38596 39356 38598
rect 39380 38596 39436 38598
rect 39460 38596 39516 38598
rect 34220 29402 34276 29404
rect 34300 29402 34356 29404
rect 34380 29402 34436 29404
rect 34460 29402 34516 29404
rect 34220 29350 34246 29402
rect 34246 29350 34276 29402
rect 34300 29350 34310 29402
rect 34310 29350 34356 29402
rect 34380 29350 34426 29402
rect 34426 29350 34436 29402
rect 34460 29350 34490 29402
rect 34490 29350 34516 29402
rect 34220 29348 34276 29350
rect 34300 29348 34356 29350
rect 34380 29348 34436 29350
rect 34460 29348 34516 29350
rect 34220 28314 34276 28316
rect 34300 28314 34356 28316
rect 34380 28314 34436 28316
rect 34460 28314 34516 28316
rect 34220 28262 34246 28314
rect 34246 28262 34276 28314
rect 34300 28262 34310 28314
rect 34310 28262 34356 28314
rect 34380 28262 34426 28314
rect 34426 28262 34436 28314
rect 34460 28262 34490 28314
rect 34490 28262 34516 28314
rect 34220 28260 34276 28262
rect 34300 28260 34356 28262
rect 34380 28260 34436 28262
rect 34460 28260 34516 28262
rect 34220 27226 34276 27228
rect 34300 27226 34356 27228
rect 34380 27226 34436 27228
rect 34460 27226 34516 27228
rect 34220 27174 34246 27226
rect 34246 27174 34276 27226
rect 34300 27174 34310 27226
rect 34310 27174 34356 27226
rect 34380 27174 34426 27226
rect 34426 27174 34436 27226
rect 34460 27174 34490 27226
rect 34490 27174 34516 27226
rect 34220 27172 34276 27174
rect 34300 27172 34356 27174
rect 34380 27172 34436 27174
rect 34460 27172 34516 27174
rect 34220 26138 34276 26140
rect 34300 26138 34356 26140
rect 34380 26138 34436 26140
rect 34460 26138 34516 26140
rect 34220 26086 34246 26138
rect 34246 26086 34276 26138
rect 34300 26086 34310 26138
rect 34310 26086 34356 26138
rect 34380 26086 34426 26138
rect 34426 26086 34436 26138
rect 34460 26086 34490 26138
rect 34490 26086 34516 26138
rect 34220 26084 34276 26086
rect 34300 26084 34356 26086
rect 34380 26084 34436 26086
rect 34460 26084 34516 26086
rect 34220 25050 34276 25052
rect 34300 25050 34356 25052
rect 34380 25050 34436 25052
rect 34460 25050 34516 25052
rect 34220 24998 34246 25050
rect 34246 24998 34276 25050
rect 34300 24998 34310 25050
rect 34310 24998 34356 25050
rect 34380 24998 34426 25050
rect 34426 24998 34436 25050
rect 34460 24998 34490 25050
rect 34490 24998 34516 25050
rect 34220 24996 34276 24998
rect 34300 24996 34356 24998
rect 34380 24996 34436 24998
rect 34460 24996 34516 24998
rect 34220 23962 34276 23964
rect 34300 23962 34356 23964
rect 34380 23962 34436 23964
rect 34460 23962 34516 23964
rect 34220 23910 34246 23962
rect 34246 23910 34276 23962
rect 34300 23910 34310 23962
rect 34310 23910 34356 23962
rect 34380 23910 34426 23962
rect 34426 23910 34436 23962
rect 34460 23910 34490 23962
rect 34490 23910 34516 23962
rect 34220 23908 34276 23910
rect 34300 23908 34356 23910
rect 34380 23908 34436 23910
rect 34460 23908 34516 23910
rect 34220 22874 34276 22876
rect 34300 22874 34356 22876
rect 34380 22874 34436 22876
rect 34460 22874 34516 22876
rect 34220 22822 34246 22874
rect 34246 22822 34276 22874
rect 34300 22822 34310 22874
rect 34310 22822 34356 22874
rect 34380 22822 34426 22874
rect 34426 22822 34436 22874
rect 34460 22822 34490 22874
rect 34490 22822 34516 22874
rect 34220 22820 34276 22822
rect 34300 22820 34356 22822
rect 34380 22820 34436 22822
rect 34460 22820 34516 22822
rect 34220 21786 34276 21788
rect 34300 21786 34356 21788
rect 34380 21786 34436 21788
rect 34460 21786 34516 21788
rect 34220 21734 34246 21786
rect 34246 21734 34276 21786
rect 34300 21734 34310 21786
rect 34310 21734 34356 21786
rect 34380 21734 34426 21786
rect 34426 21734 34436 21786
rect 34460 21734 34490 21786
rect 34490 21734 34516 21786
rect 34220 21732 34276 21734
rect 34300 21732 34356 21734
rect 34380 21732 34436 21734
rect 34460 21732 34516 21734
rect 34220 20698 34276 20700
rect 34300 20698 34356 20700
rect 34380 20698 34436 20700
rect 34460 20698 34516 20700
rect 34220 20646 34246 20698
rect 34246 20646 34276 20698
rect 34300 20646 34310 20698
rect 34310 20646 34356 20698
rect 34380 20646 34426 20698
rect 34426 20646 34436 20698
rect 34460 20646 34490 20698
rect 34490 20646 34516 20698
rect 34220 20644 34276 20646
rect 34300 20644 34356 20646
rect 34380 20644 34436 20646
rect 34460 20644 34516 20646
rect 34220 19610 34276 19612
rect 34300 19610 34356 19612
rect 34380 19610 34436 19612
rect 34460 19610 34516 19612
rect 34220 19558 34246 19610
rect 34246 19558 34276 19610
rect 34300 19558 34310 19610
rect 34310 19558 34356 19610
rect 34380 19558 34426 19610
rect 34426 19558 34436 19610
rect 34460 19558 34490 19610
rect 34490 19558 34516 19610
rect 34220 19556 34276 19558
rect 34300 19556 34356 19558
rect 34380 19556 34436 19558
rect 34460 19556 34516 19558
rect 24072 13083 24368 13219
rect 24950 6024 25006 6080
rect 32954 6024 33010 6080
rect 9220 2746 9276 2748
rect 9300 2746 9356 2748
rect 9380 2746 9436 2748
rect 9460 2746 9516 2748
rect 9220 2694 9246 2746
rect 9246 2694 9276 2746
rect 9300 2694 9310 2746
rect 9310 2694 9356 2746
rect 9380 2694 9426 2746
rect 9426 2694 9436 2746
rect 9460 2694 9490 2746
rect 9490 2694 9516 2746
rect 9220 2692 9276 2694
rect 9300 2692 9356 2694
rect 9380 2692 9436 2694
rect 9460 2692 9516 2694
rect 1398 2508 1454 2544
rect 1398 2488 1400 2508
rect 1400 2488 1452 2508
rect 1452 2488 1454 2508
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 14220 3290 14276 3292
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14220 3238 14246 3290
rect 14246 3238 14276 3290
rect 14300 3238 14310 3290
rect 14310 3238 14356 3290
rect 14380 3238 14426 3290
rect 14426 3238 14436 3290
rect 14460 3238 14490 3290
rect 14490 3238 14516 3290
rect 14220 3236 14276 3238
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 34610 6296 34666 6352
rect 37278 5888 37334 5944
rect 37922 11092 37924 11112
rect 37924 11092 37976 11112
rect 37976 11092 37978 11112
rect 37922 11056 37978 11092
rect 39220 37562 39276 37564
rect 39300 37562 39356 37564
rect 39380 37562 39436 37564
rect 39460 37562 39516 37564
rect 39220 37510 39246 37562
rect 39246 37510 39276 37562
rect 39300 37510 39310 37562
rect 39310 37510 39356 37562
rect 39380 37510 39426 37562
rect 39426 37510 39436 37562
rect 39460 37510 39490 37562
rect 39490 37510 39516 37562
rect 39220 37508 39276 37510
rect 39300 37508 39356 37510
rect 39380 37508 39436 37510
rect 39460 37508 39516 37510
rect 39220 36474 39276 36476
rect 39300 36474 39356 36476
rect 39380 36474 39436 36476
rect 39460 36474 39516 36476
rect 39220 36422 39246 36474
rect 39246 36422 39276 36474
rect 39300 36422 39310 36474
rect 39310 36422 39356 36474
rect 39380 36422 39426 36474
rect 39426 36422 39436 36474
rect 39460 36422 39490 36474
rect 39490 36422 39516 36474
rect 39220 36420 39276 36422
rect 39300 36420 39356 36422
rect 39380 36420 39436 36422
rect 39460 36420 39516 36422
rect 39220 35386 39276 35388
rect 39300 35386 39356 35388
rect 39380 35386 39436 35388
rect 39460 35386 39516 35388
rect 39220 35334 39246 35386
rect 39246 35334 39276 35386
rect 39300 35334 39310 35386
rect 39310 35334 39356 35386
rect 39380 35334 39426 35386
rect 39426 35334 39436 35386
rect 39460 35334 39490 35386
rect 39490 35334 39516 35386
rect 39220 35332 39276 35334
rect 39300 35332 39356 35334
rect 39380 35332 39436 35334
rect 39460 35332 39516 35334
rect 39220 34298 39276 34300
rect 39300 34298 39356 34300
rect 39380 34298 39436 34300
rect 39460 34298 39516 34300
rect 39220 34246 39246 34298
rect 39246 34246 39276 34298
rect 39300 34246 39310 34298
rect 39310 34246 39356 34298
rect 39380 34246 39426 34298
rect 39426 34246 39436 34298
rect 39460 34246 39490 34298
rect 39490 34246 39516 34298
rect 39220 34244 39276 34246
rect 39300 34244 39356 34246
rect 39380 34244 39436 34246
rect 39460 34244 39516 34246
rect 39220 33210 39276 33212
rect 39300 33210 39356 33212
rect 39380 33210 39436 33212
rect 39460 33210 39516 33212
rect 39220 33158 39246 33210
rect 39246 33158 39276 33210
rect 39300 33158 39310 33210
rect 39310 33158 39356 33210
rect 39380 33158 39426 33210
rect 39426 33158 39436 33210
rect 39460 33158 39490 33210
rect 39490 33158 39516 33210
rect 39220 33156 39276 33158
rect 39300 33156 39356 33158
rect 39380 33156 39436 33158
rect 39460 33156 39516 33158
rect 39220 32122 39276 32124
rect 39300 32122 39356 32124
rect 39380 32122 39436 32124
rect 39460 32122 39516 32124
rect 39220 32070 39246 32122
rect 39246 32070 39276 32122
rect 39300 32070 39310 32122
rect 39310 32070 39356 32122
rect 39380 32070 39426 32122
rect 39426 32070 39436 32122
rect 39460 32070 39490 32122
rect 39490 32070 39516 32122
rect 39220 32068 39276 32070
rect 39300 32068 39356 32070
rect 39380 32068 39436 32070
rect 39460 32068 39516 32070
rect 39220 31034 39276 31036
rect 39300 31034 39356 31036
rect 39380 31034 39436 31036
rect 39460 31034 39516 31036
rect 39220 30982 39246 31034
rect 39246 30982 39276 31034
rect 39300 30982 39310 31034
rect 39310 30982 39356 31034
rect 39380 30982 39426 31034
rect 39426 30982 39436 31034
rect 39460 30982 39490 31034
rect 39490 30982 39516 31034
rect 39220 30980 39276 30982
rect 39300 30980 39356 30982
rect 39380 30980 39436 30982
rect 39460 30980 39516 30982
rect 39220 29946 39276 29948
rect 39300 29946 39356 29948
rect 39380 29946 39436 29948
rect 39460 29946 39516 29948
rect 39220 29894 39246 29946
rect 39246 29894 39276 29946
rect 39300 29894 39310 29946
rect 39310 29894 39356 29946
rect 39380 29894 39426 29946
rect 39426 29894 39436 29946
rect 39460 29894 39490 29946
rect 39490 29894 39516 29946
rect 39220 29892 39276 29894
rect 39300 29892 39356 29894
rect 39380 29892 39436 29894
rect 39460 29892 39516 29894
rect 39220 28858 39276 28860
rect 39300 28858 39356 28860
rect 39380 28858 39436 28860
rect 39460 28858 39516 28860
rect 39220 28806 39246 28858
rect 39246 28806 39276 28858
rect 39300 28806 39310 28858
rect 39310 28806 39356 28858
rect 39380 28806 39426 28858
rect 39426 28806 39436 28858
rect 39460 28806 39490 28858
rect 39490 28806 39516 28858
rect 39220 28804 39276 28806
rect 39300 28804 39356 28806
rect 39380 28804 39436 28806
rect 39460 28804 39516 28806
rect 39220 27770 39276 27772
rect 39300 27770 39356 27772
rect 39380 27770 39436 27772
rect 39460 27770 39516 27772
rect 39220 27718 39246 27770
rect 39246 27718 39276 27770
rect 39300 27718 39310 27770
rect 39310 27718 39356 27770
rect 39380 27718 39426 27770
rect 39426 27718 39436 27770
rect 39460 27718 39490 27770
rect 39490 27718 39516 27770
rect 39220 27716 39276 27718
rect 39300 27716 39356 27718
rect 39380 27716 39436 27718
rect 39460 27716 39516 27718
rect 39220 26682 39276 26684
rect 39300 26682 39356 26684
rect 39380 26682 39436 26684
rect 39460 26682 39516 26684
rect 39220 26630 39246 26682
rect 39246 26630 39276 26682
rect 39300 26630 39310 26682
rect 39310 26630 39356 26682
rect 39380 26630 39426 26682
rect 39426 26630 39436 26682
rect 39460 26630 39490 26682
rect 39490 26630 39516 26682
rect 39220 26628 39276 26630
rect 39300 26628 39356 26630
rect 39380 26628 39436 26630
rect 39460 26628 39516 26630
rect 39220 25594 39276 25596
rect 39300 25594 39356 25596
rect 39380 25594 39436 25596
rect 39460 25594 39516 25596
rect 39220 25542 39246 25594
rect 39246 25542 39276 25594
rect 39300 25542 39310 25594
rect 39310 25542 39356 25594
rect 39380 25542 39426 25594
rect 39426 25542 39436 25594
rect 39460 25542 39490 25594
rect 39490 25542 39516 25594
rect 39220 25540 39276 25542
rect 39300 25540 39356 25542
rect 39380 25540 39436 25542
rect 39460 25540 39516 25542
rect 39220 24506 39276 24508
rect 39300 24506 39356 24508
rect 39380 24506 39436 24508
rect 39460 24506 39516 24508
rect 39220 24454 39246 24506
rect 39246 24454 39276 24506
rect 39300 24454 39310 24506
rect 39310 24454 39356 24506
rect 39380 24454 39426 24506
rect 39426 24454 39436 24506
rect 39460 24454 39490 24506
rect 39490 24454 39516 24506
rect 39220 24452 39276 24454
rect 39300 24452 39356 24454
rect 39380 24452 39436 24454
rect 39460 24452 39516 24454
rect 39220 23418 39276 23420
rect 39300 23418 39356 23420
rect 39380 23418 39436 23420
rect 39460 23418 39516 23420
rect 39220 23366 39246 23418
rect 39246 23366 39276 23418
rect 39300 23366 39310 23418
rect 39310 23366 39356 23418
rect 39380 23366 39426 23418
rect 39426 23366 39436 23418
rect 39460 23366 39490 23418
rect 39490 23366 39516 23418
rect 39220 23364 39276 23366
rect 39300 23364 39356 23366
rect 39380 23364 39436 23366
rect 39460 23364 39516 23366
rect 39220 22330 39276 22332
rect 39300 22330 39356 22332
rect 39380 22330 39436 22332
rect 39460 22330 39516 22332
rect 39220 22278 39246 22330
rect 39246 22278 39276 22330
rect 39300 22278 39310 22330
rect 39310 22278 39356 22330
rect 39380 22278 39426 22330
rect 39426 22278 39436 22330
rect 39460 22278 39490 22330
rect 39490 22278 39516 22330
rect 39220 22276 39276 22278
rect 39300 22276 39356 22278
rect 39380 22276 39436 22278
rect 39460 22276 39516 22278
rect 39220 21242 39276 21244
rect 39300 21242 39356 21244
rect 39380 21242 39436 21244
rect 39460 21242 39516 21244
rect 39220 21190 39246 21242
rect 39246 21190 39276 21242
rect 39300 21190 39310 21242
rect 39310 21190 39356 21242
rect 39380 21190 39426 21242
rect 39426 21190 39436 21242
rect 39460 21190 39490 21242
rect 39490 21190 39516 21242
rect 39220 21188 39276 21190
rect 39300 21188 39356 21190
rect 39380 21188 39436 21190
rect 39460 21188 39516 21190
rect 39220 20154 39276 20156
rect 39300 20154 39356 20156
rect 39380 20154 39436 20156
rect 39460 20154 39516 20156
rect 39220 20102 39246 20154
rect 39246 20102 39276 20154
rect 39300 20102 39310 20154
rect 39310 20102 39356 20154
rect 39380 20102 39426 20154
rect 39426 20102 39436 20154
rect 39460 20102 39490 20154
rect 39490 20102 39516 20154
rect 39220 20100 39276 20102
rect 39300 20100 39356 20102
rect 39380 20100 39436 20102
rect 39460 20100 39516 20102
rect 39220 19066 39276 19068
rect 39300 19066 39356 19068
rect 39380 19066 39436 19068
rect 39460 19066 39516 19068
rect 39220 19014 39246 19066
rect 39246 19014 39276 19066
rect 39300 19014 39310 19066
rect 39310 19014 39356 19066
rect 39380 19014 39426 19066
rect 39426 19014 39436 19066
rect 39460 19014 39490 19066
rect 39490 19014 39516 19066
rect 39220 19012 39276 19014
rect 39300 19012 39356 19014
rect 39380 19012 39436 19014
rect 39460 19012 39516 19014
rect 39220 17978 39276 17980
rect 39300 17978 39356 17980
rect 39380 17978 39436 17980
rect 39460 17978 39516 17980
rect 39220 17926 39246 17978
rect 39246 17926 39276 17978
rect 39300 17926 39310 17978
rect 39310 17926 39356 17978
rect 39380 17926 39426 17978
rect 39426 17926 39436 17978
rect 39460 17926 39490 17978
rect 39490 17926 39516 17978
rect 39220 17924 39276 17926
rect 39300 17924 39356 17926
rect 39380 17924 39436 17926
rect 39460 17924 39516 17926
rect 39220 16890 39276 16892
rect 39300 16890 39356 16892
rect 39380 16890 39436 16892
rect 39460 16890 39516 16892
rect 39220 16838 39246 16890
rect 39246 16838 39276 16890
rect 39300 16838 39310 16890
rect 39310 16838 39356 16890
rect 39380 16838 39426 16890
rect 39426 16838 39436 16890
rect 39460 16838 39490 16890
rect 39490 16838 39516 16890
rect 39220 16836 39276 16838
rect 39300 16836 39356 16838
rect 39380 16836 39436 16838
rect 39460 16836 39516 16838
rect 39220 15802 39276 15804
rect 39300 15802 39356 15804
rect 39380 15802 39436 15804
rect 39460 15802 39516 15804
rect 39220 15750 39246 15802
rect 39246 15750 39276 15802
rect 39300 15750 39310 15802
rect 39310 15750 39356 15802
rect 39380 15750 39426 15802
rect 39426 15750 39436 15802
rect 39460 15750 39490 15802
rect 39490 15750 39516 15802
rect 39220 15748 39276 15750
rect 39300 15748 39356 15750
rect 39380 15748 39436 15750
rect 39460 15748 39516 15750
rect 39220 14714 39276 14716
rect 39300 14714 39356 14716
rect 39380 14714 39436 14716
rect 39460 14714 39516 14716
rect 39220 14662 39246 14714
rect 39246 14662 39276 14714
rect 39300 14662 39310 14714
rect 39310 14662 39356 14714
rect 39380 14662 39426 14714
rect 39426 14662 39436 14714
rect 39460 14662 39490 14714
rect 39490 14662 39516 14714
rect 39220 14660 39276 14662
rect 39300 14660 39356 14662
rect 39380 14660 39436 14662
rect 39460 14660 39516 14662
rect 39220 13626 39276 13628
rect 39300 13626 39356 13628
rect 39380 13626 39436 13628
rect 39460 13626 39516 13628
rect 39220 13574 39246 13626
rect 39246 13574 39276 13626
rect 39300 13574 39310 13626
rect 39310 13574 39356 13626
rect 39380 13574 39426 13626
rect 39426 13574 39436 13626
rect 39460 13574 39490 13626
rect 39490 13574 39516 13626
rect 39220 13572 39276 13574
rect 39300 13572 39356 13574
rect 39380 13572 39436 13574
rect 39460 13572 39516 13574
rect 39220 12538 39276 12540
rect 39300 12538 39356 12540
rect 39380 12538 39436 12540
rect 39460 12538 39516 12540
rect 39220 12486 39246 12538
rect 39246 12486 39276 12538
rect 39300 12486 39310 12538
rect 39310 12486 39356 12538
rect 39380 12486 39426 12538
rect 39426 12486 39436 12538
rect 39460 12486 39490 12538
rect 39490 12486 39516 12538
rect 39220 12484 39276 12486
rect 39300 12484 39356 12486
rect 39380 12484 39436 12486
rect 39460 12484 39516 12486
rect 39220 11450 39276 11452
rect 39300 11450 39356 11452
rect 39380 11450 39436 11452
rect 39460 11450 39516 11452
rect 39220 11398 39246 11450
rect 39246 11398 39276 11450
rect 39300 11398 39310 11450
rect 39310 11398 39356 11450
rect 39380 11398 39426 11450
rect 39426 11398 39436 11450
rect 39460 11398 39490 11450
rect 39490 11398 39516 11450
rect 39220 11396 39276 11398
rect 39300 11396 39356 11398
rect 39380 11396 39436 11398
rect 39460 11396 39516 11398
rect 39220 10362 39276 10364
rect 39300 10362 39356 10364
rect 39380 10362 39436 10364
rect 39460 10362 39516 10364
rect 39220 10310 39246 10362
rect 39246 10310 39276 10362
rect 39300 10310 39310 10362
rect 39310 10310 39356 10362
rect 39380 10310 39426 10362
rect 39426 10310 39436 10362
rect 39460 10310 39490 10362
rect 39490 10310 39516 10362
rect 39220 10308 39276 10310
rect 39300 10308 39356 10310
rect 39380 10308 39436 10310
rect 39460 10308 39516 10310
rect 39220 9274 39276 9276
rect 39300 9274 39356 9276
rect 39380 9274 39436 9276
rect 39460 9274 39516 9276
rect 39220 9222 39246 9274
rect 39246 9222 39276 9274
rect 39300 9222 39310 9274
rect 39310 9222 39356 9274
rect 39380 9222 39426 9274
rect 39426 9222 39436 9274
rect 39460 9222 39490 9274
rect 39490 9222 39516 9274
rect 39220 9220 39276 9222
rect 39300 9220 39356 9222
rect 39380 9220 39436 9222
rect 39460 9220 39516 9222
rect 39220 8186 39276 8188
rect 39300 8186 39356 8188
rect 39380 8186 39436 8188
rect 39460 8186 39516 8188
rect 39220 8134 39246 8186
rect 39246 8134 39276 8186
rect 39300 8134 39310 8186
rect 39310 8134 39356 8186
rect 39380 8134 39426 8186
rect 39426 8134 39436 8186
rect 39460 8134 39490 8186
rect 39490 8134 39516 8186
rect 39220 8132 39276 8134
rect 39300 8132 39356 8134
rect 39380 8132 39436 8134
rect 39460 8132 39516 8134
rect 39220 7098 39276 7100
rect 39300 7098 39356 7100
rect 39380 7098 39436 7100
rect 39460 7098 39516 7100
rect 39220 7046 39246 7098
rect 39246 7046 39276 7098
rect 39300 7046 39310 7098
rect 39310 7046 39356 7098
rect 39380 7046 39426 7098
rect 39426 7046 39436 7098
rect 39460 7046 39490 7098
rect 39490 7046 39516 7098
rect 39220 7044 39276 7046
rect 39300 7044 39356 7046
rect 39380 7044 39436 7046
rect 39460 7044 39516 7046
rect 39220 6010 39276 6012
rect 39300 6010 39356 6012
rect 39380 6010 39436 6012
rect 39460 6010 39516 6012
rect 39220 5958 39246 6010
rect 39246 5958 39276 6010
rect 39300 5958 39310 6010
rect 39310 5958 39356 6010
rect 39380 5958 39426 6010
rect 39426 5958 39436 6010
rect 39460 5958 39490 6010
rect 39490 5958 39516 6010
rect 39220 5956 39276 5958
rect 39300 5956 39356 5958
rect 39380 5956 39436 5958
rect 39460 5956 39516 5958
rect 39220 4922 39276 4924
rect 39300 4922 39356 4924
rect 39380 4922 39436 4924
rect 39460 4922 39516 4924
rect 39220 4870 39246 4922
rect 39246 4870 39276 4922
rect 39300 4870 39310 4922
rect 39310 4870 39356 4922
rect 39380 4870 39426 4922
rect 39426 4870 39436 4922
rect 39460 4870 39490 4922
rect 39490 4870 39516 4922
rect 39220 4868 39276 4870
rect 39300 4868 39356 4870
rect 39380 4868 39436 4870
rect 39460 4868 39516 4870
rect 39220 3834 39276 3836
rect 39300 3834 39356 3836
rect 39380 3834 39436 3836
rect 39460 3834 39516 3836
rect 39220 3782 39246 3834
rect 39246 3782 39276 3834
rect 39300 3782 39310 3834
rect 39310 3782 39356 3834
rect 39380 3782 39426 3834
rect 39426 3782 39436 3834
rect 39460 3782 39490 3834
rect 39490 3782 39516 3834
rect 39220 3780 39276 3782
rect 39300 3780 39356 3782
rect 39380 3780 39436 3782
rect 39460 3780 39516 3782
rect 44220 42458 44276 42460
rect 44300 42458 44356 42460
rect 44380 42458 44436 42460
rect 44460 42458 44516 42460
rect 44220 42406 44246 42458
rect 44246 42406 44276 42458
rect 44300 42406 44310 42458
rect 44310 42406 44356 42458
rect 44380 42406 44426 42458
rect 44426 42406 44436 42458
rect 44460 42406 44490 42458
rect 44490 42406 44516 42458
rect 44220 42404 44276 42406
rect 44300 42404 44356 42406
rect 44380 42404 44436 42406
rect 44460 42404 44516 42406
rect 48134 41676 48190 41712
rect 48134 41656 48136 41676
rect 48136 41656 48188 41676
rect 48188 41656 48190 41676
rect 44220 41370 44276 41372
rect 44300 41370 44356 41372
rect 44380 41370 44436 41372
rect 44460 41370 44516 41372
rect 44220 41318 44246 41370
rect 44246 41318 44276 41370
rect 44300 41318 44310 41370
rect 44310 41318 44356 41370
rect 44380 41318 44426 41370
rect 44426 41318 44436 41370
rect 44460 41318 44490 41370
rect 44490 41318 44516 41370
rect 44220 41316 44276 41318
rect 44300 41316 44356 41318
rect 44380 41316 44436 41318
rect 44460 41316 44516 41318
rect 44220 40282 44276 40284
rect 44300 40282 44356 40284
rect 44380 40282 44436 40284
rect 44460 40282 44516 40284
rect 44220 40230 44246 40282
rect 44246 40230 44276 40282
rect 44300 40230 44310 40282
rect 44310 40230 44356 40282
rect 44380 40230 44426 40282
rect 44426 40230 44436 40282
rect 44460 40230 44490 40282
rect 44490 40230 44516 40282
rect 44220 40228 44276 40230
rect 44300 40228 44356 40230
rect 44380 40228 44436 40230
rect 44460 40228 44516 40230
rect 44220 39194 44276 39196
rect 44300 39194 44356 39196
rect 44380 39194 44436 39196
rect 44460 39194 44516 39196
rect 44220 39142 44246 39194
rect 44246 39142 44276 39194
rect 44300 39142 44310 39194
rect 44310 39142 44356 39194
rect 44380 39142 44426 39194
rect 44426 39142 44436 39194
rect 44460 39142 44490 39194
rect 44490 39142 44516 39194
rect 44220 39140 44276 39142
rect 44300 39140 44356 39142
rect 44380 39140 44436 39142
rect 44460 39140 44516 39142
rect 44220 38106 44276 38108
rect 44300 38106 44356 38108
rect 44380 38106 44436 38108
rect 44460 38106 44516 38108
rect 44220 38054 44246 38106
rect 44246 38054 44276 38106
rect 44300 38054 44310 38106
rect 44310 38054 44356 38106
rect 44380 38054 44426 38106
rect 44426 38054 44436 38106
rect 44460 38054 44490 38106
rect 44490 38054 44516 38106
rect 44220 38052 44276 38054
rect 44300 38052 44356 38054
rect 44380 38052 44436 38054
rect 44460 38052 44516 38054
rect 44220 37018 44276 37020
rect 44300 37018 44356 37020
rect 44380 37018 44436 37020
rect 44460 37018 44516 37020
rect 44220 36966 44246 37018
rect 44246 36966 44276 37018
rect 44300 36966 44310 37018
rect 44310 36966 44356 37018
rect 44380 36966 44426 37018
rect 44426 36966 44436 37018
rect 44460 36966 44490 37018
rect 44490 36966 44516 37018
rect 44220 36964 44276 36966
rect 44300 36964 44356 36966
rect 44380 36964 44436 36966
rect 44460 36964 44516 36966
rect 44220 35930 44276 35932
rect 44300 35930 44356 35932
rect 44380 35930 44436 35932
rect 44460 35930 44516 35932
rect 44220 35878 44246 35930
rect 44246 35878 44276 35930
rect 44300 35878 44310 35930
rect 44310 35878 44356 35930
rect 44380 35878 44426 35930
rect 44426 35878 44436 35930
rect 44460 35878 44490 35930
rect 44490 35878 44516 35930
rect 44220 35876 44276 35878
rect 44300 35876 44356 35878
rect 44380 35876 44436 35878
rect 44460 35876 44516 35878
rect 44220 34842 44276 34844
rect 44300 34842 44356 34844
rect 44380 34842 44436 34844
rect 44460 34842 44516 34844
rect 44220 34790 44246 34842
rect 44246 34790 44276 34842
rect 44300 34790 44310 34842
rect 44310 34790 44356 34842
rect 44380 34790 44426 34842
rect 44426 34790 44436 34842
rect 44460 34790 44490 34842
rect 44490 34790 44516 34842
rect 44220 34788 44276 34790
rect 44300 34788 44356 34790
rect 44380 34788 44436 34790
rect 44460 34788 44516 34790
rect 44220 33754 44276 33756
rect 44300 33754 44356 33756
rect 44380 33754 44436 33756
rect 44460 33754 44516 33756
rect 44220 33702 44246 33754
rect 44246 33702 44276 33754
rect 44300 33702 44310 33754
rect 44310 33702 44356 33754
rect 44380 33702 44426 33754
rect 44426 33702 44436 33754
rect 44460 33702 44490 33754
rect 44490 33702 44516 33754
rect 44220 33700 44276 33702
rect 44300 33700 44356 33702
rect 44380 33700 44436 33702
rect 44460 33700 44516 33702
rect 44220 32666 44276 32668
rect 44300 32666 44356 32668
rect 44380 32666 44436 32668
rect 44460 32666 44516 32668
rect 44220 32614 44246 32666
rect 44246 32614 44276 32666
rect 44300 32614 44310 32666
rect 44310 32614 44356 32666
rect 44380 32614 44426 32666
rect 44426 32614 44436 32666
rect 44460 32614 44490 32666
rect 44490 32614 44516 32666
rect 44220 32612 44276 32614
rect 44300 32612 44356 32614
rect 44380 32612 44436 32614
rect 44460 32612 44516 32614
rect 44220 31578 44276 31580
rect 44300 31578 44356 31580
rect 44380 31578 44436 31580
rect 44460 31578 44516 31580
rect 44220 31526 44246 31578
rect 44246 31526 44276 31578
rect 44300 31526 44310 31578
rect 44310 31526 44356 31578
rect 44380 31526 44426 31578
rect 44426 31526 44436 31578
rect 44460 31526 44490 31578
rect 44490 31526 44516 31578
rect 44220 31524 44276 31526
rect 44300 31524 44356 31526
rect 44380 31524 44436 31526
rect 44460 31524 44516 31526
rect 44220 30490 44276 30492
rect 44300 30490 44356 30492
rect 44380 30490 44436 30492
rect 44460 30490 44516 30492
rect 44220 30438 44246 30490
rect 44246 30438 44276 30490
rect 44300 30438 44310 30490
rect 44310 30438 44356 30490
rect 44380 30438 44426 30490
rect 44426 30438 44436 30490
rect 44460 30438 44490 30490
rect 44490 30438 44516 30490
rect 44220 30436 44276 30438
rect 44300 30436 44356 30438
rect 44380 30436 44436 30438
rect 44460 30436 44516 30438
rect 44220 29402 44276 29404
rect 44300 29402 44356 29404
rect 44380 29402 44436 29404
rect 44460 29402 44516 29404
rect 44220 29350 44246 29402
rect 44246 29350 44276 29402
rect 44300 29350 44310 29402
rect 44310 29350 44356 29402
rect 44380 29350 44426 29402
rect 44426 29350 44436 29402
rect 44460 29350 44490 29402
rect 44490 29350 44516 29402
rect 44220 29348 44276 29350
rect 44300 29348 44356 29350
rect 44380 29348 44436 29350
rect 44460 29348 44516 29350
rect 44220 28314 44276 28316
rect 44300 28314 44356 28316
rect 44380 28314 44436 28316
rect 44460 28314 44516 28316
rect 44220 28262 44246 28314
rect 44246 28262 44276 28314
rect 44300 28262 44310 28314
rect 44310 28262 44356 28314
rect 44380 28262 44426 28314
rect 44426 28262 44436 28314
rect 44460 28262 44490 28314
rect 44490 28262 44516 28314
rect 44220 28260 44276 28262
rect 44300 28260 44356 28262
rect 44380 28260 44436 28262
rect 44460 28260 44516 28262
rect 44220 27226 44276 27228
rect 44300 27226 44356 27228
rect 44380 27226 44436 27228
rect 44460 27226 44516 27228
rect 44220 27174 44246 27226
rect 44246 27174 44276 27226
rect 44300 27174 44310 27226
rect 44310 27174 44356 27226
rect 44380 27174 44426 27226
rect 44426 27174 44436 27226
rect 44460 27174 44490 27226
rect 44490 27174 44516 27226
rect 44220 27172 44276 27174
rect 44300 27172 44356 27174
rect 44380 27172 44436 27174
rect 44460 27172 44516 27174
rect 44220 26138 44276 26140
rect 44300 26138 44356 26140
rect 44380 26138 44436 26140
rect 44460 26138 44516 26140
rect 44220 26086 44246 26138
rect 44246 26086 44276 26138
rect 44300 26086 44310 26138
rect 44310 26086 44356 26138
rect 44380 26086 44426 26138
rect 44426 26086 44436 26138
rect 44460 26086 44490 26138
rect 44490 26086 44516 26138
rect 44220 26084 44276 26086
rect 44300 26084 44356 26086
rect 44380 26084 44436 26086
rect 44460 26084 44516 26086
rect 44220 25050 44276 25052
rect 44300 25050 44356 25052
rect 44380 25050 44436 25052
rect 44460 25050 44516 25052
rect 44220 24998 44246 25050
rect 44246 24998 44276 25050
rect 44300 24998 44310 25050
rect 44310 24998 44356 25050
rect 44380 24998 44426 25050
rect 44426 24998 44436 25050
rect 44460 24998 44490 25050
rect 44490 24998 44516 25050
rect 44220 24996 44276 24998
rect 44300 24996 44356 24998
rect 44380 24996 44436 24998
rect 44460 24996 44516 24998
rect 44220 23962 44276 23964
rect 44300 23962 44356 23964
rect 44380 23962 44436 23964
rect 44460 23962 44516 23964
rect 44220 23910 44246 23962
rect 44246 23910 44276 23962
rect 44300 23910 44310 23962
rect 44310 23910 44356 23962
rect 44380 23910 44426 23962
rect 44426 23910 44436 23962
rect 44460 23910 44490 23962
rect 44490 23910 44516 23962
rect 44220 23908 44276 23910
rect 44300 23908 44356 23910
rect 44380 23908 44436 23910
rect 44460 23908 44516 23910
rect 44220 22874 44276 22876
rect 44300 22874 44356 22876
rect 44380 22874 44436 22876
rect 44460 22874 44516 22876
rect 44220 22822 44246 22874
rect 44246 22822 44276 22874
rect 44300 22822 44310 22874
rect 44310 22822 44356 22874
rect 44380 22822 44426 22874
rect 44426 22822 44436 22874
rect 44460 22822 44490 22874
rect 44490 22822 44516 22874
rect 44220 22820 44276 22822
rect 44300 22820 44356 22822
rect 44380 22820 44436 22822
rect 44460 22820 44516 22822
rect 44220 21786 44276 21788
rect 44300 21786 44356 21788
rect 44380 21786 44436 21788
rect 44460 21786 44516 21788
rect 44220 21734 44246 21786
rect 44246 21734 44276 21786
rect 44300 21734 44310 21786
rect 44310 21734 44356 21786
rect 44380 21734 44426 21786
rect 44426 21734 44436 21786
rect 44460 21734 44490 21786
rect 44490 21734 44516 21786
rect 44220 21732 44276 21734
rect 44300 21732 44356 21734
rect 44380 21732 44436 21734
rect 44460 21732 44516 21734
rect 44220 20698 44276 20700
rect 44300 20698 44356 20700
rect 44380 20698 44436 20700
rect 44460 20698 44516 20700
rect 44220 20646 44246 20698
rect 44246 20646 44276 20698
rect 44300 20646 44310 20698
rect 44310 20646 44356 20698
rect 44380 20646 44426 20698
rect 44426 20646 44436 20698
rect 44460 20646 44490 20698
rect 44490 20646 44516 20698
rect 44220 20644 44276 20646
rect 44300 20644 44356 20646
rect 44380 20644 44436 20646
rect 44460 20644 44516 20646
rect 44220 19610 44276 19612
rect 44300 19610 44356 19612
rect 44380 19610 44436 19612
rect 44460 19610 44516 19612
rect 44220 19558 44246 19610
rect 44246 19558 44276 19610
rect 44300 19558 44310 19610
rect 44310 19558 44356 19610
rect 44380 19558 44426 19610
rect 44426 19558 44436 19610
rect 44460 19558 44490 19610
rect 44490 19558 44516 19610
rect 44220 19556 44276 19558
rect 44300 19556 44356 19558
rect 44380 19556 44436 19558
rect 44460 19556 44516 19558
rect 44220 18522 44276 18524
rect 44300 18522 44356 18524
rect 44380 18522 44436 18524
rect 44460 18522 44516 18524
rect 44220 18470 44246 18522
rect 44246 18470 44276 18522
rect 44300 18470 44310 18522
rect 44310 18470 44356 18522
rect 44380 18470 44426 18522
rect 44426 18470 44436 18522
rect 44460 18470 44490 18522
rect 44490 18470 44516 18522
rect 44220 18468 44276 18470
rect 44300 18468 44356 18470
rect 44380 18468 44436 18470
rect 44460 18468 44516 18470
rect 44220 17434 44276 17436
rect 44300 17434 44356 17436
rect 44380 17434 44436 17436
rect 44460 17434 44516 17436
rect 44220 17382 44246 17434
rect 44246 17382 44276 17434
rect 44300 17382 44310 17434
rect 44310 17382 44356 17434
rect 44380 17382 44426 17434
rect 44426 17382 44436 17434
rect 44460 17382 44490 17434
rect 44490 17382 44516 17434
rect 44220 17380 44276 17382
rect 44300 17380 44356 17382
rect 44380 17380 44436 17382
rect 44460 17380 44516 17382
rect 44220 16346 44276 16348
rect 44300 16346 44356 16348
rect 44380 16346 44436 16348
rect 44460 16346 44516 16348
rect 44220 16294 44246 16346
rect 44246 16294 44276 16346
rect 44300 16294 44310 16346
rect 44310 16294 44356 16346
rect 44380 16294 44426 16346
rect 44426 16294 44436 16346
rect 44460 16294 44490 16346
rect 44490 16294 44516 16346
rect 44220 16292 44276 16294
rect 44300 16292 44356 16294
rect 44380 16292 44436 16294
rect 44460 16292 44516 16294
rect 44220 15258 44276 15260
rect 44300 15258 44356 15260
rect 44380 15258 44436 15260
rect 44460 15258 44516 15260
rect 44220 15206 44246 15258
rect 44246 15206 44276 15258
rect 44300 15206 44310 15258
rect 44310 15206 44356 15258
rect 44380 15206 44426 15258
rect 44426 15206 44436 15258
rect 44460 15206 44490 15258
rect 44490 15206 44516 15258
rect 44220 15204 44276 15206
rect 44300 15204 44356 15206
rect 44380 15204 44436 15206
rect 44460 15204 44516 15206
rect 44220 14170 44276 14172
rect 44300 14170 44356 14172
rect 44380 14170 44436 14172
rect 44460 14170 44516 14172
rect 44220 14118 44246 14170
rect 44246 14118 44276 14170
rect 44300 14118 44310 14170
rect 44310 14118 44356 14170
rect 44380 14118 44426 14170
rect 44426 14118 44436 14170
rect 44460 14118 44490 14170
rect 44490 14118 44516 14170
rect 44220 14116 44276 14118
rect 44300 14116 44356 14118
rect 44380 14116 44436 14118
rect 44460 14116 44516 14118
rect 44220 13082 44276 13084
rect 44300 13082 44356 13084
rect 44380 13082 44436 13084
rect 44460 13082 44516 13084
rect 44220 13030 44246 13082
rect 44246 13030 44276 13082
rect 44300 13030 44310 13082
rect 44310 13030 44356 13082
rect 44380 13030 44426 13082
rect 44426 13030 44436 13082
rect 44460 13030 44490 13082
rect 44490 13030 44516 13082
rect 44220 13028 44276 13030
rect 44300 13028 44356 13030
rect 44380 13028 44436 13030
rect 44460 13028 44516 13030
rect 44220 11994 44276 11996
rect 44300 11994 44356 11996
rect 44380 11994 44436 11996
rect 44460 11994 44516 11996
rect 44220 11942 44246 11994
rect 44246 11942 44276 11994
rect 44300 11942 44310 11994
rect 44310 11942 44356 11994
rect 44380 11942 44426 11994
rect 44426 11942 44436 11994
rect 44460 11942 44490 11994
rect 44490 11942 44516 11994
rect 44220 11940 44276 11942
rect 44300 11940 44356 11942
rect 44380 11940 44436 11942
rect 44460 11940 44516 11942
rect 44220 10906 44276 10908
rect 44300 10906 44356 10908
rect 44380 10906 44436 10908
rect 44460 10906 44516 10908
rect 44220 10854 44246 10906
rect 44246 10854 44276 10906
rect 44300 10854 44310 10906
rect 44310 10854 44356 10906
rect 44380 10854 44426 10906
rect 44426 10854 44436 10906
rect 44460 10854 44490 10906
rect 44490 10854 44516 10906
rect 44220 10852 44276 10854
rect 44300 10852 44356 10854
rect 44380 10852 44436 10854
rect 44460 10852 44516 10854
rect 44220 9818 44276 9820
rect 44300 9818 44356 9820
rect 44380 9818 44436 9820
rect 44460 9818 44516 9820
rect 44220 9766 44246 9818
rect 44246 9766 44276 9818
rect 44300 9766 44310 9818
rect 44310 9766 44356 9818
rect 44380 9766 44426 9818
rect 44426 9766 44436 9818
rect 44460 9766 44490 9818
rect 44490 9766 44516 9818
rect 44220 9764 44276 9766
rect 44300 9764 44356 9766
rect 44380 9764 44436 9766
rect 44460 9764 44516 9766
rect 44220 8730 44276 8732
rect 44300 8730 44356 8732
rect 44380 8730 44436 8732
rect 44460 8730 44516 8732
rect 44220 8678 44246 8730
rect 44246 8678 44276 8730
rect 44300 8678 44310 8730
rect 44310 8678 44356 8730
rect 44380 8678 44426 8730
rect 44426 8678 44436 8730
rect 44460 8678 44490 8730
rect 44490 8678 44516 8730
rect 44220 8676 44276 8678
rect 44300 8676 44356 8678
rect 44380 8676 44436 8678
rect 44460 8676 44516 8678
rect 44220 7642 44276 7644
rect 44300 7642 44356 7644
rect 44380 7642 44436 7644
rect 44460 7642 44516 7644
rect 44220 7590 44246 7642
rect 44246 7590 44276 7642
rect 44300 7590 44310 7642
rect 44310 7590 44356 7642
rect 44380 7590 44426 7642
rect 44426 7590 44436 7642
rect 44460 7590 44490 7642
rect 44490 7590 44516 7642
rect 44220 7588 44276 7590
rect 44300 7588 44356 7590
rect 44380 7588 44436 7590
rect 44460 7588 44516 7590
rect 44220 6554 44276 6556
rect 44300 6554 44356 6556
rect 44380 6554 44436 6556
rect 44460 6554 44516 6556
rect 44220 6502 44246 6554
rect 44246 6502 44276 6554
rect 44300 6502 44310 6554
rect 44310 6502 44356 6554
rect 44380 6502 44426 6554
rect 44426 6502 44436 6554
rect 44460 6502 44490 6554
rect 44490 6502 44516 6554
rect 44220 6500 44276 6502
rect 44300 6500 44356 6502
rect 44380 6500 44436 6502
rect 44460 6500 44516 6502
rect 44220 5466 44276 5468
rect 44300 5466 44356 5468
rect 44380 5466 44436 5468
rect 44460 5466 44516 5468
rect 44220 5414 44246 5466
rect 44246 5414 44276 5466
rect 44300 5414 44310 5466
rect 44310 5414 44356 5466
rect 44380 5414 44426 5466
rect 44426 5414 44436 5466
rect 44460 5414 44490 5466
rect 44490 5414 44516 5466
rect 44220 5412 44276 5414
rect 44300 5412 44356 5414
rect 44380 5412 44436 5414
rect 44460 5412 44516 5414
rect 44220 4378 44276 4380
rect 44300 4378 44356 4380
rect 44380 4378 44436 4380
rect 44460 4378 44516 4380
rect 44220 4326 44246 4378
rect 44246 4326 44276 4378
rect 44300 4326 44310 4378
rect 44310 4326 44356 4378
rect 44380 4326 44426 4378
rect 44426 4326 44436 4378
rect 44460 4326 44490 4378
rect 44490 4326 44516 4378
rect 44220 4324 44276 4326
rect 44300 4324 44356 4326
rect 44380 4324 44436 4326
rect 44460 4324 44516 4326
rect 44220 3290 44276 3292
rect 44300 3290 44356 3292
rect 44380 3290 44436 3292
rect 44460 3290 44516 3292
rect 44220 3238 44246 3290
rect 44246 3238 44276 3290
rect 44300 3238 44310 3290
rect 44310 3238 44356 3290
rect 44380 3238 44426 3290
rect 44426 3238 44436 3290
rect 44460 3238 44490 3290
rect 44490 3238 44516 3290
rect 44220 3236 44276 3238
rect 44300 3236 44356 3238
rect 44380 3236 44436 3238
rect 44460 3236 44516 3238
rect 48134 24928 48190 24984
rect 48134 8336 48190 8392
rect 39220 2746 39276 2748
rect 39300 2746 39356 2748
rect 39380 2746 39436 2748
rect 39460 2746 39516 2748
rect 39220 2694 39246 2746
rect 39246 2694 39276 2746
rect 39300 2694 39310 2746
rect 39310 2694 39356 2746
rect 39380 2694 39426 2746
rect 39426 2694 39436 2746
rect 39460 2694 39490 2746
rect 39490 2694 39516 2746
rect 39220 2692 39276 2694
rect 39300 2692 39356 2694
rect 39380 2692 39436 2694
rect 39460 2692 39516 2694
rect 14220 2202 14276 2204
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14220 2150 14246 2202
rect 14246 2150 14276 2202
rect 14300 2150 14310 2202
rect 14310 2150 14356 2202
rect 14380 2150 14426 2202
rect 14426 2150 14436 2202
rect 14460 2150 14490 2202
rect 14490 2150 14516 2202
rect 14220 2148 14276 2150
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 44220 2202 44276 2204
rect 44300 2202 44356 2204
rect 44380 2202 44436 2204
rect 44460 2202 44516 2204
rect 44220 2150 44246 2202
rect 44246 2150 44276 2202
rect 44300 2150 44310 2202
rect 44310 2150 44356 2202
rect 44380 2150 44426 2202
rect 44426 2150 44436 2202
rect 44460 2150 44490 2202
rect 44490 2150 44516 2202
rect 44220 2148 44276 2150
rect 44300 2148 44356 2150
rect 44380 2148 44436 2150
rect 44460 2148 44516 2150
<< metal3 >>
rect 0 47562 800 47592
rect 1853 47562 1919 47565
rect 0 47560 1919 47562
rect 0 47504 1858 47560
rect 1914 47504 1919 47560
rect 0 47502 1919 47504
rect 0 47472 800 47502
rect 1853 47499 1919 47502
rect 9208 47360 9528 47361
rect 9208 47296 9216 47360
rect 9280 47296 9296 47360
rect 9360 47296 9376 47360
rect 9440 47296 9456 47360
rect 9520 47296 9528 47360
rect 9208 47295 9528 47296
rect 19208 47360 19528 47361
rect 19208 47296 19216 47360
rect 19280 47296 19296 47360
rect 19360 47296 19376 47360
rect 19440 47296 19456 47360
rect 19520 47296 19528 47360
rect 19208 47295 19528 47296
rect 29208 47360 29528 47361
rect 29208 47296 29216 47360
rect 29280 47296 29296 47360
rect 29360 47296 29376 47360
rect 29440 47296 29456 47360
rect 29520 47296 29528 47360
rect 29208 47295 29528 47296
rect 39208 47360 39528 47361
rect 39208 47296 39216 47360
rect 39280 47296 39296 47360
rect 39360 47296 39376 47360
rect 39440 47296 39456 47360
rect 39520 47296 39528 47360
rect 39208 47295 39528 47296
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 14208 46816 14528 46817
rect 14208 46752 14216 46816
rect 14280 46752 14296 46816
rect 14360 46752 14376 46816
rect 14440 46752 14456 46816
rect 14520 46752 14528 46816
rect 14208 46751 14528 46752
rect 24208 46816 24528 46817
rect 24208 46752 24216 46816
rect 24280 46752 24296 46816
rect 24360 46752 24376 46816
rect 24440 46752 24456 46816
rect 24520 46752 24528 46816
rect 24208 46751 24528 46752
rect 34208 46816 34528 46817
rect 34208 46752 34216 46816
rect 34280 46752 34296 46816
rect 34360 46752 34376 46816
rect 34440 46752 34456 46816
rect 34520 46752 34528 46816
rect 34208 46751 34528 46752
rect 44208 46816 44528 46817
rect 44208 46752 44216 46816
rect 44280 46752 44296 46816
rect 44360 46752 44376 46816
rect 44440 46752 44456 46816
rect 44520 46752 44528 46816
rect 44208 46751 44528 46752
rect 9208 46272 9528 46273
rect 9208 46208 9216 46272
rect 9280 46208 9296 46272
rect 9360 46208 9376 46272
rect 9440 46208 9456 46272
rect 9520 46208 9528 46272
rect 9208 46207 9528 46208
rect 19208 46272 19528 46273
rect 19208 46208 19216 46272
rect 19280 46208 19296 46272
rect 19360 46208 19376 46272
rect 19440 46208 19456 46272
rect 19520 46208 19528 46272
rect 19208 46207 19528 46208
rect 29208 46272 29528 46273
rect 29208 46208 29216 46272
rect 29280 46208 29296 46272
rect 29360 46208 29376 46272
rect 29440 46208 29456 46272
rect 29520 46208 29528 46272
rect 29208 46207 29528 46208
rect 39208 46272 39528 46273
rect 39208 46208 39216 46272
rect 39280 46208 39296 46272
rect 39360 46208 39376 46272
rect 39440 46208 39456 46272
rect 39520 46208 39528 46272
rect 39208 46207 39528 46208
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 14208 45728 14528 45729
rect 14208 45664 14216 45728
rect 14280 45664 14296 45728
rect 14360 45664 14376 45728
rect 14440 45664 14456 45728
rect 14520 45664 14528 45728
rect 14208 45663 14528 45664
rect 24208 45728 24528 45729
rect 24208 45664 24216 45728
rect 24280 45664 24296 45728
rect 24360 45664 24376 45728
rect 24440 45664 24456 45728
rect 24520 45664 24528 45728
rect 24208 45663 24528 45664
rect 34208 45728 34528 45729
rect 34208 45664 34216 45728
rect 34280 45664 34296 45728
rect 34360 45664 34376 45728
rect 34440 45664 34456 45728
rect 34520 45664 34528 45728
rect 34208 45663 34528 45664
rect 44208 45728 44528 45729
rect 44208 45664 44216 45728
rect 44280 45664 44296 45728
rect 44360 45664 44376 45728
rect 44440 45664 44456 45728
rect 44520 45664 44528 45728
rect 44208 45663 44528 45664
rect 9208 45184 9528 45185
rect 9208 45120 9216 45184
rect 9280 45120 9296 45184
rect 9360 45120 9376 45184
rect 9440 45120 9456 45184
rect 9520 45120 9528 45184
rect 9208 45119 9528 45120
rect 19208 45184 19528 45185
rect 19208 45120 19216 45184
rect 19280 45120 19296 45184
rect 19360 45120 19376 45184
rect 19440 45120 19456 45184
rect 19520 45120 19528 45184
rect 19208 45119 19528 45120
rect 29208 45184 29528 45185
rect 29208 45120 29216 45184
rect 29280 45120 29296 45184
rect 29360 45120 29376 45184
rect 29440 45120 29456 45184
rect 29520 45120 29528 45184
rect 29208 45119 29528 45120
rect 39208 45184 39528 45185
rect 39208 45120 39216 45184
rect 39280 45120 39296 45184
rect 39360 45120 39376 45184
rect 39440 45120 39456 45184
rect 39520 45120 39528 45184
rect 39208 45119 39528 45120
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 14208 44640 14528 44641
rect 14208 44576 14216 44640
rect 14280 44576 14296 44640
rect 14360 44576 14376 44640
rect 14440 44576 14456 44640
rect 14520 44576 14528 44640
rect 14208 44575 14528 44576
rect 24208 44640 24528 44641
rect 24208 44576 24216 44640
rect 24280 44576 24296 44640
rect 24360 44576 24376 44640
rect 24440 44576 24456 44640
rect 24520 44576 24528 44640
rect 24208 44575 24528 44576
rect 34208 44640 34528 44641
rect 34208 44576 34216 44640
rect 34280 44576 34296 44640
rect 34360 44576 34376 44640
rect 34440 44576 34456 44640
rect 34520 44576 34528 44640
rect 34208 44575 34528 44576
rect 44208 44640 44528 44641
rect 44208 44576 44216 44640
rect 44280 44576 44296 44640
rect 44360 44576 44376 44640
rect 44440 44576 44456 44640
rect 44520 44576 44528 44640
rect 44208 44575 44528 44576
rect 9208 44096 9528 44097
rect 9208 44032 9216 44096
rect 9280 44032 9296 44096
rect 9360 44032 9376 44096
rect 9440 44032 9456 44096
rect 9520 44032 9528 44096
rect 9208 44031 9528 44032
rect 19208 44096 19528 44097
rect 19208 44032 19216 44096
rect 19280 44032 19296 44096
rect 19360 44032 19376 44096
rect 19440 44032 19456 44096
rect 19520 44032 19528 44096
rect 19208 44031 19528 44032
rect 29208 44096 29528 44097
rect 29208 44032 29216 44096
rect 29280 44032 29296 44096
rect 29360 44032 29376 44096
rect 29440 44032 29456 44096
rect 29520 44032 29528 44096
rect 29208 44031 29528 44032
rect 39208 44096 39528 44097
rect 39208 44032 39216 44096
rect 39280 44032 39296 44096
rect 39360 44032 39376 44096
rect 39440 44032 39456 44096
rect 39520 44032 39528 44096
rect 39208 44031 39528 44032
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 14208 43552 14528 43553
rect 14208 43488 14216 43552
rect 14280 43488 14296 43552
rect 14360 43488 14376 43552
rect 14440 43488 14456 43552
rect 14520 43488 14528 43552
rect 14208 43487 14528 43488
rect 24208 43552 24528 43553
rect 24208 43488 24216 43552
rect 24280 43488 24296 43552
rect 24360 43488 24376 43552
rect 24440 43488 24456 43552
rect 24520 43488 24528 43552
rect 24208 43487 24528 43488
rect 34208 43552 34528 43553
rect 34208 43488 34216 43552
rect 34280 43488 34296 43552
rect 34360 43488 34376 43552
rect 34440 43488 34456 43552
rect 34520 43488 34528 43552
rect 34208 43487 34528 43488
rect 44208 43552 44528 43553
rect 44208 43488 44216 43552
rect 44280 43488 44296 43552
rect 44360 43488 44376 43552
rect 44440 43488 44456 43552
rect 44520 43488 44528 43552
rect 44208 43487 44528 43488
rect 9208 43008 9528 43009
rect 9208 42944 9216 43008
rect 9280 42944 9296 43008
rect 9360 42944 9376 43008
rect 9440 42944 9456 43008
rect 9520 42944 9528 43008
rect 9208 42943 9528 42944
rect 19208 43008 19528 43009
rect 19208 42944 19216 43008
rect 19280 42944 19296 43008
rect 19360 42944 19376 43008
rect 19440 42944 19456 43008
rect 19520 42944 19528 43008
rect 19208 42943 19528 42944
rect 29208 43008 29528 43009
rect 29208 42944 29216 43008
rect 29280 42944 29296 43008
rect 29360 42944 29376 43008
rect 29440 42944 29456 43008
rect 29520 42944 29528 43008
rect 29208 42943 29528 42944
rect 39208 43008 39528 43009
rect 39208 42944 39216 43008
rect 39280 42944 39296 43008
rect 39360 42944 39376 43008
rect 39440 42944 39456 43008
rect 39520 42944 39528 43008
rect 39208 42943 39528 42944
rect 0 42530 800 42560
rect 1853 42530 1919 42533
rect 0 42528 1919 42530
rect 0 42472 1858 42528
rect 1914 42472 1919 42528
rect 0 42470 1919 42472
rect 0 42440 800 42470
rect 1853 42467 1919 42470
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 14208 42464 14528 42465
rect 14208 42400 14216 42464
rect 14280 42400 14296 42464
rect 14360 42400 14376 42464
rect 14440 42400 14456 42464
rect 14520 42400 14528 42464
rect 14208 42399 14528 42400
rect 24208 42464 24528 42465
rect 24208 42400 24216 42464
rect 24280 42400 24296 42464
rect 24360 42400 24376 42464
rect 24440 42400 24456 42464
rect 24520 42400 24528 42464
rect 24208 42399 24528 42400
rect 34208 42464 34528 42465
rect 34208 42400 34216 42464
rect 34280 42400 34296 42464
rect 34360 42400 34376 42464
rect 34440 42400 34456 42464
rect 34520 42400 34528 42464
rect 34208 42399 34528 42400
rect 44208 42464 44528 42465
rect 44208 42400 44216 42464
rect 44280 42400 44296 42464
rect 44360 42400 44376 42464
rect 44440 42400 44456 42464
rect 44520 42400 44528 42464
rect 44208 42399 44528 42400
rect 9208 41920 9528 41921
rect 9208 41856 9216 41920
rect 9280 41856 9296 41920
rect 9360 41856 9376 41920
rect 9440 41856 9456 41920
rect 9520 41856 9528 41920
rect 9208 41855 9528 41856
rect 19208 41920 19528 41921
rect 19208 41856 19216 41920
rect 19280 41856 19296 41920
rect 19360 41856 19376 41920
rect 19440 41856 19456 41920
rect 19520 41856 19528 41920
rect 19208 41855 19528 41856
rect 29208 41920 29528 41921
rect 29208 41856 29216 41920
rect 29280 41856 29296 41920
rect 29360 41856 29376 41920
rect 29440 41856 29456 41920
rect 29520 41856 29528 41920
rect 29208 41855 29528 41856
rect 39208 41920 39528 41921
rect 39208 41856 39216 41920
rect 39280 41856 39296 41920
rect 39360 41856 39376 41920
rect 39440 41856 39456 41920
rect 39520 41856 39528 41920
rect 39208 41855 39528 41856
rect 48129 41714 48195 41717
rect 49200 41714 50000 41744
rect 48129 41712 50000 41714
rect 48129 41656 48134 41712
rect 48190 41656 50000 41712
rect 48129 41654 50000 41656
rect 48129 41651 48195 41654
rect 49200 41624 50000 41654
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 14208 41376 14528 41377
rect 14208 41312 14216 41376
rect 14280 41312 14296 41376
rect 14360 41312 14376 41376
rect 14440 41312 14456 41376
rect 14520 41312 14528 41376
rect 14208 41311 14528 41312
rect 24208 41376 24528 41377
rect 24208 41312 24216 41376
rect 24280 41312 24296 41376
rect 24360 41312 24376 41376
rect 24440 41312 24456 41376
rect 24520 41312 24528 41376
rect 24208 41311 24528 41312
rect 34208 41376 34528 41377
rect 34208 41312 34216 41376
rect 34280 41312 34296 41376
rect 34360 41312 34376 41376
rect 34440 41312 34456 41376
rect 34520 41312 34528 41376
rect 34208 41311 34528 41312
rect 44208 41376 44528 41377
rect 44208 41312 44216 41376
rect 44280 41312 44296 41376
rect 44360 41312 44376 41376
rect 44440 41312 44456 41376
rect 44520 41312 44528 41376
rect 44208 41311 44528 41312
rect 9208 40832 9528 40833
rect 9208 40768 9216 40832
rect 9280 40768 9296 40832
rect 9360 40768 9376 40832
rect 9440 40768 9456 40832
rect 9520 40768 9528 40832
rect 9208 40767 9528 40768
rect 19208 40832 19528 40833
rect 19208 40768 19216 40832
rect 19280 40768 19296 40832
rect 19360 40768 19376 40832
rect 19440 40768 19456 40832
rect 19520 40768 19528 40832
rect 19208 40767 19528 40768
rect 29208 40832 29528 40833
rect 29208 40768 29216 40832
rect 29280 40768 29296 40832
rect 29360 40768 29376 40832
rect 29440 40768 29456 40832
rect 29520 40768 29528 40832
rect 29208 40767 29528 40768
rect 39208 40832 39528 40833
rect 39208 40768 39216 40832
rect 39280 40768 39296 40832
rect 39360 40768 39376 40832
rect 39440 40768 39456 40832
rect 39520 40768 39528 40832
rect 39208 40767 39528 40768
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 14208 40288 14528 40289
rect 14208 40224 14216 40288
rect 14280 40224 14296 40288
rect 14360 40224 14376 40288
rect 14440 40224 14456 40288
rect 14520 40224 14528 40288
rect 14208 40223 14528 40224
rect 24208 40288 24528 40289
rect 24208 40224 24216 40288
rect 24280 40224 24296 40288
rect 24360 40224 24376 40288
rect 24440 40224 24456 40288
rect 24520 40224 24528 40288
rect 24208 40223 24528 40224
rect 34208 40288 34528 40289
rect 34208 40224 34216 40288
rect 34280 40224 34296 40288
rect 34360 40224 34376 40288
rect 34440 40224 34456 40288
rect 34520 40224 34528 40288
rect 34208 40223 34528 40224
rect 44208 40288 44528 40289
rect 44208 40224 44216 40288
rect 44280 40224 44296 40288
rect 44360 40224 44376 40288
rect 44440 40224 44456 40288
rect 44520 40224 44528 40288
rect 44208 40223 44528 40224
rect 9208 39744 9528 39745
rect 9208 39680 9216 39744
rect 9280 39680 9296 39744
rect 9360 39680 9376 39744
rect 9440 39680 9456 39744
rect 9520 39680 9528 39744
rect 9208 39679 9528 39680
rect 19208 39744 19528 39745
rect 19208 39680 19216 39744
rect 19280 39680 19296 39744
rect 19360 39680 19376 39744
rect 19440 39680 19456 39744
rect 19520 39680 19528 39744
rect 19208 39679 19528 39680
rect 29208 39744 29528 39745
rect 29208 39680 29216 39744
rect 29280 39680 29296 39744
rect 29360 39680 29376 39744
rect 29440 39680 29456 39744
rect 29520 39680 29528 39744
rect 29208 39679 29528 39680
rect 39208 39744 39528 39745
rect 39208 39680 39216 39744
rect 39280 39680 39296 39744
rect 39360 39680 39376 39744
rect 39440 39680 39456 39744
rect 39520 39680 39528 39744
rect 39208 39679 39528 39680
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 14208 39200 14528 39201
rect 14208 39136 14216 39200
rect 14280 39136 14296 39200
rect 14360 39136 14376 39200
rect 14440 39136 14456 39200
rect 14520 39136 14528 39200
rect 14208 39135 14528 39136
rect 24208 39200 24528 39201
rect 24208 39136 24216 39200
rect 24280 39136 24296 39200
rect 24360 39136 24376 39200
rect 24440 39136 24456 39200
rect 24520 39136 24528 39200
rect 24208 39135 24528 39136
rect 34208 39200 34528 39201
rect 34208 39136 34216 39200
rect 34280 39136 34296 39200
rect 34360 39136 34376 39200
rect 34440 39136 34456 39200
rect 34520 39136 34528 39200
rect 34208 39135 34528 39136
rect 44208 39200 44528 39201
rect 44208 39136 44216 39200
rect 44280 39136 44296 39200
rect 44360 39136 44376 39200
rect 44440 39136 44456 39200
rect 44520 39136 44528 39200
rect 44208 39135 44528 39136
rect 9208 38656 9528 38657
rect 9208 38592 9216 38656
rect 9280 38592 9296 38656
rect 9360 38592 9376 38656
rect 9440 38592 9456 38656
rect 9520 38592 9528 38656
rect 9208 38591 9528 38592
rect 19208 38656 19528 38657
rect 19208 38592 19216 38656
rect 19280 38592 19296 38656
rect 19360 38592 19376 38656
rect 19440 38592 19456 38656
rect 19520 38592 19528 38656
rect 19208 38591 19528 38592
rect 29208 38656 29528 38657
rect 29208 38592 29216 38656
rect 29280 38592 29296 38656
rect 29360 38592 29376 38656
rect 29440 38592 29456 38656
rect 29520 38592 29528 38656
rect 29208 38591 29528 38592
rect 39208 38656 39528 38657
rect 39208 38592 39216 38656
rect 39280 38592 39296 38656
rect 39360 38592 39376 38656
rect 39440 38592 39456 38656
rect 39520 38592 39528 38656
rect 39208 38591 39528 38592
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 14208 38112 14528 38113
rect 14208 38048 14216 38112
rect 14280 38048 14296 38112
rect 14360 38048 14376 38112
rect 14440 38048 14456 38112
rect 14520 38048 14528 38112
rect 14208 38047 14528 38048
rect 24208 38112 24528 38113
rect 24208 38048 24216 38112
rect 24280 38048 24296 38112
rect 24360 38048 24376 38112
rect 24440 38048 24456 38112
rect 24520 38048 24528 38112
rect 24208 38047 24528 38048
rect 34208 38112 34528 38113
rect 34208 38048 34216 38112
rect 34280 38048 34296 38112
rect 34360 38048 34376 38112
rect 34440 38048 34456 38112
rect 34520 38048 34528 38112
rect 34208 38047 34528 38048
rect 44208 38112 44528 38113
rect 44208 38048 44216 38112
rect 44280 38048 44296 38112
rect 44360 38048 44376 38112
rect 44440 38048 44456 38112
rect 44520 38048 44528 38112
rect 44208 38047 44528 38048
rect 9208 37568 9528 37569
rect 0 37498 800 37528
rect 9208 37504 9216 37568
rect 9280 37504 9296 37568
rect 9360 37504 9376 37568
rect 9440 37504 9456 37568
rect 9520 37504 9528 37568
rect 9208 37503 9528 37504
rect 19208 37568 19528 37569
rect 19208 37504 19216 37568
rect 19280 37504 19296 37568
rect 19360 37504 19376 37568
rect 19440 37504 19456 37568
rect 19520 37504 19528 37568
rect 19208 37503 19528 37504
rect 29208 37568 29528 37569
rect 29208 37504 29216 37568
rect 29280 37504 29296 37568
rect 29360 37504 29376 37568
rect 29440 37504 29456 37568
rect 29520 37504 29528 37568
rect 29208 37503 29528 37504
rect 39208 37568 39528 37569
rect 39208 37504 39216 37568
rect 39280 37504 39296 37568
rect 39360 37504 39376 37568
rect 39440 37504 39456 37568
rect 39520 37504 39528 37568
rect 39208 37503 39528 37504
rect 1853 37498 1919 37501
rect 0 37496 1919 37498
rect 0 37440 1858 37496
rect 1914 37440 1919 37496
rect 0 37438 1919 37440
rect 0 37408 800 37438
rect 1853 37435 1919 37438
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 14208 37024 14528 37025
rect 14208 36960 14216 37024
rect 14280 36960 14296 37024
rect 14360 36960 14376 37024
rect 14440 36960 14456 37024
rect 14520 36960 14528 37024
rect 14208 36959 14528 36960
rect 24208 37024 24528 37025
rect 24208 36960 24216 37024
rect 24280 36960 24296 37024
rect 24360 36960 24376 37024
rect 24440 36960 24456 37024
rect 24520 36960 24528 37024
rect 24208 36959 24528 36960
rect 34208 37024 34528 37025
rect 34208 36960 34216 37024
rect 34280 36960 34296 37024
rect 34360 36960 34376 37024
rect 34440 36960 34456 37024
rect 34520 36960 34528 37024
rect 34208 36959 34528 36960
rect 44208 37024 44528 37025
rect 44208 36960 44216 37024
rect 44280 36960 44296 37024
rect 44360 36960 44376 37024
rect 44440 36960 44456 37024
rect 44520 36960 44528 37024
rect 44208 36959 44528 36960
rect 9208 36480 9528 36481
rect 9208 36416 9216 36480
rect 9280 36416 9296 36480
rect 9360 36416 9376 36480
rect 9440 36416 9456 36480
rect 9520 36416 9528 36480
rect 9208 36415 9528 36416
rect 19208 36480 19528 36481
rect 19208 36416 19216 36480
rect 19280 36416 19296 36480
rect 19360 36416 19376 36480
rect 19440 36416 19456 36480
rect 19520 36416 19528 36480
rect 19208 36415 19528 36416
rect 29208 36480 29528 36481
rect 29208 36416 29216 36480
rect 29280 36416 29296 36480
rect 29360 36416 29376 36480
rect 29440 36416 29456 36480
rect 29520 36416 29528 36480
rect 29208 36415 29528 36416
rect 39208 36480 39528 36481
rect 39208 36416 39216 36480
rect 39280 36416 39296 36480
rect 39360 36416 39376 36480
rect 39440 36416 39456 36480
rect 39520 36416 39528 36480
rect 39208 36415 39528 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 14208 35936 14528 35937
rect 14208 35872 14216 35936
rect 14280 35872 14296 35936
rect 14360 35872 14376 35936
rect 14440 35872 14456 35936
rect 14520 35872 14528 35936
rect 14208 35871 14528 35872
rect 24208 35936 24528 35937
rect 24208 35872 24216 35936
rect 24280 35872 24296 35936
rect 24360 35872 24376 35936
rect 24440 35872 24456 35936
rect 24520 35872 24528 35936
rect 24208 35871 24528 35872
rect 34208 35936 34528 35937
rect 34208 35872 34216 35936
rect 34280 35872 34296 35936
rect 34360 35872 34376 35936
rect 34440 35872 34456 35936
rect 34520 35872 34528 35936
rect 34208 35871 34528 35872
rect 44208 35936 44528 35937
rect 44208 35872 44216 35936
rect 44280 35872 44296 35936
rect 44360 35872 44376 35936
rect 44440 35872 44456 35936
rect 44520 35872 44528 35936
rect 44208 35871 44528 35872
rect 9208 35392 9528 35393
rect 9208 35328 9216 35392
rect 9280 35328 9296 35392
rect 9360 35328 9376 35392
rect 9440 35328 9456 35392
rect 9520 35328 9528 35392
rect 9208 35327 9528 35328
rect 19208 35392 19528 35393
rect 19208 35328 19216 35392
rect 19280 35328 19296 35392
rect 19360 35328 19376 35392
rect 19440 35328 19456 35392
rect 19520 35328 19528 35392
rect 19208 35327 19528 35328
rect 29208 35392 29528 35393
rect 29208 35328 29216 35392
rect 29280 35328 29296 35392
rect 29360 35328 29376 35392
rect 29440 35328 29456 35392
rect 29520 35328 29528 35392
rect 29208 35327 29528 35328
rect 39208 35392 39528 35393
rect 39208 35328 39216 35392
rect 39280 35328 39296 35392
rect 39360 35328 39376 35392
rect 39440 35328 39456 35392
rect 39520 35328 39528 35392
rect 39208 35327 39528 35328
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 14208 34848 14528 34849
rect 14208 34784 14216 34848
rect 14280 34784 14296 34848
rect 14360 34784 14376 34848
rect 14440 34784 14456 34848
rect 14520 34784 14528 34848
rect 14208 34783 14528 34784
rect 24208 34848 24528 34849
rect 24208 34784 24216 34848
rect 24280 34784 24296 34848
rect 24360 34784 24376 34848
rect 24440 34784 24456 34848
rect 24520 34784 24528 34848
rect 24208 34783 24528 34784
rect 34208 34848 34528 34849
rect 34208 34784 34216 34848
rect 34280 34784 34296 34848
rect 34360 34784 34376 34848
rect 34440 34784 34456 34848
rect 34520 34784 34528 34848
rect 34208 34783 34528 34784
rect 44208 34848 44528 34849
rect 44208 34784 44216 34848
rect 44280 34784 44296 34848
rect 44360 34784 44376 34848
rect 44440 34784 44456 34848
rect 44520 34784 44528 34848
rect 44208 34783 44528 34784
rect 9208 34304 9528 34305
rect 9208 34240 9216 34304
rect 9280 34240 9296 34304
rect 9360 34240 9376 34304
rect 9440 34240 9456 34304
rect 9520 34240 9528 34304
rect 9208 34239 9528 34240
rect 19208 34304 19528 34305
rect 19208 34240 19216 34304
rect 19280 34240 19296 34304
rect 19360 34240 19376 34304
rect 19440 34240 19456 34304
rect 19520 34240 19528 34304
rect 19208 34239 19528 34240
rect 29208 34304 29528 34305
rect 29208 34240 29216 34304
rect 29280 34240 29296 34304
rect 29360 34240 29376 34304
rect 29440 34240 29456 34304
rect 29520 34240 29528 34304
rect 29208 34239 29528 34240
rect 39208 34304 39528 34305
rect 39208 34240 39216 34304
rect 39280 34240 39296 34304
rect 39360 34240 39376 34304
rect 39440 34240 39456 34304
rect 39520 34240 39528 34304
rect 39208 34239 39528 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 14208 33760 14528 33761
rect 14208 33696 14216 33760
rect 14280 33696 14296 33760
rect 14360 33696 14376 33760
rect 14440 33696 14456 33760
rect 14520 33696 14528 33760
rect 14208 33695 14528 33696
rect 24208 33760 24528 33761
rect 24208 33696 24216 33760
rect 24280 33696 24296 33760
rect 24360 33696 24376 33760
rect 24440 33696 24456 33760
rect 24520 33696 24528 33760
rect 24208 33695 24528 33696
rect 34208 33760 34528 33761
rect 34208 33696 34216 33760
rect 34280 33696 34296 33760
rect 34360 33696 34376 33760
rect 34440 33696 34456 33760
rect 34520 33696 34528 33760
rect 34208 33695 34528 33696
rect 44208 33760 44528 33761
rect 44208 33696 44216 33760
rect 44280 33696 44296 33760
rect 44360 33696 44376 33760
rect 44440 33696 44456 33760
rect 44520 33696 44528 33760
rect 44208 33695 44528 33696
rect 9208 33216 9528 33217
rect 9208 33152 9216 33216
rect 9280 33152 9296 33216
rect 9360 33152 9376 33216
rect 9440 33152 9456 33216
rect 9520 33152 9528 33216
rect 9208 33151 9528 33152
rect 19208 33216 19528 33217
rect 19208 33152 19216 33216
rect 19280 33152 19296 33216
rect 19360 33152 19376 33216
rect 19440 33152 19456 33216
rect 19520 33152 19528 33216
rect 19208 33151 19528 33152
rect 29208 33216 29528 33217
rect 29208 33152 29216 33216
rect 29280 33152 29296 33216
rect 29360 33152 29376 33216
rect 29440 33152 29456 33216
rect 29520 33152 29528 33216
rect 29208 33151 29528 33152
rect 39208 33216 39528 33217
rect 39208 33152 39216 33216
rect 39280 33152 39296 33216
rect 39360 33152 39376 33216
rect 39440 33152 39456 33216
rect 39520 33152 39528 33216
rect 39208 33151 39528 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 14208 32672 14528 32673
rect 14208 32608 14216 32672
rect 14280 32608 14296 32672
rect 14360 32608 14376 32672
rect 14440 32608 14456 32672
rect 14520 32608 14528 32672
rect 14208 32607 14528 32608
rect 24208 32672 24528 32673
rect 24208 32608 24216 32672
rect 24280 32608 24296 32672
rect 24360 32608 24376 32672
rect 24440 32608 24456 32672
rect 24520 32608 24528 32672
rect 24208 32607 24528 32608
rect 34208 32672 34528 32673
rect 34208 32608 34216 32672
rect 34280 32608 34296 32672
rect 34360 32608 34376 32672
rect 34440 32608 34456 32672
rect 34520 32608 34528 32672
rect 34208 32607 34528 32608
rect 44208 32672 44528 32673
rect 44208 32608 44216 32672
rect 44280 32608 44296 32672
rect 44360 32608 44376 32672
rect 44440 32608 44456 32672
rect 44520 32608 44528 32672
rect 44208 32607 44528 32608
rect 0 32466 800 32496
rect 1761 32466 1827 32469
rect 0 32464 1827 32466
rect 0 32408 1766 32464
rect 1822 32408 1827 32464
rect 0 32406 1827 32408
rect 0 32376 800 32406
rect 1761 32403 1827 32406
rect 9208 32128 9528 32129
rect 9208 32064 9216 32128
rect 9280 32064 9296 32128
rect 9360 32064 9376 32128
rect 9440 32064 9456 32128
rect 9520 32064 9528 32128
rect 9208 32063 9528 32064
rect 19208 32128 19528 32129
rect 19208 32064 19216 32128
rect 19280 32064 19296 32128
rect 19360 32064 19376 32128
rect 19440 32064 19456 32128
rect 19520 32064 19528 32128
rect 19208 32063 19528 32064
rect 29208 32128 29528 32129
rect 29208 32064 29216 32128
rect 29280 32064 29296 32128
rect 29360 32064 29376 32128
rect 29440 32064 29456 32128
rect 29520 32064 29528 32128
rect 29208 32063 29528 32064
rect 39208 32128 39528 32129
rect 39208 32064 39216 32128
rect 39280 32064 39296 32128
rect 39360 32064 39376 32128
rect 39440 32064 39456 32128
rect 39520 32064 39528 32128
rect 39208 32063 39528 32064
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 14208 31584 14528 31585
rect 14208 31520 14216 31584
rect 14280 31520 14296 31584
rect 14360 31520 14376 31584
rect 14440 31520 14456 31584
rect 14520 31520 14528 31584
rect 14208 31519 14528 31520
rect 24208 31584 24528 31585
rect 24208 31520 24216 31584
rect 24280 31520 24296 31584
rect 24360 31520 24376 31584
rect 24440 31520 24456 31584
rect 24520 31520 24528 31584
rect 24208 31519 24528 31520
rect 34208 31584 34528 31585
rect 34208 31520 34216 31584
rect 34280 31520 34296 31584
rect 34360 31520 34376 31584
rect 34440 31520 34456 31584
rect 34520 31520 34528 31584
rect 34208 31519 34528 31520
rect 44208 31584 44528 31585
rect 44208 31520 44216 31584
rect 44280 31520 44296 31584
rect 44360 31520 44376 31584
rect 44440 31520 44456 31584
rect 44520 31520 44528 31584
rect 44208 31519 44528 31520
rect 9208 31040 9528 31041
rect 9208 30976 9216 31040
rect 9280 30976 9296 31040
rect 9360 30976 9376 31040
rect 9440 30976 9456 31040
rect 9520 30976 9528 31040
rect 9208 30975 9528 30976
rect 19208 31040 19528 31041
rect 19208 30976 19216 31040
rect 19280 30976 19296 31040
rect 19360 30976 19376 31040
rect 19440 30976 19456 31040
rect 19520 30976 19528 31040
rect 19208 30975 19528 30976
rect 29208 31040 29528 31041
rect 29208 30976 29216 31040
rect 29280 30976 29296 31040
rect 29360 30976 29376 31040
rect 29440 30976 29456 31040
rect 29520 30976 29528 31040
rect 29208 30975 29528 30976
rect 39208 31040 39528 31041
rect 39208 30976 39216 31040
rect 39280 30976 39296 31040
rect 39360 30976 39376 31040
rect 39440 30976 39456 31040
rect 39520 30976 39528 31040
rect 39208 30975 39528 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 14208 30496 14528 30497
rect 14208 30432 14216 30496
rect 14280 30432 14296 30496
rect 14360 30432 14376 30496
rect 14440 30432 14456 30496
rect 14520 30432 14528 30496
rect 14208 30431 14528 30432
rect 24208 30496 24528 30497
rect 24208 30432 24216 30496
rect 24280 30432 24296 30496
rect 24360 30432 24376 30496
rect 24440 30432 24456 30496
rect 24520 30432 24528 30496
rect 24208 30431 24528 30432
rect 34208 30496 34528 30497
rect 34208 30432 34216 30496
rect 34280 30432 34296 30496
rect 34360 30432 34376 30496
rect 34440 30432 34456 30496
rect 34520 30432 34528 30496
rect 34208 30431 34528 30432
rect 44208 30496 44528 30497
rect 44208 30432 44216 30496
rect 44280 30432 44296 30496
rect 44360 30432 44376 30496
rect 44440 30432 44456 30496
rect 44520 30432 44528 30496
rect 44208 30431 44528 30432
rect 9208 29952 9528 29953
rect 9208 29888 9216 29952
rect 9280 29888 9296 29952
rect 9360 29888 9376 29952
rect 9440 29888 9456 29952
rect 9520 29888 9528 29952
rect 9208 29887 9528 29888
rect 19208 29952 19528 29953
rect 19208 29888 19216 29952
rect 19280 29888 19296 29952
rect 19360 29888 19376 29952
rect 19440 29888 19456 29952
rect 19520 29888 19528 29952
rect 19208 29887 19528 29888
rect 29208 29952 29528 29953
rect 29208 29888 29216 29952
rect 29280 29888 29296 29952
rect 29360 29888 29376 29952
rect 29440 29888 29456 29952
rect 29520 29888 29528 29952
rect 29208 29887 29528 29888
rect 39208 29952 39528 29953
rect 39208 29888 39216 29952
rect 39280 29888 39296 29952
rect 39360 29888 39376 29952
rect 39440 29888 39456 29952
rect 39520 29888 39528 29952
rect 39208 29887 39528 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 14208 29408 14528 29409
rect 14208 29344 14216 29408
rect 14280 29344 14296 29408
rect 14360 29344 14376 29408
rect 14440 29344 14456 29408
rect 14520 29344 14528 29408
rect 14208 29343 14528 29344
rect 24208 29408 24528 29409
rect 24208 29344 24216 29408
rect 24280 29344 24296 29408
rect 24360 29344 24376 29408
rect 24440 29344 24456 29408
rect 24520 29344 24528 29408
rect 24208 29343 24528 29344
rect 34208 29408 34528 29409
rect 34208 29344 34216 29408
rect 34280 29344 34296 29408
rect 34360 29344 34376 29408
rect 34440 29344 34456 29408
rect 34520 29344 34528 29408
rect 34208 29343 34528 29344
rect 44208 29408 44528 29409
rect 44208 29344 44216 29408
rect 44280 29344 44296 29408
rect 44360 29344 44376 29408
rect 44440 29344 44456 29408
rect 44520 29344 44528 29408
rect 44208 29343 44528 29344
rect 9208 28864 9528 28865
rect 9208 28800 9216 28864
rect 9280 28800 9296 28864
rect 9360 28800 9376 28864
rect 9440 28800 9456 28864
rect 9520 28800 9528 28864
rect 9208 28799 9528 28800
rect 19208 28864 19528 28865
rect 19208 28800 19216 28864
rect 19280 28800 19296 28864
rect 19360 28800 19376 28864
rect 19440 28800 19456 28864
rect 19520 28800 19528 28864
rect 19208 28799 19528 28800
rect 29208 28864 29528 28865
rect 29208 28800 29216 28864
rect 29280 28800 29296 28864
rect 29360 28800 29376 28864
rect 29440 28800 29456 28864
rect 29520 28800 29528 28864
rect 29208 28799 29528 28800
rect 39208 28864 39528 28865
rect 39208 28800 39216 28864
rect 39280 28800 39296 28864
rect 39360 28800 39376 28864
rect 39440 28800 39456 28864
rect 39520 28800 39528 28864
rect 39208 28799 39528 28800
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 14208 28320 14528 28321
rect 14208 28256 14216 28320
rect 14280 28256 14296 28320
rect 14360 28256 14376 28320
rect 14440 28256 14456 28320
rect 14520 28256 14528 28320
rect 14208 28255 14528 28256
rect 24208 28320 24528 28321
rect 24208 28256 24216 28320
rect 24280 28256 24296 28320
rect 24360 28256 24376 28320
rect 24440 28256 24456 28320
rect 24520 28256 24528 28320
rect 24208 28255 24528 28256
rect 34208 28320 34528 28321
rect 34208 28256 34216 28320
rect 34280 28256 34296 28320
rect 34360 28256 34376 28320
rect 34440 28256 34456 28320
rect 34520 28256 34528 28320
rect 34208 28255 34528 28256
rect 44208 28320 44528 28321
rect 44208 28256 44216 28320
rect 44280 28256 44296 28320
rect 44360 28256 44376 28320
rect 44440 28256 44456 28320
rect 44520 28256 44528 28320
rect 44208 28255 44528 28256
rect 9208 27776 9528 27777
rect 9208 27712 9216 27776
rect 9280 27712 9296 27776
rect 9360 27712 9376 27776
rect 9440 27712 9456 27776
rect 9520 27712 9528 27776
rect 9208 27711 9528 27712
rect 19208 27776 19528 27777
rect 19208 27712 19216 27776
rect 19280 27712 19296 27776
rect 19360 27712 19376 27776
rect 19440 27712 19456 27776
rect 19520 27712 19528 27776
rect 19208 27711 19528 27712
rect 29208 27776 29528 27777
rect 29208 27712 29216 27776
rect 29280 27712 29296 27776
rect 29360 27712 29376 27776
rect 29440 27712 29456 27776
rect 29520 27712 29528 27776
rect 29208 27711 29528 27712
rect 39208 27776 39528 27777
rect 39208 27712 39216 27776
rect 39280 27712 39296 27776
rect 39360 27712 39376 27776
rect 39440 27712 39456 27776
rect 39520 27712 39528 27776
rect 39208 27711 39528 27712
rect 0 27570 800 27600
rect 1761 27570 1827 27573
rect 0 27568 1827 27570
rect 0 27512 1766 27568
rect 1822 27512 1827 27568
rect 0 27510 1827 27512
rect 0 27480 800 27510
rect 1761 27507 1827 27510
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 14208 27232 14528 27233
rect 14208 27168 14216 27232
rect 14280 27168 14296 27232
rect 14360 27168 14376 27232
rect 14440 27168 14456 27232
rect 14520 27168 14528 27232
rect 14208 27167 14528 27168
rect 24208 27232 24528 27233
rect 24208 27168 24216 27232
rect 24280 27168 24296 27232
rect 24360 27168 24376 27232
rect 24440 27168 24456 27232
rect 24520 27168 24528 27232
rect 24208 27167 24528 27168
rect 34208 27232 34528 27233
rect 34208 27168 34216 27232
rect 34280 27168 34296 27232
rect 34360 27168 34376 27232
rect 34440 27168 34456 27232
rect 34520 27168 34528 27232
rect 34208 27167 34528 27168
rect 44208 27232 44528 27233
rect 44208 27168 44216 27232
rect 44280 27168 44296 27232
rect 44360 27168 44376 27232
rect 44440 27168 44456 27232
rect 44520 27168 44528 27232
rect 44208 27167 44528 27168
rect 9208 26688 9528 26689
rect 9208 26624 9216 26688
rect 9280 26624 9296 26688
rect 9360 26624 9376 26688
rect 9440 26624 9456 26688
rect 9520 26624 9528 26688
rect 9208 26623 9528 26624
rect 19208 26688 19528 26689
rect 19208 26624 19216 26688
rect 19280 26624 19296 26688
rect 19360 26624 19376 26688
rect 19440 26624 19456 26688
rect 19520 26624 19528 26688
rect 19208 26623 19528 26624
rect 29208 26688 29528 26689
rect 29208 26624 29216 26688
rect 29280 26624 29296 26688
rect 29360 26624 29376 26688
rect 29440 26624 29456 26688
rect 29520 26624 29528 26688
rect 29208 26623 29528 26624
rect 39208 26688 39528 26689
rect 39208 26624 39216 26688
rect 39280 26624 39296 26688
rect 39360 26624 39376 26688
rect 39440 26624 39456 26688
rect 39520 26624 39528 26688
rect 39208 26623 39528 26624
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 14208 26144 14528 26145
rect 14208 26080 14216 26144
rect 14280 26080 14296 26144
rect 14360 26080 14376 26144
rect 14440 26080 14456 26144
rect 14520 26080 14528 26144
rect 14208 26079 14528 26080
rect 24208 26144 24528 26145
rect 24208 26080 24216 26144
rect 24280 26080 24296 26144
rect 24360 26080 24376 26144
rect 24440 26080 24456 26144
rect 24520 26080 24528 26144
rect 24208 26079 24528 26080
rect 34208 26144 34528 26145
rect 34208 26080 34216 26144
rect 34280 26080 34296 26144
rect 34360 26080 34376 26144
rect 34440 26080 34456 26144
rect 34520 26080 34528 26144
rect 34208 26079 34528 26080
rect 44208 26144 44528 26145
rect 44208 26080 44216 26144
rect 44280 26080 44296 26144
rect 44360 26080 44376 26144
rect 44440 26080 44456 26144
rect 44520 26080 44528 26144
rect 44208 26079 44528 26080
rect 9208 25600 9528 25601
rect 9208 25536 9216 25600
rect 9280 25536 9296 25600
rect 9360 25536 9376 25600
rect 9440 25536 9456 25600
rect 9520 25536 9528 25600
rect 9208 25535 9528 25536
rect 19208 25600 19528 25601
rect 19208 25536 19216 25600
rect 19280 25536 19296 25600
rect 19360 25536 19376 25600
rect 19440 25536 19456 25600
rect 19520 25536 19528 25600
rect 19208 25535 19528 25536
rect 29208 25600 29528 25601
rect 29208 25536 29216 25600
rect 29280 25536 29296 25600
rect 29360 25536 29376 25600
rect 29440 25536 29456 25600
rect 29520 25536 29528 25600
rect 29208 25535 29528 25536
rect 39208 25600 39528 25601
rect 39208 25536 39216 25600
rect 39280 25536 39296 25600
rect 39360 25536 39376 25600
rect 39440 25536 39456 25600
rect 39520 25536 39528 25600
rect 39208 25535 39528 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 14208 25056 14528 25057
rect 14208 24992 14216 25056
rect 14280 24992 14296 25056
rect 14360 24992 14376 25056
rect 14440 24992 14456 25056
rect 14520 24992 14528 25056
rect 14208 24991 14528 24992
rect 24208 25056 24528 25057
rect 24208 24992 24216 25056
rect 24280 24992 24296 25056
rect 24360 24992 24376 25056
rect 24440 24992 24456 25056
rect 24520 24992 24528 25056
rect 24208 24991 24528 24992
rect 34208 25056 34528 25057
rect 34208 24992 34216 25056
rect 34280 24992 34296 25056
rect 34360 24992 34376 25056
rect 34440 24992 34456 25056
rect 34520 24992 34528 25056
rect 34208 24991 34528 24992
rect 44208 25056 44528 25057
rect 44208 24992 44216 25056
rect 44280 24992 44296 25056
rect 44360 24992 44376 25056
rect 44440 24992 44456 25056
rect 44520 24992 44528 25056
rect 44208 24991 44528 24992
rect 48129 24986 48195 24989
rect 49200 24986 50000 25016
rect 48129 24984 50000 24986
rect 48129 24928 48134 24984
rect 48190 24928 50000 24984
rect 48129 24926 50000 24928
rect 48129 24923 48195 24926
rect 49200 24896 50000 24926
rect 9208 24512 9528 24513
rect 9208 24448 9216 24512
rect 9280 24448 9296 24512
rect 9360 24448 9376 24512
rect 9440 24448 9456 24512
rect 9520 24448 9528 24512
rect 9208 24447 9528 24448
rect 19208 24512 19528 24513
rect 19208 24448 19216 24512
rect 19280 24448 19296 24512
rect 19360 24448 19376 24512
rect 19440 24448 19456 24512
rect 19520 24448 19528 24512
rect 19208 24447 19528 24448
rect 29208 24512 29528 24513
rect 29208 24448 29216 24512
rect 29280 24448 29296 24512
rect 29360 24448 29376 24512
rect 29440 24448 29456 24512
rect 29520 24448 29528 24512
rect 29208 24447 29528 24448
rect 39208 24512 39528 24513
rect 39208 24448 39216 24512
rect 39280 24448 39296 24512
rect 39360 24448 39376 24512
rect 39440 24448 39456 24512
rect 39520 24448 39528 24512
rect 39208 24447 39528 24448
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 14208 23968 14528 23969
rect 14208 23904 14216 23968
rect 14280 23904 14296 23968
rect 14360 23904 14376 23968
rect 14440 23904 14456 23968
rect 14520 23904 14528 23968
rect 14208 23903 14528 23904
rect 24208 23968 24528 23969
rect 24208 23904 24216 23968
rect 24280 23904 24296 23968
rect 24360 23904 24376 23968
rect 24440 23904 24456 23968
rect 24520 23904 24528 23968
rect 24208 23903 24528 23904
rect 34208 23968 34528 23969
rect 34208 23904 34216 23968
rect 34280 23904 34296 23968
rect 34360 23904 34376 23968
rect 34440 23904 34456 23968
rect 34520 23904 34528 23968
rect 34208 23903 34528 23904
rect 44208 23968 44528 23969
rect 44208 23904 44216 23968
rect 44280 23904 44296 23968
rect 44360 23904 44376 23968
rect 44440 23904 44456 23968
rect 44520 23904 44528 23968
rect 44208 23903 44528 23904
rect 9208 23424 9528 23425
rect 9208 23360 9216 23424
rect 9280 23360 9296 23424
rect 9360 23360 9376 23424
rect 9440 23360 9456 23424
rect 9520 23360 9528 23424
rect 9208 23359 9528 23360
rect 19208 23424 19528 23425
rect 19208 23360 19216 23424
rect 19280 23360 19296 23424
rect 19360 23360 19376 23424
rect 19440 23360 19456 23424
rect 19520 23360 19528 23424
rect 19208 23359 19528 23360
rect 29208 23424 29528 23425
rect 29208 23360 29216 23424
rect 29280 23360 29296 23424
rect 29360 23360 29376 23424
rect 29440 23360 29456 23424
rect 29520 23360 29528 23424
rect 29208 23359 29528 23360
rect 39208 23424 39528 23425
rect 39208 23360 39216 23424
rect 39280 23360 39296 23424
rect 39360 23360 39376 23424
rect 39440 23360 39456 23424
rect 39520 23360 39528 23424
rect 39208 23359 39528 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 14208 22880 14528 22881
rect 14208 22816 14216 22880
rect 14280 22816 14296 22880
rect 14360 22816 14376 22880
rect 14440 22816 14456 22880
rect 14520 22816 14528 22880
rect 14208 22815 14528 22816
rect 24208 22880 24528 22881
rect 24208 22816 24216 22880
rect 24280 22816 24296 22880
rect 24360 22816 24376 22880
rect 24440 22816 24456 22880
rect 24520 22816 24528 22880
rect 24208 22815 24528 22816
rect 34208 22880 34528 22881
rect 34208 22816 34216 22880
rect 34280 22816 34296 22880
rect 34360 22816 34376 22880
rect 34440 22816 34456 22880
rect 34520 22816 34528 22880
rect 34208 22815 34528 22816
rect 44208 22880 44528 22881
rect 44208 22816 44216 22880
rect 44280 22816 44296 22880
rect 44360 22816 44376 22880
rect 44440 22816 44456 22880
rect 44520 22816 44528 22880
rect 44208 22815 44528 22816
rect 0 22538 800 22568
rect 1761 22538 1827 22541
rect 0 22536 1827 22538
rect 0 22480 1766 22536
rect 1822 22480 1827 22536
rect 0 22478 1827 22480
rect 0 22448 800 22478
rect 1761 22475 1827 22478
rect 9208 22336 9528 22337
rect 9208 22272 9216 22336
rect 9280 22272 9296 22336
rect 9360 22272 9376 22336
rect 9440 22272 9456 22336
rect 9520 22272 9528 22336
rect 9208 22271 9528 22272
rect 19208 22336 19528 22337
rect 19208 22272 19216 22336
rect 19280 22272 19296 22336
rect 19360 22272 19376 22336
rect 19440 22272 19456 22336
rect 19520 22272 19528 22336
rect 19208 22271 19528 22272
rect 29208 22336 29528 22337
rect 29208 22272 29216 22336
rect 29280 22272 29296 22336
rect 29360 22272 29376 22336
rect 29440 22272 29456 22336
rect 29520 22272 29528 22336
rect 29208 22271 29528 22272
rect 39208 22336 39528 22337
rect 39208 22272 39216 22336
rect 39280 22272 39296 22336
rect 39360 22272 39376 22336
rect 39440 22272 39456 22336
rect 39520 22272 39528 22336
rect 39208 22271 39528 22272
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 14208 21792 14528 21793
rect 14208 21728 14216 21792
rect 14280 21728 14296 21792
rect 14360 21728 14376 21792
rect 14440 21728 14456 21792
rect 14520 21728 14528 21792
rect 14208 21727 14528 21728
rect 24208 21792 24528 21793
rect 24208 21728 24216 21792
rect 24280 21728 24296 21792
rect 24360 21728 24376 21792
rect 24440 21728 24456 21792
rect 24520 21728 24528 21792
rect 24208 21727 24528 21728
rect 34208 21792 34528 21793
rect 34208 21728 34216 21792
rect 34280 21728 34296 21792
rect 34360 21728 34376 21792
rect 34440 21728 34456 21792
rect 34520 21728 34528 21792
rect 34208 21727 34528 21728
rect 44208 21792 44528 21793
rect 44208 21728 44216 21792
rect 44280 21728 44296 21792
rect 44360 21728 44376 21792
rect 44440 21728 44456 21792
rect 44520 21728 44528 21792
rect 44208 21727 44528 21728
rect 9208 21248 9528 21249
rect 9208 21184 9216 21248
rect 9280 21184 9296 21248
rect 9360 21184 9376 21248
rect 9440 21184 9456 21248
rect 9520 21184 9528 21248
rect 9208 21183 9528 21184
rect 19208 21248 19528 21249
rect 19208 21184 19216 21248
rect 19280 21184 19296 21248
rect 19360 21184 19376 21248
rect 19440 21184 19456 21248
rect 19520 21184 19528 21248
rect 19208 21183 19528 21184
rect 29208 21248 29528 21249
rect 29208 21184 29216 21248
rect 29280 21184 29296 21248
rect 29360 21184 29376 21248
rect 29440 21184 29456 21248
rect 29520 21184 29528 21248
rect 29208 21183 29528 21184
rect 39208 21248 39528 21249
rect 39208 21184 39216 21248
rect 39280 21184 39296 21248
rect 39360 21184 39376 21248
rect 39440 21184 39456 21248
rect 39520 21184 39528 21248
rect 39208 21183 39528 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 14208 20704 14528 20705
rect 14208 20640 14216 20704
rect 14280 20640 14296 20704
rect 14360 20640 14376 20704
rect 14440 20640 14456 20704
rect 14520 20640 14528 20704
rect 14208 20639 14528 20640
rect 24208 20704 24528 20705
rect 24208 20640 24216 20704
rect 24280 20640 24296 20704
rect 24360 20640 24376 20704
rect 24440 20640 24456 20704
rect 24520 20640 24528 20704
rect 24208 20639 24528 20640
rect 34208 20704 34528 20705
rect 34208 20640 34216 20704
rect 34280 20640 34296 20704
rect 34360 20640 34376 20704
rect 34440 20640 34456 20704
rect 34520 20640 34528 20704
rect 34208 20639 34528 20640
rect 44208 20704 44528 20705
rect 44208 20640 44216 20704
rect 44280 20640 44296 20704
rect 44360 20640 44376 20704
rect 44440 20640 44456 20704
rect 44520 20640 44528 20704
rect 44208 20639 44528 20640
rect 9208 20160 9528 20161
rect 9208 20096 9216 20160
rect 9280 20096 9296 20160
rect 9360 20096 9376 20160
rect 9440 20096 9456 20160
rect 9520 20096 9528 20160
rect 9208 20095 9528 20096
rect 19208 20160 19528 20161
rect 19208 20096 19216 20160
rect 19280 20096 19296 20160
rect 19360 20096 19376 20160
rect 19440 20096 19456 20160
rect 19520 20096 19528 20160
rect 19208 20095 19528 20096
rect 29208 20160 29528 20161
rect 29208 20096 29216 20160
rect 29280 20096 29296 20160
rect 29360 20096 29376 20160
rect 29440 20096 29456 20160
rect 29520 20096 29528 20160
rect 29208 20095 29528 20096
rect 39208 20160 39528 20161
rect 39208 20096 39216 20160
rect 39280 20096 39296 20160
rect 39360 20096 39376 20160
rect 39440 20096 39456 20160
rect 39520 20096 39528 20160
rect 39208 20095 39528 20096
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 14208 19616 14528 19617
rect 14208 19552 14216 19616
rect 14280 19552 14296 19616
rect 14360 19552 14376 19616
rect 14440 19552 14456 19616
rect 14520 19552 14528 19616
rect 14208 19551 14528 19552
rect 24208 19616 24528 19617
rect 24208 19552 24216 19616
rect 24280 19552 24296 19616
rect 24360 19552 24376 19616
rect 24440 19552 24456 19616
rect 24520 19552 24528 19616
rect 24208 19551 24528 19552
rect 34208 19616 34528 19617
rect 34208 19552 34216 19616
rect 34280 19552 34296 19616
rect 34360 19552 34376 19616
rect 34440 19552 34456 19616
rect 34520 19552 34528 19616
rect 34208 19551 34528 19552
rect 44208 19616 44528 19617
rect 44208 19552 44216 19616
rect 44280 19552 44296 19616
rect 44360 19552 44376 19616
rect 44440 19552 44456 19616
rect 44520 19552 44528 19616
rect 44208 19551 44528 19552
rect 9208 19072 9528 19073
rect 9208 19008 9216 19072
rect 9280 19008 9296 19072
rect 9360 19008 9376 19072
rect 9440 19008 9456 19072
rect 9520 19008 9528 19072
rect 9208 19007 9528 19008
rect 39208 19072 39528 19073
rect 39208 19008 39216 19072
rect 39280 19008 39296 19072
rect 39360 19008 39376 19072
rect 39440 19008 39456 19072
rect 39520 19008 39528 19072
rect 39208 19007 39528 19008
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 14208 18528 14528 18529
rect 14208 18464 14216 18528
rect 14280 18464 14296 18528
rect 14360 18464 14376 18528
rect 14440 18464 14456 18528
rect 14520 18464 14528 18528
rect 14208 18463 14528 18464
rect 44208 18528 44528 18529
rect 44208 18464 44216 18528
rect 44280 18464 44296 18528
rect 44360 18464 44376 18528
rect 44440 18464 44456 18528
rect 44520 18464 44528 18528
rect 44208 18463 44528 18464
rect 9208 17984 9528 17985
rect 9208 17920 9216 17984
rect 9280 17920 9296 17984
rect 9360 17920 9376 17984
rect 9440 17920 9456 17984
rect 9520 17920 9528 17984
rect 9208 17919 9528 17920
rect 39208 17984 39528 17985
rect 39208 17920 39216 17984
rect 39280 17920 39296 17984
rect 39360 17920 39376 17984
rect 39440 17920 39456 17984
rect 39520 17920 39528 17984
rect 39208 17919 39528 17920
rect 0 17506 800 17536
rect 1853 17506 1919 17509
rect 0 17504 1919 17506
rect 0 17448 1858 17504
rect 1914 17448 1919 17504
rect 0 17446 1919 17448
rect 0 17416 800 17446
rect 1853 17443 1919 17446
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 14208 17440 14528 17441
rect 14208 17376 14216 17440
rect 14280 17376 14296 17440
rect 14360 17376 14376 17440
rect 14440 17376 14456 17440
rect 14520 17376 14528 17440
rect 14208 17375 14528 17376
rect 44208 17440 44528 17441
rect 44208 17376 44216 17440
rect 44280 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44528 17440
rect 44208 17375 44528 17376
rect 9208 16896 9528 16897
rect 9208 16832 9216 16896
rect 9280 16832 9296 16896
rect 9360 16832 9376 16896
rect 9440 16832 9456 16896
rect 9520 16832 9528 16896
rect 9208 16831 9528 16832
rect 39208 16896 39528 16897
rect 39208 16832 39216 16896
rect 39280 16832 39296 16896
rect 39360 16832 39376 16896
rect 39440 16832 39456 16896
rect 39520 16832 39528 16896
rect 39208 16831 39528 16832
rect 29208 16438 29528 16476
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 14208 16352 14528 16353
rect 14208 16288 14216 16352
rect 14280 16288 14296 16352
rect 14360 16288 14376 16352
rect 14440 16288 14456 16352
rect 14520 16288 14528 16352
rect 14208 16287 14528 16288
rect 29208 16054 29216 16438
rect 29520 16054 29528 16438
rect 44208 16352 44528 16353
rect 44208 16288 44216 16352
rect 44280 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44528 16352
rect 44208 16287 44528 16288
rect 29208 16016 29528 16054
rect 9208 15808 9528 15809
rect 9208 15744 9216 15808
rect 9280 15744 9296 15808
rect 9360 15744 9376 15808
rect 9440 15744 9456 15808
rect 9520 15744 9528 15808
rect 9208 15743 9528 15744
rect 39208 15808 39528 15809
rect 39208 15744 39216 15808
rect 39280 15744 39296 15808
rect 39360 15744 39376 15808
rect 39440 15744 39456 15808
rect 39520 15744 39528 15808
rect 39208 15743 39528 15744
rect 24208 15638 24528 15676
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 14208 15264 14528 15265
rect 14208 15200 14216 15264
rect 14280 15200 14296 15264
rect 14360 15200 14376 15264
rect 14440 15200 14456 15264
rect 14520 15200 14528 15264
rect 24208 15254 24216 15638
rect 24520 15254 24528 15638
rect 24208 15216 24528 15254
rect 44208 15264 44528 15265
rect 14208 15199 14528 15200
rect 44208 15200 44216 15264
rect 44280 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44528 15264
rect 44208 15199 44528 15200
rect 9208 14720 9528 14721
rect 9208 14656 9216 14720
rect 9280 14656 9296 14720
rect 9360 14656 9376 14720
rect 9440 14656 9456 14720
rect 9520 14656 9528 14720
rect 9208 14655 9528 14656
rect 39208 14720 39528 14721
rect 39208 14656 39216 14720
rect 39280 14656 39296 14720
rect 39360 14656 39376 14720
rect 39440 14656 39456 14720
rect 39520 14656 39528 14720
rect 39208 14655 39528 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 14208 14176 14528 14177
rect 14208 14112 14216 14176
rect 14280 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14528 14176
rect 14208 14111 14528 14112
rect 44208 14176 44528 14177
rect 44208 14112 44216 14176
rect 44280 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44528 14176
rect 44208 14111 44528 14112
rect 9208 13632 9528 13633
rect 9208 13568 9216 13632
rect 9280 13568 9296 13632
rect 9360 13568 9376 13632
rect 9440 13568 9456 13632
rect 9520 13568 9528 13632
rect 9208 13567 9528 13568
rect 39208 13632 39528 13633
rect 39208 13568 39216 13632
rect 39280 13568 39296 13632
rect 39360 13568 39376 13632
rect 39440 13568 39456 13632
rect 39520 13568 39528 13632
rect 39208 13567 39528 13568
rect 22799 13224 24426 13253
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 14208 13088 14528 13089
rect 14208 13024 14216 13088
rect 14280 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14528 13088
rect 14208 13023 14528 13024
rect 22799 13088 22840 13224
rect 23216 13219 24426 13224
rect 22799 12932 22841 13088
rect 23216 13083 24072 13219
rect 24368 13083 24426 13219
rect 23216 13068 24426 13083
rect 23217 12932 24426 13068
rect 44208 13088 44528 13089
rect 44208 13024 44216 13088
rect 44280 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44528 13088
rect 44208 13023 44528 13024
rect 22799 12902 24426 12932
rect 22799 12846 22842 12902
rect 22799 12690 22843 12846
rect 23218 12826 24426 12902
rect 23219 12690 24426 12826
rect 22799 12620 24426 12690
rect 9208 12544 9528 12545
rect 0 12474 800 12504
rect 9208 12480 9216 12544
rect 9280 12480 9296 12544
rect 9360 12480 9376 12544
rect 9440 12480 9456 12544
rect 9520 12480 9528 12544
rect 9208 12479 9528 12480
rect 39208 12544 39528 12545
rect 39208 12480 39216 12544
rect 39280 12480 39296 12544
rect 39360 12480 39376 12544
rect 39440 12480 39456 12544
rect 39520 12480 39528 12544
rect 39208 12479 39528 12480
rect 1853 12474 1919 12477
rect 0 12472 1919 12474
rect 0 12416 1858 12472
rect 1914 12416 1919 12472
rect 0 12414 1919 12416
rect 0 12384 800 12414
rect 1853 12411 1919 12414
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 14208 12000 14528 12001
rect 14208 11936 14216 12000
rect 14280 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14528 12000
rect 14208 11935 14528 11936
rect 44208 12000 44528 12001
rect 44208 11936 44216 12000
rect 44280 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44528 12000
rect 44208 11935 44528 11936
rect 24208 11907 24528 11935
rect 24208 11603 24216 11907
rect 24520 11603 24528 11907
rect 24208 11575 24528 11603
rect 34208 11907 34528 11935
rect 34208 11603 34216 11907
rect 34520 11603 34528 11907
rect 34208 11575 34528 11603
rect 9208 11456 9528 11457
rect 9208 11392 9216 11456
rect 9280 11392 9296 11456
rect 9360 11392 9376 11456
rect 9440 11392 9456 11456
rect 9520 11392 9528 11456
rect 9208 11391 9528 11392
rect 39208 11456 39528 11457
rect 39208 11392 39216 11456
rect 39280 11392 39296 11456
rect 39360 11392 39376 11456
rect 39440 11392 39456 11456
rect 39520 11392 39528 11456
rect 39208 11391 39528 11392
rect 16021 11114 16087 11117
rect 37917 11114 37983 11117
rect 16021 11112 37983 11114
rect 16021 11056 16026 11112
rect 16082 11056 37922 11112
rect 37978 11056 37983 11112
rect 16021 11054 37983 11056
rect 16021 11051 16087 11054
rect 37917 11051 37983 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 14208 10912 14528 10913
rect 14208 10848 14216 10912
rect 14280 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14528 10912
rect 14208 10847 14528 10848
rect 44208 10912 44528 10913
rect 44208 10848 44216 10912
rect 44280 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44528 10912
rect 44208 10847 44528 10848
rect 29208 10633 29528 10661
rect 9208 10368 9528 10369
rect 9208 10304 9216 10368
rect 9280 10304 9296 10368
rect 9360 10304 9376 10368
rect 9440 10304 9456 10368
rect 9520 10304 9528 10368
rect 9208 10303 9528 10304
rect 29208 10329 29216 10633
rect 29520 10329 29528 10633
rect 29208 10301 29528 10329
rect 39208 10368 39528 10369
rect 39208 10304 39216 10368
rect 39280 10304 39296 10368
rect 39360 10304 39376 10368
rect 39440 10304 39456 10368
rect 39520 10304 39528 10368
rect 39208 10303 39528 10304
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 14208 9824 14528 9825
rect 14208 9760 14216 9824
rect 14280 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14528 9824
rect 14208 9759 14528 9760
rect 44208 9824 44528 9825
rect 44208 9760 44216 9824
rect 44280 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44528 9824
rect 44208 9759 44528 9760
rect 24208 9358 24528 9386
rect 9208 9280 9528 9281
rect 9208 9216 9216 9280
rect 9280 9216 9296 9280
rect 9360 9216 9376 9280
rect 9440 9216 9456 9280
rect 9520 9216 9528 9280
rect 9208 9215 9528 9216
rect 24208 9054 24216 9358
rect 24520 9054 24528 9358
rect 24208 9026 24528 9054
rect 34208 9358 34528 9386
rect 34208 9054 34216 9358
rect 34520 9054 34528 9358
rect 39208 9280 39528 9281
rect 39208 9216 39216 9280
rect 39280 9216 39296 9280
rect 39360 9216 39376 9280
rect 39440 9216 39456 9280
rect 39520 9216 39528 9280
rect 39208 9215 39528 9216
rect 34208 9026 34528 9054
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 14208 8736 14528 8737
rect 14208 8672 14216 8736
rect 14280 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14528 8736
rect 14208 8671 14528 8672
rect 44208 8736 44528 8737
rect 44208 8672 44216 8736
rect 44280 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44528 8736
rect 44208 8671 44528 8672
rect 48129 8394 48195 8397
rect 49200 8394 50000 8424
rect 48129 8392 50000 8394
rect 48129 8336 48134 8392
rect 48190 8336 50000 8392
rect 48129 8334 50000 8336
rect 48129 8331 48195 8334
rect 49200 8304 50000 8334
rect 9208 8192 9528 8193
rect 9208 8128 9216 8192
rect 9280 8128 9296 8192
rect 9360 8128 9376 8192
rect 9440 8128 9456 8192
rect 9520 8128 9528 8192
rect 9208 8127 9528 8128
rect 39208 8192 39528 8193
rect 39208 8128 39216 8192
rect 39280 8128 39296 8192
rect 39360 8128 39376 8192
rect 39440 8128 39456 8192
rect 39520 8128 39528 8192
rect 39208 8127 39528 8128
rect 29208 8083 29528 8111
rect 29208 7779 29216 8083
rect 29520 7779 29528 8083
rect 29208 7751 29528 7779
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 14208 7648 14528 7649
rect 14208 7584 14216 7648
rect 14280 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14528 7648
rect 14208 7583 14528 7584
rect 44208 7648 44528 7649
rect 44208 7584 44216 7648
rect 44280 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44528 7648
rect 44208 7583 44528 7584
rect 0 7442 800 7472
rect 1761 7442 1827 7445
rect 0 7440 1827 7442
rect 0 7384 1766 7440
rect 1822 7384 1827 7440
rect 0 7382 1827 7384
rect 0 7352 800 7382
rect 1761 7379 1827 7382
rect 9208 7104 9528 7105
rect 9208 7040 9216 7104
rect 9280 7040 9296 7104
rect 9360 7040 9376 7104
rect 9440 7040 9456 7104
rect 9520 7040 9528 7104
rect 9208 7039 9528 7040
rect 39208 7104 39528 7105
rect 39208 7040 39216 7104
rect 39280 7040 39296 7104
rect 39360 7040 39376 7104
rect 39440 7040 39456 7104
rect 39520 7040 39528 7104
rect 39208 7039 39528 7040
rect 18045 7034 18111 7037
rect 21817 7034 21883 7037
rect 18045 7032 21883 7034
rect 18045 6976 18050 7032
rect 18106 6976 21822 7032
rect 21878 6976 21883 7032
rect 18045 6974 21883 6976
rect 18045 6971 18111 6974
rect 21817 6971 21883 6974
rect 24208 6809 24528 6837
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 14208 6560 14528 6561
rect 14208 6496 14216 6560
rect 14280 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14528 6560
rect 14208 6495 14528 6496
rect 24208 6505 24216 6809
rect 24520 6505 24528 6809
rect 24208 6477 24528 6505
rect 34208 6809 34528 6837
rect 34208 6505 34216 6809
rect 34520 6505 34528 6809
rect 34208 6477 34528 6505
rect 44208 6560 44528 6561
rect 44208 6496 44216 6560
rect 44280 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44528 6560
rect 44208 6495 44528 6496
rect 21817 6354 21883 6357
rect 34605 6354 34671 6357
rect 21817 6352 34671 6354
rect 21817 6296 21822 6352
rect 21878 6296 34610 6352
rect 34666 6296 34671 6352
rect 21817 6294 34671 6296
rect 21817 6291 21883 6294
rect 34605 6291 34671 6294
rect 21725 6218 21791 6221
rect 21725 6216 22110 6218
rect 21725 6160 21730 6216
rect 21786 6160 22110 6216
rect 21725 6158 22110 6160
rect 21725 6155 21791 6158
rect 9208 6016 9528 6017
rect 9208 5952 9216 6016
rect 9280 5952 9296 6016
rect 9360 5952 9376 6016
rect 9440 5952 9456 6016
rect 9520 5952 9528 6016
rect 9208 5951 9528 5952
rect 22050 5946 22110 6158
rect 24945 6082 25011 6085
rect 32949 6082 33015 6085
rect 24945 6080 33015 6082
rect 24945 6024 24950 6080
rect 25006 6024 32954 6080
rect 33010 6024 33015 6080
rect 24945 6022 33015 6024
rect 24945 6019 25011 6022
rect 32949 6019 33015 6022
rect 39208 6016 39528 6017
rect 39208 5952 39216 6016
rect 39280 5952 39296 6016
rect 39360 5952 39376 6016
rect 39440 5952 39456 6016
rect 39520 5952 39528 6016
rect 39208 5951 39528 5952
rect 37273 5946 37339 5949
rect 22050 5944 37339 5946
rect 22050 5888 37278 5944
rect 37334 5888 37339 5944
rect 22050 5886 37339 5888
rect 37273 5883 37339 5886
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 14208 5472 14528 5473
rect 14208 5408 14216 5472
rect 14280 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14528 5472
rect 14208 5407 14528 5408
rect 44208 5472 44528 5473
rect 44208 5408 44216 5472
rect 44280 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44528 5472
rect 44208 5407 44528 5408
rect 9208 4928 9528 4929
rect 9208 4864 9216 4928
rect 9280 4864 9296 4928
rect 9360 4864 9376 4928
rect 9440 4864 9456 4928
rect 9520 4864 9528 4928
rect 9208 4863 9528 4864
rect 39208 4928 39528 4929
rect 39208 4864 39216 4928
rect 39280 4864 39296 4928
rect 39360 4864 39376 4928
rect 39440 4864 39456 4928
rect 39520 4864 39528 4928
rect 39208 4863 39528 4864
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 14208 4384 14528 4385
rect 14208 4320 14216 4384
rect 14280 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14528 4384
rect 14208 4319 14528 4320
rect 44208 4384 44528 4385
rect 44208 4320 44216 4384
rect 44280 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44528 4384
rect 44208 4319 44528 4320
rect 9208 3840 9528 3841
rect 9208 3776 9216 3840
rect 9280 3776 9296 3840
rect 9360 3776 9376 3840
rect 9440 3776 9456 3840
rect 9520 3776 9528 3840
rect 9208 3775 9528 3776
rect 39208 3840 39528 3841
rect 39208 3776 39216 3840
rect 39280 3776 39296 3840
rect 39360 3776 39376 3840
rect 39440 3776 39456 3840
rect 39520 3776 39528 3840
rect 39208 3775 39528 3776
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 14208 3296 14528 3297
rect 14208 3232 14216 3296
rect 14280 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14528 3296
rect 44208 3296 44528 3297
rect 14208 3231 14528 3232
rect 24208 3222 24528 3260
rect 44208 3232 44216 3296
rect 44280 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44528 3296
rect 44208 3231 44528 3232
rect 24208 2838 24216 3222
rect 24520 2838 24528 3222
rect 24208 2800 24528 2838
rect 9208 2752 9528 2753
rect 9208 2688 9216 2752
rect 9280 2688 9296 2752
rect 9360 2688 9376 2752
rect 9440 2688 9456 2752
rect 9520 2688 9528 2752
rect 9208 2687 9528 2688
rect 39208 2752 39528 2753
rect 39208 2688 39216 2752
rect 39280 2688 39296 2752
rect 39360 2688 39376 2752
rect 39440 2688 39456 2752
rect 39520 2688 39528 2752
rect 39208 2687 39528 2688
rect 0 2546 800 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 0 2456 800 2486
rect 1393 2483 1459 2486
rect 29208 2430 29528 2460
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 14208 2208 14528 2209
rect 14208 2144 14216 2208
rect 14280 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14528 2208
rect 29208 2206 29216 2430
rect 29520 2206 29528 2430
rect 29208 2176 29528 2206
rect 44208 2208 44528 2209
rect 14208 2143 14528 2144
rect 44208 2144 44216 2208
rect 44280 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44528 2208
rect 44208 2143 44528 2144
<< via3 >>
rect 9216 47356 9280 47360
rect 9216 47300 9220 47356
rect 9220 47300 9276 47356
rect 9276 47300 9280 47356
rect 9216 47296 9280 47300
rect 9296 47356 9360 47360
rect 9296 47300 9300 47356
rect 9300 47300 9356 47356
rect 9356 47300 9360 47356
rect 9296 47296 9360 47300
rect 9376 47356 9440 47360
rect 9376 47300 9380 47356
rect 9380 47300 9436 47356
rect 9436 47300 9440 47356
rect 9376 47296 9440 47300
rect 9456 47356 9520 47360
rect 9456 47300 9460 47356
rect 9460 47300 9516 47356
rect 9516 47300 9520 47356
rect 9456 47296 9520 47300
rect 19216 47356 19280 47360
rect 19216 47300 19220 47356
rect 19220 47300 19276 47356
rect 19276 47300 19280 47356
rect 19216 47296 19280 47300
rect 19296 47356 19360 47360
rect 19296 47300 19300 47356
rect 19300 47300 19356 47356
rect 19356 47300 19360 47356
rect 19296 47296 19360 47300
rect 19376 47356 19440 47360
rect 19376 47300 19380 47356
rect 19380 47300 19436 47356
rect 19436 47300 19440 47356
rect 19376 47296 19440 47300
rect 19456 47356 19520 47360
rect 19456 47300 19460 47356
rect 19460 47300 19516 47356
rect 19516 47300 19520 47356
rect 19456 47296 19520 47300
rect 29216 47356 29280 47360
rect 29216 47300 29220 47356
rect 29220 47300 29276 47356
rect 29276 47300 29280 47356
rect 29216 47296 29280 47300
rect 29296 47356 29360 47360
rect 29296 47300 29300 47356
rect 29300 47300 29356 47356
rect 29356 47300 29360 47356
rect 29296 47296 29360 47300
rect 29376 47356 29440 47360
rect 29376 47300 29380 47356
rect 29380 47300 29436 47356
rect 29436 47300 29440 47356
rect 29376 47296 29440 47300
rect 29456 47356 29520 47360
rect 29456 47300 29460 47356
rect 29460 47300 29516 47356
rect 29516 47300 29520 47356
rect 29456 47296 29520 47300
rect 39216 47356 39280 47360
rect 39216 47300 39220 47356
rect 39220 47300 39276 47356
rect 39276 47300 39280 47356
rect 39216 47296 39280 47300
rect 39296 47356 39360 47360
rect 39296 47300 39300 47356
rect 39300 47300 39356 47356
rect 39356 47300 39360 47356
rect 39296 47296 39360 47300
rect 39376 47356 39440 47360
rect 39376 47300 39380 47356
rect 39380 47300 39436 47356
rect 39436 47300 39440 47356
rect 39376 47296 39440 47300
rect 39456 47356 39520 47360
rect 39456 47300 39460 47356
rect 39460 47300 39516 47356
rect 39516 47300 39520 47356
rect 39456 47296 39520 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 14216 46812 14280 46816
rect 14216 46756 14220 46812
rect 14220 46756 14276 46812
rect 14276 46756 14280 46812
rect 14216 46752 14280 46756
rect 14296 46812 14360 46816
rect 14296 46756 14300 46812
rect 14300 46756 14356 46812
rect 14356 46756 14360 46812
rect 14296 46752 14360 46756
rect 14376 46812 14440 46816
rect 14376 46756 14380 46812
rect 14380 46756 14436 46812
rect 14436 46756 14440 46812
rect 14376 46752 14440 46756
rect 14456 46812 14520 46816
rect 14456 46756 14460 46812
rect 14460 46756 14516 46812
rect 14516 46756 14520 46812
rect 14456 46752 14520 46756
rect 24216 46812 24280 46816
rect 24216 46756 24220 46812
rect 24220 46756 24276 46812
rect 24276 46756 24280 46812
rect 24216 46752 24280 46756
rect 24296 46812 24360 46816
rect 24296 46756 24300 46812
rect 24300 46756 24356 46812
rect 24356 46756 24360 46812
rect 24296 46752 24360 46756
rect 24376 46812 24440 46816
rect 24376 46756 24380 46812
rect 24380 46756 24436 46812
rect 24436 46756 24440 46812
rect 24376 46752 24440 46756
rect 24456 46812 24520 46816
rect 24456 46756 24460 46812
rect 24460 46756 24516 46812
rect 24516 46756 24520 46812
rect 24456 46752 24520 46756
rect 34216 46812 34280 46816
rect 34216 46756 34220 46812
rect 34220 46756 34276 46812
rect 34276 46756 34280 46812
rect 34216 46752 34280 46756
rect 34296 46812 34360 46816
rect 34296 46756 34300 46812
rect 34300 46756 34356 46812
rect 34356 46756 34360 46812
rect 34296 46752 34360 46756
rect 34376 46812 34440 46816
rect 34376 46756 34380 46812
rect 34380 46756 34436 46812
rect 34436 46756 34440 46812
rect 34376 46752 34440 46756
rect 34456 46812 34520 46816
rect 34456 46756 34460 46812
rect 34460 46756 34516 46812
rect 34516 46756 34520 46812
rect 34456 46752 34520 46756
rect 44216 46812 44280 46816
rect 44216 46756 44220 46812
rect 44220 46756 44276 46812
rect 44276 46756 44280 46812
rect 44216 46752 44280 46756
rect 44296 46812 44360 46816
rect 44296 46756 44300 46812
rect 44300 46756 44356 46812
rect 44356 46756 44360 46812
rect 44296 46752 44360 46756
rect 44376 46812 44440 46816
rect 44376 46756 44380 46812
rect 44380 46756 44436 46812
rect 44436 46756 44440 46812
rect 44376 46752 44440 46756
rect 44456 46812 44520 46816
rect 44456 46756 44460 46812
rect 44460 46756 44516 46812
rect 44516 46756 44520 46812
rect 44456 46752 44520 46756
rect 9216 46268 9280 46272
rect 9216 46212 9220 46268
rect 9220 46212 9276 46268
rect 9276 46212 9280 46268
rect 9216 46208 9280 46212
rect 9296 46268 9360 46272
rect 9296 46212 9300 46268
rect 9300 46212 9356 46268
rect 9356 46212 9360 46268
rect 9296 46208 9360 46212
rect 9376 46268 9440 46272
rect 9376 46212 9380 46268
rect 9380 46212 9436 46268
rect 9436 46212 9440 46268
rect 9376 46208 9440 46212
rect 9456 46268 9520 46272
rect 9456 46212 9460 46268
rect 9460 46212 9516 46268
rect 9516 46212 9520 46268
rect 9456 46208 9520 46212
rect 19216 46268 19280 46272
rect 19216 46212 19220 46268
rect 19220 46212 19276 46268
rect 19276 46212 19280 46268
rect 19216 46208 19280 46212
rect 19296 46268 19360 46272
rect 19296 46212 19300 46268
rect 19300 46212 19356 46268
rect 19356 46212 19360 46268
rect 19296 46208 19360 46212
rect 19376 46268 19440 46272
rect 19376 46212 19380 46268
rect 19380 46212 19436 46268
rect 19436 46212 19440 46268
rect 19376 46208 19440 46212
rect 19456 46268 19520 46272
rect 19456 46212 19460 46268
rect 19460 46212 19516 46268
rect 19516 46212 19520 46268
rect 19456 46208 19520 46212
rect 29216 46268 29280 46272
rect 29216 46212 29220 46268
rect 29220 46212 29276 46268
rect 29276 46212 29280 46268
rect 29216 46208 29280 46212
rect 29296 46268 29360 46272
rect 29296 46212 29300 46268
rect 29300 46212 29356 46268
rect 29356 46212 29360 46268
rect 29296 46208 29360 46212
rect 29376 46268 29440 46272
rect 29376 46212 29380 46268
rect 29380 46212 29436 46268
rect 29436 46212 29440 46268
rect 29376 46208 29440 46212
rect 29456 46268 29520 46272
rect 29456 46212 29460 46268
rect 29460 46212 29516 46268
rect 29516 46212 29520 46268
rect 29456 46208 29520 46212
rect 39216 46268 39280 46272
rect 39216 46212 39220 46268
rect 39220 46212 39276 46268
rect 39276 46212 39280 46268
rect 39216 46208 39280 46212
rect 39296 46268 39360 46272
rect 39296 46212 39300 46268
rect 39300 46212 39356 46268
rect 39356 46212 39360 46268
rect 39296 46208 39360 46212
rect 39376 46268 39440 46272
rect 39376 46212 39380 46268
rect 39380 46212 39436 46268
rect 39436 46212 39440 46268
rect 39376 46208 39440 46212
rect 39456 46268 39520 46272
rect 39456 46212 39460 46268
rect 39460 46212 39516 46268
rect 39516 46212 39520 46268
rect 39456 46208 39520 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 14216 45724 14280 45728
rect 14216 45668 14220 45724
rect 14220 45668 14276 45724
rect 14276 45668 14280 45724
rect 14216 45664 14280 45668
rect 14296 45724 14360 45728
rect 14296 45668 14300 45724
rect 14300 45668 14356 45724
rect 14356 45668 14360 45724
rect 14296 45664 14360 45668
rect 14376 45724 14440 45728
rect 14376 45668 14380 45724
rect 14380 45668 14436 45724
rect 14436 45668 14440 45724
rect 14376 45664 14440 45668
rect 14456 45724 14520 45728
rect 14456 45668 14460 45724
rect 14460 45668 14516 45724
rect 14516 45668 14520 45724
rect 14456 45664 14520 45668
rect 24216 45724 24280 45728
rect 24216 45668 24220 45724
rect 24220 45668 24276 45724
rect 24276 45668 24280 45724
rect 24216 45664 24280 45668
rect 24296 45724 24360 45728
rect 24296 45668 24300 45724
rect 24300 45668 24356 45724
rect 24356 45668 24360 45724
rect 24296 45664 24360 45668
rect 24376 45724 24440 45728
rect 24376 45668 24380 45724
rect 24380 45668 24436 45724
rect 24436 45668 24440 45724
rect 24376 45664 24440 45668
rect 24456 45724 24520 45728
rect 24456 45668 24460 45724
rect 24460 45668 24516 45724
rect 24516 45668 24520 45724
rect 24456 45664 24520 45668
rect 34216 45724 34280 45728
rect 34216 45668 34220 45724
rect 34220 45668 34276 45724
rect 34276 45668 34280 45724
rect 34216 45664 34280 45668
rect 34296 45724 34360 45728
rect 34296 45668 34300 45724
rect 34300 45668 34356 45724
rect 34356 45668 34360 45724
rect 34296 45664 34360 45668
rect 34376 45724 34440 45728
rect 34376 45668 34380 45724
rect 34380 45668 34436 45724
rect 34436 45668 34440 45724
rect 34376 45664 34440 45668
rect 34456 45724 34520 45728
rect 34456 45668 34460 45724
rect 34460 45668 34516 45724
rect 34516 45668 34520 45724
rect 34456 45664 34520 45668
rect 44216 45724 44280 45728
rect 44216 45668 44220 45724
rect 44220 45668 44276 45724
rect 44276 45668 44280 45724
rect 44216 45664 44280 45668
rect 44296 45724 44360 45728
rect 44296 45668 44300 45724
rect 44300 45668 44356 45724
rect 44356 45668 44360 45724
rect 44296 45664 44360 45668
rect 44376 45724 44440 45728
rect 44376 45668 44380 45724
rect 44380 45668 44436 45724
rect 44436 45668 44440 45724
rect 44376 45664 44440 45668
rect 44456 45724 44520 45728
rect 44456 45668 44460 45724
rect 44460 45668 44516 45724
rect 44516 45668 44520 45724
rect 44456 45664 44520 45668
rect 9216 45180 9280 45184
rect 9216 45124 9220 45180
rect 9220 45124 9276 45180
rect 9276 45124 9280 45180
rect 9216 45120 9280 45124
rect 9296 45180 9360 45184
rect 9296 45124 9300 45180
rect 9300 45124 9356 45180
rect 9356 45124 9360 45180
rect 9296 45120 9360 45124
rect 9376 45180 9440 45184
rect 9376 45124 9380 45180
rect 9380 45124 9436 45180
rect 9436 45124 9440 45180
rect 9376 45120 9440 45124
rect 9456 45180 9520 45184
rect 9456 45124 9460 45180
rect 9460 45124 9516 45180
rect 9516 45124 9520 45180
rect 9456 45120 9520 45124
rect 19216 45180 19280 45184
rect 19216 45124 19220 45180
rect 19220 45124 19276 45180
rect 19276 45124 19280 45180
rect 19216 45120 19280 45124
rect 19296 45180 19360 45184
rect 19296 45124 19300 45180
rect 19300 45124 19356 45180
rect 19356 45124 19360 45180
rect 19296 45120 19360 45124
rect 19376 45180 19440 45184
rect 19376 45124 19380 45180
rect 19380 45124 19436 45180
rect 19436 45124 19440 45180
rect 19376 45120 19440 45124
rect 19456 45180 19520 45184
rect 19456 45124 19460 45180
rect 19460 45124 19516 45180
rect 19516 45124 19520 45180
rect 19456 45120 19520 45124
rect 29216 45180 29280 45184
rect 29216 45124 29220 45180
rect 29220 45124 29276 45180
rect 29276 45124 29280 45180
rect 29216 45120 29280 45124
rect 29296 45180 29360 45184
rect 29296 45124 29300 45180
rect 29300 45124 29356 45180
rect 29356 45124 29360 45180
rect 29296 45120 29360 45124
rect 29376 45180 29440 45184
rect 29376 45124 29380 45180
rect 29380 45124 29436 45180
rect 29436 45124 29440 45180
rect 29376 45120 29440 45124
rect 29456 45180 29520 45184
rect 29456 45124 29460 45180
rect 29460 45124 29516 45180
rect 29516 45124 29520 45180
rect 29456 45120 29520 45124
rect 39216 45180 39280 45184
rect 39216 45124 39220 45180
rect 39220 45124 39276 45180
rect 39276 45124 39280 45180
rect 39216 45120 39280 45124
rect 39296 45180 39360 45184
rect 39296 45124 39300 45180
rect 39300 45124 39356 45180
rect 39356 45124 39360 45180
rect 39296 45120 39360 45124
rect 39376 45180 39440 45184
rect 39376 45124 39380 45180
rect 39380 45124 39436 45180
rect 39436 45124 39440 45180
rect 39376 45120 39440 45124
rect 39456 45180 39520 45184
rect 39456 45124 39460 45180
rect 39460 45124 39516 45180
rect 39516 45124 39520 45180
rect 39456 45120 39520 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 14216 44636 14280 44640
rect 14216 44580 14220 44636
rect 14220 44580 14276 44636
rect 14276 44580 14280 44636
rect 14216 44576 14280 44580
rect 14296 44636 14360 44640
rect 14296 44580 14300 44636
rect 14300 44580 14356 44636
rect 14356 44580 14360 44636
rect 14296 44576 14360 44580
rect 14376 44636 14440 44640
rect 14376 44580 14380 44636
rect 14380 44580 14436 44636
rect 14436 44580 14440 44636
rect 14376 44576 14440 44580
rect 14456 44636 14520 44640
rect 14456 44580 14460 44636
rect 14460 44580 14516 44636
rect 14516 44580 14520 44636
rect 14456 44576 14520 44580
rect 24216 44636 24280 44640
rect 24216 44580 24220 44636
rect 24220 44580 24276 44636
rect 24276 44580 24280 44636
rect 24216 44576 24280 44580
rect 24296 44636 24360 44640
rect 24296 44580 24300 44636
rect 24300 44580 24356 44636
rect 24356 44580 24360 44636
rect 24296 44576 24360 44580
rect 24376 44636 24440 44640
rect 24376 44580 24380 44636
rect 24380 44580 24436 44636
rect 24436 44580 24440 44636
rect 24376 44576 24440 44580
rect 24456 44636 24520 44640
rect 24456 44580 24460 44636
rect 24460 44580 24516 44636
rect 24516 44580 24520 44636
rect 24456 44576 24520 44580
rect 34216 44636 34280 44640
rect 34216 44580 34220 44636
rect 34220 44580 34276 44636
rect 34276 44580 34280 44636
rect 34216 44576 34280 44580
rect 34296 44636 34360 44640
rect 34296 44580 34300 44636
rect 34300 44580 34356 44636
rect 34356 44580 34360 44636
rect 34296 44576 34360 44580
rect 34376 44636 34440 44640
rect 34376 44580 34380 44636
rect 34380 44580 34436 44636
rect 34436 44580 34440 44636
rect 34376 44576 34440 44580
rect 34456 44636 34520 44640
rect 34456 44580 34460 44636
rect 34460 44580 34516 44636
rect 34516 44580 34520 44636
rect 34456 44576 34520 44580
rect 44216 44636 44280 44640
rect 44216 44580 44220 44636
rect 44220 44580 44276 44636
rect 44276 44580 44280 44636
rect 44216 44576 44280 44580
rect 44296 44636 44360 44640
rect 44296 44580 44300 44636
rect 44300 44580 44356 44636
rect 44356 44580 44360 44636
rect 44296 44576 44360 44580
rect 44376 44636 44440 44640
rect 44376 44580 44380 44636
rect 44380 44580 44436 44636
rect 44436 44580 44440 44636
rect 44376 44576 44440 44580
rect 44456 44636 44520 44640
rect 44456 44580 44460 44636
rect 44460 44580 44516 44636
rect 44516 44580 44520 44636
rect 44456 44576 44520 44580
rect 9216 44092 9280 44096
rect 9216 44036 9220 44092
rect 9220 44036 9276 44092
rect 9276 44036 9280 44092
rect 9216 44032 9280 44036
rect 9296 44092 9360 44096
rect 9296 44036 9300 44092
rect 9300 44036 9356 44092
rect 9356 44036 9360 44092
rect 9296 44032 9360 44036
rect 9376 44092 9440 44096
rect 9376 44036 9380 44092
rect 9380 44036 9436 44092
rect 9436 44036 9440 44092
rect 9376 44032 9440 44036
rect 9456 44092 9520 44096
rect 9456 44036 9460 44092
rect 9460 44036 9516 44092
rect 9516 44036 9520 44092
rect 9456 44032 9520 44036
rect 19216 44092 19280 44096
rect 19216 44036 19220 44092
rect 19220 44036 19276 44092
rect 19276 44036 19280 44092
rect 19216 44032 19280 44036
rect 19296 44092 19360 44096
rect 19296 44036 19300 44092
rect 19300 44036 19356 44092
rect 19356 44036 19360 44092
rect 19296 44032 19360 44036
rect 19376 44092 19440 44096
rect 19376 44036 19380 44092
rect 19380 44036 19436 44092
rect 19436 44036 19440 44092
rect 19376 44032 19440 44036
rect 19456 44092 19520 44096
rect 19456 44036 19460 44092
rect 19460 44036 19516 44092
rect 19516 44036 19520 44092
rect 19456 44032 19520 44036
rect 29216 44092 29280 44096
rect 29216 44036 29220 44092
rect 29220 44036 29276 44092
rect 29276 44036 29280 44092
rect 29216 44032 29280 44036
rect 29296 44092 29360 44096
rect 29296 44036 29300 44092
rect 29300 44036 29356 44092
rect 29356 44036 29360 44092
rect 29296 44032 29360 44036
rect 29376 44092 29440 44096
rect 29376 44036 29380 44092
rect 29380 44036 29436 44092
rect 29436 44036 29440 44092
rect 29376 44032 29440 44036
rect 29456 44092 29520 44096
rect 29456 44036 29460 44092
rect 29460 44036 29516 44092
rect 29516 44036 29520 44092
rect 29456 44032 29520 44036
rect 39216 44092 39280 44096
rect 39216 44036 39220 44092
rect 39220 44036 39276 44092
rect 39276 44036 39280 44092
rect 39216 44032 39280 44036
rect 39296 44092 39360 44096
rect 39296 44036 39300 44092
rect 39300 44036 39356 44092
rect 39356 44036 39360 44092
rect 39296 44032 39360 44036
rect 39376 44092 39440 44096
rect 39376 44036 39380 44092
rect 39380 44036 39436 44092
rect 39436 44036 39440 44092
rect 39376 44032 39440 44036
rect 39456 44092 39520 44096
rect 39456 44036 39460 44092
rect 39460 44036 39516 44092
rect 39516 44036 39520 44092
rect 39456 44032 39520 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 14216 43548 14280 43552
rect 14216 43492 14220 43548
rect 14220 43492 14276 43548
rect 14276 43492 14280 43548
rect 14216 43488 14280 43492
rect 14296 43548 14360 43552
rect 14296 43492 14300 43548
rect 14300 43492 14356 43548
rect 14356 43492 14360 43548
rect 14296 43488 14360 43492
rect 14376 43548 14440 43552
rect 14376 43492 14380 43548
rect 14380 43492 14436 43548
rect 14436 43492 14440 43548
rect 14376 43488 14440 43492
rect 14456 43548 14520 43552
rect 14456 43492 14460 43548
rect 14460 43492 14516 43548
rect 14516 43492 14520 43548
rect 14456 43488 14520 43492
rect 24216 43548 24280 43552
rect 24216 43492 24220 43548
rect 24220 43492 24276 43548
rect 24276 43492 24280 43548
rect 24216 43488 24280 43492
rect 24296 43548 24360 43552
rect 24296 43492 24300 43548
rect 24300 43492 24356 43548
rect 24356 43492 24360 43548
rect 24296 43488 24360 43492
rect 24376 43548 24440 43552
rect 24376 43492 24380 43548
rect 24380 43492 24436 43548
rect 24436 43492 24440 43548
rect 24376 43488 24440 43492
rect 24456 43548 24520 43552
rect 24456 43492 24460 43548
rect 24460 43492 24516 43548
rect 24516 43492 24520 43548
rect 24456 43488 24520 43492
rect 34216 43548 34280 43552
rect 34216 43492 34220 43548
rect 34220 43492 34276 43548
rect 34276 43492 34280 43548
rect 34216 43488 34280 43492
rect 34296 43548 34360 43552
rect 34296 43492 34300 43548
rect 34300 43492 34356 43548
rect 34356 43492 34360 43548
rect 34296 43488 34360 43492
rect 34376 43548 34440 43552
rect 34376 43492 34380 43548
rect 34380 43492 34436 43548
rect 34436 43492 34440 43548
rect 34376 43488 34440 43492
rect 34456 43548 34520 43552
rect 34456 43492 34460 43548
rect 34460 43492 34516 43548
rect 34516 43492 34520 43548
rect 34456 43488 34520 43492
rect 44216 43548 44280 43552
rect 44216 43492 44220 43548
rect 44220 43492 44276 43548
rect 44276 43492 44280 43548
rect 44216 43488 44280 43492
rect 44296 43548 44360 43552
rect 44296 43492 44300 43548
rect 44300 43492 44356 43548
rect 44356 43492 44360 43548
rect 44296 43488 44360 43492
rect 44376 43548 44440 43552
rect 44376 43492 44380 43548
rect 44380 43492 44436 43548
rect 44436 43492 44440 43548
rect 44376 43488 44440 43492
rect 44456 43548 44520 43552
rect 44456 43492 44460 43548
rect 44460 43492 44516 43548
rect 44516 43492 44520 43548
rect 44456 43488 44520 43492
rect 9216 43004 9280 43008
rect 9216 42948 9220 43004
rect 9220 42948 9276 43004
rect 9276 42948 9280 43004
rect 9216 42944 9280 42948
rect 9296 43004 9360 43008
rect 9296 42948 9300 43004
rect 9300 42948 9356 43004
rect 9356 42948 9360 43004
rect 9296 42944 9360 42948
rect 9376 43004 9440 43008
rect 9376 42948 9380 43004
rect 9380 42948 9436 43004
rect 9436 42948 9440 43004
rect 9376 42944 9440 42948
rect 9456 43004 9520 43008
rect 9456 42948 9460 43004
rect 9460 42948 9516 43004
rect 9516 42948 9520 43004
rect 9456 42944 9520 42948
rect 19216 43004 19280 43008
rect 19216 42948 19220 43004
rect 19220 42948 19276 43004
rect 19276 42948 19280 43004
rect 19216 42944 19280 42948
rect 19296 43004 19360 43008
rect 19296 42948 19300 43004
rect 19300 42948 19356 43004
rect 19356 42948 19360 43004
rect 19296 42944 19360 42948
rect 19376 43004 19440 43008
rect 19376 42948 19380 43004
rect 19380 42948 19436 43004
rect 19436 42948 19440 43004
rect 19376 42944 19440 42948
rect 19456 43004 19520 43008
rect 19456 42948 19460 43004
rect 19460 42948 19516 43004
rect 19516 42948 19520 43004
rect 19456 42944 19520 42948
rect 29216 43004 29280 43008
rect 29216 42948 29220 43004
rect 29220 42948 29276 43004
rect 29276 42948 29280 43004
rect 29216 42944 29280 42948
rect 29296 43004 29360 43008
rect 29296 42948 29300 43004
rect 29300 42948 29356 43004
rect 29356 42948 29360 43004
rect 29296 42944 29360 42948
rect 29376 43004 29440 43008
rect 29376 42948 29380 43004
rect 29380 42948 29436 43004
rect 29436 42948 29440 43004
rect 29376 42944 29440 42948
rect 29456 43004 29520 43008
rect 29456 42948 29460 43004
rect 29460 42948 29516 43004
rect 29516 42948 29520 43004
rect 29456 42944 29520 42948
rect 39216 43004 39280 43008
rect 39216 42948 39220 43004
rect 39220 42948 39276 43004
rect 39276 42948 39280 43004
rect 39216 42944 39280 42948
rect 39296 43004 39360 43008
rect 39296 42948 39300 43004
rect 39300 42948 39356 43004
rect 39356 42948 39360 43004
rect 39296 42944 39360 42948
rect 39376 43004 39440 43008
rect 39376 42948 39380 43004
rect 39380 42948 39436 43004
rect 39436 42948 39440 43004
rect 39376 42944 39440 42948
rect 39456 43004 39520 43008
rect 39456 42948 39460 43004
rect 39460 42948 39516 43004
rect 39516 42948 39520 43004
rect 39456 42944 39520 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 14216 42460 14280 42464
rect 14216 42404 14220 42460
rect 14220 42404 14276 42460
rect 14276 42404 14280 42460
rect 14216 42400 14280 42404
rect 14296 42460 14360 42464
rect 14296 42404 14300 42460
rect 14300 42404 14356 42460
rect 14356 42404 14360 42460
rect 14296 42400 14360 42404
rect 14376 42460 14440 42464
rect 14376 42404 14380 42460
rect 14380 42404 14436 42460
rect 14436 42404 14440 42460
rect 14376 42400 14440 42404
rect 14456 42460 14520 42464
rect 14456 42404 14460 42460
rect 14460 42404 14516 42460
rect 14516 42404 14520 42460
rect 14456 42400 14520 42404
rect 24216 42460 24280 42464
rect 24216 42404 24220 42460
rect 24220 42404 24276 42460
rect 24276 42404 24280 42460
rect 24216 42400 24280 42404
rect 24296 42460 24360 42464
rect 24296 42404 24300 42460
rect 24300 42404 24356 42460
rect 24356 42404 24360 42460
rect 24296 42400 24360 42404
rect 24376 42460 24440 42464
rect 24376 42404 24380 42460
rect 24380 42404 24436 42460
rect 24436 42404 24440 42460
rect 24376 42400 24440 42404
rect 24456 42460 24520 42464
rect 24456 42404 24460 42460
rect 24460 42404 24516 42460
rect 24516 42404 24520 42460
rect 24456 42400 24520 42404
rect 34216 42460 34280 42464
rect 34216 42404 34220 42460
rect 34220 42404 34276 42460
rect 34276 42404 34280 42460
rect 34216 42400 34280 42404
rect 34296 42460 34360 42464
rect 34296 42404 34300 42460
rect 34300 42404 34356 42460
rect 34356 42404 34360 42460
rect 34296 42400 34360 42404
rect 34376 42460 34440 42464
rect 34376 42404 34380 42460
rect 34380 42404 34436 42460
rect 34436 42404 34440 42460
rect 34376 42400 34440 42404
rect 34456 42460 34520 42464
rect 34456 42404 34460 42460
rect 34460 42404 34516 42460
rect 34516 42404 34520 42460
rect 34456 42400 34520 42404
rect 44216 42460 44280 42464
rect 44216 42404 44220 42460
rect 44220 42404 44276 42460
rect 44276 42404 44280 42460
rect 44216 42400 44280 42404
rect 44296 42460 44360 42464
rect 44296 42404 44300 42460
rect 44300 42404 44356 42460
rect 44356 42404 44360 42460
rect 44296 42400 44360 42404
rect 44376 42460 44440 42464
rect 44376 42404 44380 42460
rect 44380 42404 44436 42460
rect 44436 42404 44440 42460
rect 44376 42400 44440 42404
rect 44456 42460 44520 42464
rect 44456 42404 44460 42460
rect 44460 42404 44516 42460
rect 44516 42404 44520 42460
rect 44456 42400 44520 42404
rect 9216 41916 9280 41920
rect 9216 41860 9220 41916
rect 9220 41860 9276 41916
rect 9276 41860 9280 41916
rect 9216 41856 9280 41860
rect 9296 41916 9360 41920
rect 9296 41860 9300 41916
rect 9300 41860 9356 41916
rect 9356 41860 9360 41916
rect 9296 41856 9360 41860
rect 9376 41916 9440 41920
rect 9376 41860 9380 41916
rect 9380 41860 9436 41916
rect 9436 41860 9440 41916
rect 9376 41856 9440 41860
rect 9456 41916 9520 41920
rect 9456 41860 9460 41916
rect 9460 41860 9516 41916
rect 9516 41860 9520 41916
rect 9456 41856 9520 41860
rect 19216 41916 19280 41920
rect 19216 41860 19220 41916
rect 19220 41860 19276 41916
rect 19276 41860 19280 41916
rect 19216 41856 19280 41860
rect 19296 41916 19360 41920
rect 19296 41860 19300 41916
rect 19300 41860 19356 41916
rect 19356 41860 19360 41916
rect 19296 41856 19360 41860
rect 19376 41916 19440 41920
rect 19376 41860 19380 41916
rect 19380 41860 19436 41916
rect 19436 41860 19440 41916
rect 19376 41856 19440 41860
rect 19456 41916 19520 41920
rect 19456 41860 19460 41916
rect 19460 41860 19516 41916
rect 19516 41860 19520 41916
rect 19456 41856 19520 41860
rect 29216 41916 29280 41920
rect 29216 41860 29220 41916
rect 29220 41860 29276 41916
rect 29276 41860 29280 41916
rect 29216 41856 29280 41860
rect 29296 41916 29360 41920
rect 29296 41860 29300 41916
rect 29300 41860 29356 41916
rect 29356 41860 29360 41916
rect 29296 41856 29360 41860
rect 29376 41916 29440 41920
rect 29376 41860 29380 41916
rect 29380 41860 29436 41916
rect 29436 41860 29440 41916
rect 29376 41856 29440 41860
rect 29456 41916 29520 41920
rect 29456 41860 29460 41916
rect 29460 41860 29516 41916
rect 29516 41860 29520 41916
rect 29456 41856 29520 41860
rect 39216 41916 39280 41920
rect 39216 41860 39220 41916
rect 39220 41860 39276 41916
rect 39276 41860 39280 41916
rect 39216 41856 39280 41860
rect 39296 41916 39360 41920
rect 39296 41860 39300 41916
rect 39300 41860 39356 41916
rect 39356 41860 39360 41916
rect 39296 41856 39360 41860
rect 39376 41916 39440 41920
rect 39376 41860 39380 41916
rect 39380 41860 39436 41916
rect 39436 41860 39440 41916
rect 39376 41856 39440 41860
rect 39456 41916 39520 41920
rect 39456 41860 39460 41916
rect 39460 41860 39516 41916
rect 39516 41860 39520 41916
rect 39456 41856 39520 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 14216 41372 14280 41376
rect 14216 41316 14220 41372
rect 14220 41316 14276 41372
rect 14276 41316 14280 41372
rect 14216 41312 14280 41316
rect 14296 41372 14360 41376
rect 14296 41316 14300 41372
rect 14300 41316 14356 41372
rect 14356 41316 14360 41372
rect 14296 41312 14360 41316
rect 14376 41372 14440 41376
rect 14376 41316 14380 41372
rect 14380 41316 14436 41372
rect 14436 41316 14440 41372
rect 14376 41312 14440 41316
rect 14456 41372 14520 41376
rect 14456 41316 14460 41372
rect 14460 41316 14516 41372
rect 14516 41316 14520 41372
rect 14456 41312 14520 41316
rect 24216 41372 24280 41376
rect 24216 41316 24220 41372
rect 24220 41316 24276 41372
rect 24276 41316 24280 41372
rect 24216 41312 24280 41316
rect 24296 41372 24360 41376
rect 24296 41316 24300 41372
rect 24300 41316 24356 41372
rect 24356 41316 24360 41372
rect 24296 41312 24360 41316
rect 24376 41372 24440 41376
rect 24376 41316 24380 41372
rect 24380 41316 24436 41372
rect 24436 41316 24440 41372
rect 24376 41312 24440 41316
rect 24456 41372 24520 41376
rect 24456 41316 24460 41372
rect 24460 41316 24516 41372
rect 24516 41316 24520 41372
rect 24456 41312 24520 41316
rect 34216 41372 34280 41376
rect 34216 41316 34220 41372
rect 34220 41316 34276 41372
rect 34276 41316 34280 41372
rect 34216 41312 34280 41316
rect 34296 41372 34360 41376
rect 34296 41316 34300 41372
rect 34300 41316 34356 41372
rect 34356 41316 34360 41372
rect 34296 41312 34360 41316
rect 34376 41372 34440 41376
rect 34376 41316 34380 41372
rect 34380 41316 34436 41372
rect 34436 41316 34440 41372
rect 34376 41312 34440 41316
rect 34456 41372 34520 41376
rect 34456 41316 34460 41372
rect 34460 41316 34516 41372
rect 34516 41316 34520 41372
rect 34456 41312 34520 41316
rect 44216 41372 44280 41376
rect 44216 41316 44220 41372
rect 44220 41316 44276 41372
rect 44276 41316 44280 41372
rect 44216 41312 44280 41316
rect 44296 41372 44360 41376
rect 44296 41316 44300 41372
rect 44300 41316 44356 41372
rect 44356 41316 44360 41372
rect 44296 41312 44360 41316
rect 44376 41372 44440 41376
rect 44376 41316 44380 41372
rect 44380 41316 44436 41372
rect 44436 41316 44440 41372
rect 44376 41312 44440 41316
rect 44456 41372 44520 41376
rect 44456 41316 44460 41372
rect 44460 41316 44516 41372
rect 44516 41316 44520 41372
rect 44456 41312 44520 41316
rect 9216 40828 9280 40832
rect 9216 40772 9220 40828
rect 9220 40772 9276 40828
rect 9276 40772 9280 40828
rect 9216 40768 9280 40772
rect 9296 40828 9360 40832
rect 9296 40772 9300 40828
rect 9300 40772 9356 40828
rect 9356 40772 9360 40828
rect 9296 40768 9360 40772
rect 9376 40828 9440 40832
rect 9376 40772 9380 40828
rect 9380 40772 9436 40828
rect 9436 40772 9440 40828
rect 9376 40768 9440 40772
rect 9456 40828 9520 40832
rect 9456 40772 9460 40828
rect 9460 40772 9516 40828
rect 9516 40772 9520 40828
rect 9456 40768 9520 40772
rect 19216 40828 19280 40832
rect 19216 40772 19220 40828
rect 19220 40772 19276 40828
rect 19276 40772 19280 40828
rect 19216 40768 19280 40772
rect 19296 40828 19360 40832
rect 19296 40772 19300 40828
rect 19300 40772 19356 40828
rect 19356 40772 19360 40828
rect 19296 40768 19360 40772
rect 19376 40828 19440 40832
rect 19376 40772 19380 40828
rect 19380 40772 19436 40828
rect 19436 40772 19440 40828
rect 19376 40768 19440 40772
rect 19456 40828 19520 40832
rect 19456 40772 19460 40828
rect 19460 40772 19516 40828
rect 19516 40772 19520 40828
rect 19456 40768 19520 40772
rect 29216 40828 29280 40832
rect 29216 40772 29220 40828
rect 29220 40772 29276 40828
rect 29276 40772 29280 40828
rect 29216 40768 29280 40772
rect 29296 40828 29360 40832
rect 29296 40772 29300 40828
rect 29300 40772 29356 40828
rect 29356 40772 29360 40828
rect 29296 40768 29360 40772
rect 29376 40828 29440 40832
rect 29376 40772 29380 40828
rect 29380 40772 29436 40828
rect 29436 40772 29440 40828
rect 29376 40768 29440 40772
rect 29456 40828 29520 40832
rect 29456 40772 29460 40828
rect 29460 40772 29516 40828
rect 29516 40772 29520 40828
rect 29456 40768 29520 40772
rect 39216 40828 39280 40832
rect 39216 40772 39220 40828
rect 39220 40772 39276 40828
rect 39276 40772 39280 40828
rect 39216 40768 39280 40772
rect 39296 40828 39360 40832
rect 39296 40772 39300 40828
rect 39300 40772 39356 40828
rect 39356 40772 39360 40828
rect 39296 40768 39360 40772
rect 39376 40828 39440 40832
rect 39376 40772 39380 40828
rect 39380 40772 39436 40828
rect 39436 40772 39440 40828
rect 39376 40768 39440 40772
rect 39456 40828 39520 40832
rect 39456 40772 39460 40828
rect 39460 40772 39516 40828
rect 39516 40772 39520 40828
rect 39456 40768 39520 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 14216 40284 14280 40288
rect 14216 40228 14220 40284
rect 14220 40228 14276 40284
rect 14276 40228 14280 40284
rect 14216 40224 14280 40228
rect 14296 40284 14360 40288
rect 14296 40228 14300 40284
rect 14300 40228 14356 40284
rect 14356 40228 14360 40284
rect 14296 40224 14360 40228
rect 14376 40284 14440 40288
rect 14376 40228 14380 40284
rect 14380 40228 14436 40284
rect 14436 40228 14440 40284
rect 14376 40224 14440 40228
rect 14456 40284 14520 40288
rect 14456 40228 14460 40284
rect 14460 40228 14516 40284
rect 14516 40228 14520 40284
rect 14456 40224 14520 40228
rect 24216 40284 24280 40288
rect 24216 40228 24220 40284
rect 24220 40228 24276 40284
rect 24276 40228 24280 40284
rect 24216 40224 24280 40228
rect 24296 40284 24360 40288
rect 24296 40228 24300 40284
rect 24300 40228 24356 40284
rect 24356 40228 24360 40284
rect 24296 40224 24360 40228
rect 24376 40284 24440 40288
rect 24376 40228 24380 40284
rect 24380 40228 24436 40284
rect 24436 40228 24440 40284
rect 24376 40224 24440 40228
rect 24456 40284 24520 40288
rect 24456 40228 24460 40284
rect 24460 40228 24516 40284
rect 24516 40228 24520 40284
rect 24456 40224 24520 40228
rect 34216 40284 34280 40288
rect 34216 40228 34220 40284
rect 34220 40228 34276 40284
rect 34276 40228 34280 40284
rect 34216 40224 34280 40228
rect 34296 40284 34360 40288
rect 34296 40228 34300 40284
rect 34300 40228 34356 40284
rect 34356 40228 34360 40284
rect 34296 40224 34360 40228
rect 34376 40284 34440 40288
rect 34376 40228 34380 40284
rect 34380 40228 34436 40284
rect 34436 40228 34440 40284
rect 34376 40224 34440 40228
rect 34456 40284 34520 40288
rect 34456 40228 34460 40284
rect 34460 40228 34516 40284
rect 34516 40228 34520 40284
rect 34456 40224 34520 40228
rect 44216 40284 44280 40288
rect 44216 40228 44220 40284
rect 44220 40228 44276 40284
rect 44276 40228 44280 40284
rect 44216 40224 44280 40228
rect 44296 40284 44360 40288
rect 44296 40228 44300 40284
rect 44300 40228 44356 40284
rect 44356 40228 44360 40284
rect 44296 40224 44360 40228
rect 44376 40284 44440 40288
rect 44376 40228 44380 40284
rect 44380 40228 44436 40284
rect 44436 40228 44440 40284
rect 44376 40224 44440 40228
rect 44456 40284 44520 40288
rect 44456 40228 44460 40284
rect 44460 40228 44516 40284
rect 44516 40228 44520 40284
rect 44456 40224 44520 40228
rect 9216 39740 9280 39744
rect 9216 39684 9220 39740
rect 9220 39684 9276 39740
rect 9276 39684 9280 39740
rect 9216 39680 9280 39684
rect 9296 39740 9360 39744
rect 9296 39684 9300 39740
rect 9300 39684 9356 39740
rect 9356 39684 9360 39740
rect 9296 39680 9360 39684
rect 9376 39740 9440 39744
rect 9376 39684 9380 39740
rect 9380 39684 9436 39740
rect 9436 39684 9440 39740
rect 9376 39680 9440 39684
rect 9456 39740 9520 39744
rect 9456 39684 9460 39740
rect 9460 39684 9516 39740
rect 9516 39684 9520 39740
rect 9456 39680 9520 39684
rect 19216 39740 19280 39744
rect 19216 39684 19220 39740
rect 19220 39684 19276 39740
rect 19276 39684 19280 39740
rect 19216 39680 19280 39684
rect 19296 39740 19360 39744
rect 19296 39684 19300 39740
rect 19300 39684 19356 39740
rect 19356 39684 19360 39740
rect 19296 39680 19360 39684
rect 19376 39740 19440 39744
rect 19376 39684 19380 39740
rect 19380 39684 19436 39740
rect 19436 39684 19440 39740
rect 19376 39680 19440 39684
rect 19456 39740 19520 39744
rect 19456 39684 19460 39740
rect 19460 39684 19516 39740
rect 19516 39684 19520 39740
rect 19456 39680 19520 39684
rect 29216 39740 29280 39744
rect 29216 39684 29220 39740
rect 29220 39684 29276 39740
rect 29276 39684 29280 39740
rect 29216 39680 29280 39684
rect 29296 39740 29360 39744
rect 29296 39684 29300 39740
rect 29300 39684 29356 39740
rect 29356 39684 29360 39740
rect 29296 39680 29360 39684
rect 29376 39740 29440 39744
rect 29376 39684 29380 39740
rect 29380 39684 29436 39740
rect 29436 39684 29440 39740
rect 29376 39680 29440 39684
rect 29456 39740 29520 39744
rect 29456 39684 29460 39740
rect 29460 39684 29516 39740
rect 29516 39684 29520 39740
rect 29456 39680 29520 39684
rect 39216 39740 39280 39744
rect 39216 39684 39220 39740
rect 39220 39684 39276 39740
rect 39276 39684 39280 39740
rect 39216 39680 39280 39684
rect 39296 39740 39360 39744
rect 39296 39684 39300 39740
rect 39300 39684 39356 39740
rect 39356 39684 39360 39740
rect 39296 39680 39360 39684
rect 39376 39740 39440 39744
rect 39376 39684 39380 39740
rect 39380 39684 39436 39740
rect 39436 39684 39440 39740
rect 39376 39680 39440 39684
rect 39456 39740 39520 39744
rect 39456 39684 39460 39740
rect 39460 39684 39516 39740
rect 39516 39684 39520 39740
rect 39456 39680 39520 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 14216 39196 14280 39200
rect 14216 39140 14220 39196
rect 14220 39140 14276 39196
rect 14276 39140 14280 39196
rect 14216 39136 14280 39140
rect 14296 39196 14360 39200
rect 14296 39140 14300 39196
rect 14300 39140 14356 39196
rect 14356 39140 14360 39196
rect 14296 39136 14360 39140
rect 14376 39196 14440 39200
rect 14376 39140 14380 39196
rect 14380 39140 14436 39196
rect 14436 39140 14440 39196
rect 14376 39136 14440 39140
rect 14456 39196 14520 39200
rect 14456 39140 14460 39196
rect 14460 39140 14516 39196
rect 14516 39140 14520 39196
rect 14456 39136 14520 39140
rect 24216 39196 24280 39200
rect 24216 39140 24220 39196
rect 24220 39140 24276 39196
rect 24276 39140 24280 39196
rect 24216 39136 24280 39140
rect 24296 39196 24360 39200
rect 24296 39140 24300 39196
rect 24300 39140 24356 39196
rect 24356 39140 24360 39196
rect 24296 39136 24360 39140
rect 24376 39196 24440 39200
rect 24376 39140 24380 39196
rect 24380 39140 24436 39196
rect 24436 39140 24440 39196
rect 24376 39136 24440 39140
rect 24456 39196 24520 39200
rect 24456 39140 24460 39196
rect 24460 39140 24516 39196
rect 24516 39140 24520 39196
rect 24456 39136 24520 39140
rect 34216 39196 34280 39200
rect 34216 39140 34220 39196
rect 34220 39140 34276 39196
rect 34276 39140 34280 39196
rect 34216 39136 34280 39140
rect 34296 39196 34360 39200
rect 34296 39140 34300 39196
rect 34300 39140 34356 39196
rect 34356 39140 34360 39196
rect 34296 39136 34360 39140
rect 34376 39196 34440 39200
rect 34376 39140 34380 39196
rect 34380 39140 34436 39196
rect 34436 39140 34440 39196
rect 34376 39136 34440 39140
rect 34456 39196 34520 39200
rect 34456 39140 34460 39196
rect 34460 39140 34516 39196
rect 34516 39140 34520 39196
rect 34456 39136 34520 39140
rect 44216 39196 44280 39200
rect 44216 39140 44220 39196
rect 44220 39140 44276 39196
rect 44276 39140 44280 39196
rect 44216 39136 44280 39140
rect 44296 39196 44360 39200
rect 44296 39140 44300 39196
rect 44300 39140 44356 39196
rect 44356 39140 44360 39196
rect 44296 39136 44360 39140
rect 44376 39196 44440 39200
rect 44376 39140 44380 39196
rect 44380 39140 44436 39196
rect 44436 39140 44440 39196
rect 44376 39136 44440 39140
rect 44456 39196 44520 39200
rect 44456 39140 44460 39196
rect 44460 39140 44516 39196
rect 44516 39140 44520 39196
rect 44456 39136 44520 39140
rect 9216 38652 9280 38656
rect 9216 38596 9220 38652
rect 9220 38596 9276 38652
rect 9276 38596 9280 38652
rect 9216 38592 9280 38596
rect 9296 38652 9360 38656
rect 9296 38596 9300 38652
rect 9300 38596 9356 38652
rect 9356 38596 9360 38652
rect 9296 38592 9360 38596
rect 9376 38652 9440 38656
rect 9376 38596 9380 38652
rect 9380 38596 9436 38652
rect 9436 38596 9440 38652
rect 9376 38592 9440 38596
rect 9456 38652 9520 38656
rect 9456 38596 9460 38652
rect 9460 38596 9516 38652
rect 9516 38596 9520 38652
rect 9456 38592 9520 38596
rect 19216 38652 19280 38656
rect 19216 38596 19220 38652
rect 19220 38596 19276 38652
rect 19276 38596 19280 38652
rect 19216 38592 19280 38596
rect 19296 38652 19360 38656
rect 19296 38596 19300 38652
rect 19300 38596 19356 38652
rect 19356 38596 19360 38652
rect 19296 38592 19360 38596
rect 19376 38652 19440 38656
rect 19376 38596 19380 38652
rect 19380 38596 19436 38652
rect 19436 38596 19440 38652
rect 19376 38592 19440 38596
rect 19456 38652 19520 38656
rect 19456 38596 19460 38652
rect 19460 38596 19516 38652
rect 19516 38596 19520 38652
rect 19456 38592 19520 38596
rect 29216 38652 29280 38656
rect 29216 38596 29220 38652
rect 29220 38596 29276 38652
rect 29276 38596 29280 38652
rect 29216 38592 29280 38596
rect 29296 38652 29360 38656
rect 29296 38596 29300 38652
rect 29300 38596 29356 38652
rect 29356 38596 29360 38652
rect 29296 38592 29360 38596
rect 29376 38652 29440 38656
rect 29376 38596 29380 38652
rect 29380 38596 29436 38652
rect 29436 38596 29440 38652
rect 29376 38592 29440 38596
rect 29456 38652 29520 38656
rect 29456 38596 29460 38652
rect 29460 38596 29516 38652
rect 29516 38596 29520 38652
rect 29456 38592 29520 38596
rect 39216 38652 39280 38656
rect 39216 38596 39220 38652
rect 39220 38596 39276 38652
rect 39276 38596 39280 38652
rect 39216 38592 39280 38596
rect 39296 38652 39360 38656
rect 39296 38596 39300 38652
rect 39300 38596 39356 38652
rect 39356 38596 39360 38652
rect 39296 38592 39360 38596
rect 39376 38652 39440 38656
rect 39376 38596 39380 38652
rect 39380 38596 39436 38652
rect 39436 38596 39440 38652
rect 39376 38592 39440 38596
rect 39456 38652 39520 38656
rect 39456 38596 39460 38652
rect 39460 38596 39516 38652
rect 39516 38596 39520 38652
rect 39456 38592 39520 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 14216 38108 14280 38112
rect 14216 38052 14220 38108
rect 14220 38052 14276 38108
rect 14276 38052 14280 38108
rect 14216 38048 14280 38052
rect 14296 38108 14360 38112
rect 14296 38052 14300 38108
rect 14300 38052 14356 38108
rect 14356 38052 14360 38108
rect 14296 38048 14360 38052
rect 14376 38108 14440 38112
rect 14376 38052 14380 38108
rect 14380 38052 14436 38108
rect 14436 38052 14440 38108
rect 14376 38048 14440 38052
rect 14456 38108 14520 38112
rect 14456 38052 14460 38108
rect 14460 38052 14516 38108
rect 14516 38052 14520 38108
rect 14456 38048 14520 38052
rect 24216 38108 24280 38112
rect 24216 38052 24220 38108
rect 24220 38052 24276 38108
rect 24276 38052 24280 38108
rect 24216 38048 24280 38052
rect 24296 38108 24360 38112
rect 24296 38052 24300 38108
rect 24300 38052 24356 38108
rect 24356 38052 24360 38108
rect 24296 38048 24360 38052
rect 24376 38108 24440 38112
rect 24376 38052 24380 38108
rect 24380 38052 24436 38108
rect 24436 38052 24440 38108
rect 24376 38048 24440 38052
rect 24456 38108 24520 38112
rect 24456 38052 24460 38108
rect 24460 38052 24516 38108
rect 24516 38052 24520 38108
rect 24456 38048 24520 38052
rect 34216 38108 34280 38112
rect 34216 38052 34220 38108
rect 34220 38052 34276 38108
rect 34276 38052 34280 38108
rect 34216 38048 34280 38052
rect 34296 38108 34360 38112
rect 34296 38052 34300 38108
rect 34300 38052 34356 38108
rect 34356 38052 34360 38108
rect 34296 38048 34360 38052
rect 34376 38108 34440 38112
rect 34376 38052 34380 38108
rect 34380 38052 34436 38108
rect 34436 38052 34440 38108
rect 34376 38048 34440 38052
rect 34456 38108 34520 38112
rect 34456 38052 34460 38108
rect 34460 38052 34516 38108
rect 34516 38052 34520 38108
rect 34456 38048 34520 38052
rect 44216 38108 44280 38112
rect 44216 38052 44220 38108
rect 44220 38052 44276 38108
rect 44276 38052 44280 38108
rect 44216 38048 44280 38052
rect 44296 38108 44360 38112
rect 44296 38052 44300 38108
rect 44300 38052 44356 38108
rect 44356 38052 44360 38108
rect 44296 38048 44360 38052
rect 44376 38108 44440 38112
rect 44376 38052 44380 38108
rect 44380 38052 44436 38108
rect 44436 38052 44440 38108
rect 44376 38048 44440 38052
rect 44456 38108 44520 38112
rect 44456 38052 44460 38108
rect 44460 38052 44516 38108
rect 44516 38052 44520 38108
rect 44456 38048 44520 38052
rect 9216 37564 9280 37568
rect 9216 37508 9220 37564
rect 9220 37508 9276 37564
rect 9276 37508 9280 37564
rect 9216 37504 9280 37508
rect 9296 37564 9360 37568
rect 9296 37508 9300 37564
rect 9300 37508 9356 37564
rect 9356 37508 9360 37564
rect 9296 37504 9360 37508
rect 9376 37564 9440 37568
rect 9376 37508 9380 37564
rect 9380 37508 9436 37564
rect 9436 37508 9440 37564
rect 9376 37504 9440 37508
rect 9456 37564 9520 37568
rect 9456 37508 9460 37564
rect 9460 37508 9516 37564
rect 9516 37508 9520 37564
rect 9456 37504 9520 37508
rect 19216 37564 19280 37568
rect 19216 37508 19220 37564
rect 19220 37508 19276 37564
rect 19276 37508 19280 37564
rect 19216 37504 19280 37508
rect 19296 37564 19360 37568
rect 19296 37508 19300 37564
rect 19300 37508 19356 37564
rect 19356 37508 19360 37564
rect 19296 37504 19360 37508
rect 19376 37564 19440 37568
rect 19376 37508 19380 37564
rect 19380 37508 19436 37564
rect 19436 37508 19440 37564
rect 19376 37504 19440 37508
rect 19456 37564 19520 37568
rect 19456 37508 19460 37564
rect 19460 37508 19516 37564
rect 19516 37508 19520 37564
rect 19456 37504 19520 37508
rect 29216 37564 29280 37568
rect 29216 37508 29220 37564
rect 29220 37508 29276 37564
rect 29276 37508 29280 37564
rect 29216 37504 29280 37508
rect 29296 37564 29360 37568
rect 29296 37508 29300 37564
rect 29300 37508 29356 37564
rect 29356 37508 29360 37564
rect 29296 37504 29360 37508
rect 29376 37564 29440 37568
rect 29376 37508 29380 37564
rect 29380 37508 29436 37564
rect 29436 37508 29440 37564
rect 29376 37504 29440 37508
rect 29456 37564 29520 37568
rect 29456 37508 29460 37564
rect 29460 37508 29516 37564
rect 29516 37508 29520 37564
rect 29456 37504 29520 37508
rect 39216 37564 39280 37568
rect 39216 37508 39220 37564
rect 39220 37508 39276 37564
rect 39276 37508 39280 37564
rect 39216 37504 39280 37508
rect 39296 37564 39360 37568
rect 39296 37508 39300 37564
rect 39300 37508 39356 37564
rect 39356 37508 39360 37564
rect 39296 37504 39360 37508
rect 39376 37564 39440 37568
rect 39376 37508 39380 37564
rect 39380 37508 39436 37564
rect 39436 37508 39440 37564
rect 39376 37504 39440 37508
rect 39456 37564 39520 37568
rect 39456 37508 39460 37564
rect 39460 37508 39516 37564
rect 39516 37508 39520 37564
rect 39456 37504 39520 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 14216 37020 14280 37024
rect 14216 36964 14220 37020
rect 14220 36964 14276 37020
rect 14276 36964 14280 37020
rect 14216 36960 14280 36964
rect 14296 37020 14360 37024
rect 14296 36964 14300 37020
rect 14300 36964 14356 37020
rect 14356 36964 14360 37020
rect 14296 36960 14360 36964
rect 14376 37020 14440 37024
rect 14376 36964 14380 37020
rect 14380 36964 14436 37020
rect 14436 36964 14440 37020
rect 14376 36960 14440 36964
rect 14456 37020 14520 37024
rect 14456 36964 14460 37020
rect 14460 36964 14516 37020
rect 14516 36964 14520 37020
rect 14456 36960 14520 36964
rect 24216 37020 24280 37024
rect 24216 36964 24220 37020
rect 24220 36964 24276 37020
rect 24276 36964 24280 37020
rect 24216 36960 24280 36964
rect 24296 37020 24360 37024
rect 24296 36964 24300 37020
rect 24300 36964 24356 37020
rect 24356 36964 24360 37020
rect 24296 36960 24360 36964
rect 24376 37020 24440 37024
rect 24376 36964 24380 37020
rect 24380 36964 24436 37020
rect 24436 36964 24440 37020
rect 24376 36960 24440 36964
rect 24456 37020 24520 37024
rect 24456 36964 24460 37020
rect 24460 36964 24516 37020
rect 24516 36964 24520 37020
rect 24456 36960 24520 36964
rect 34216 37020 34280 37024
rect 34216 36964 34220 37020
rect 34220 36964 34276 37020
rect 34276 36964 34280 37020
rect 34216 36960 34280 36964
rect 34296 37020 34360 37024
rect 34296 36964 34300 37020
rect 34300 36964 34356 37020
rect 34356 36964 34360 37020
rect 34296 36960 34360 36964
rect 34376 37020 34440 37024
rect 34376 36964 34380 37020
rect 34380 36964 34436 37020
rect 34436 36964 34440 37020
rect 34376 36960 34440 36964
rect 34456 37020 34520 37024
rect 34456 36964 34460 37020
rect 34460 36964 34516 37020
rect 34516 36964 34520 37020
rect 34456 36960 34520 36964
rect 44216 37020 44280 37024
rect 44216 36964 44220 37020
rect 44220 36964 44276 37020
rect 44276 36964 44280 37020
rect 44216 36960 44280 36964
rect 44296 37020 44360 37024
rect 44296 36964 44300 37020
rect 44300 36964 44356 37020
rect 44356 36964 44360 37020
rect 44296 36960 44360 36964
rect 44376 37020 44440 37024
rect 44376 36964 44380 37020
rect 44380 36964 44436 37020
rect 44436 36964 44440 37020
rect 44376 36960 44440 36964
rect 44456 37020 44520 37024
rect 44456 36964 44460 37020
rect 44460 36964 44516 37020
rect 44516 36964 44520 37020
rect 44456 36960 44520 36964
rect 9216 36476 9280 36480
rect 9216 36420 9220 36476
rect 9220 36420 9276 36476
rect 9276 36420 9280 36476
rect 9216 36416 9280 36420
rect 9296 36476 9360 36480
rect 9296 36420 9300 36476
rect 9300 36420 9356 36476
rect 9356 36420 9360 36476
rect 9296 36416 9360 36420
rect 9376 36476 9440 36480
rect 9376 36420 9380 36476
rect 9380 36420 9436 36476
rect 9436 36420 9440 36476
rect 9376 36416 9440 36420
rect 9456 36476 9520 36480
rect 9456 36420 9460 36476
rect 9460 36420 9516 36476
rect 9516 36420 9520 36476
rect 9456 36416 9520 36420
rect 19216 36476 19280 36480
rect 19216 36420 19220 36476
rect 19220 36420 19276 36476
rect 19276 36420 19280 36476
rect 19216 36416 19280 36420
rect 19296 36476 19360 36480
rect 19296 36420 19300 36476
rect 19300 36420 19356 36476
rect 19356 36420 19360 36476
rect 19296 36416 19360 36420
rect 19376 36476 19440 36480
rect 19376 36420 19380 36476
rect 19380 36420 19436 36476
rect 19436 36420 19440 36476
rect 19376 36416 19440 36420
rect 19456 36476 19520 36480
rect 19456 36420 19460 36476
rect 19460 36420 19516 36476
rect 19516 36420 19520 36476
rect 19456 36416 19520 36420
rect 29216 36476 29280 36480
rect 29216 36420 29220 36476
rect 29220 36420 29276 36476
rect 29276 36420 29280 36476
rect 29216 36416 29280 36420
rect 29296 36476 29360 36480
rect 29296 36420 29300 36476
rect 29300 36420 29356 36476
rect 29356 36420 29360 36476
rect 29296 36416 29360 36420
rect 29376 36476 29440 36480
rect 29376 36420 29380 36476
rect 29380 36420 29436 36476
rect 29436 36420 29440 36476
rect 29376 36416 29440 36420
rect 29456 36476 29520 36480
rect 29456 36420 29460 36476
rect 29460 36420 29516 36476
rect 29516 36420 29520 36476
rect 29456 36416 29520 36420
rect 39216 36476 39280 36480
rect 39216 36420 39220 36476
rect 39220 36420 39276 36476
rect 39276 36420 39280 36476
rect 39216 36416 39280 36420
rect 39296 36476 39360 36480
rect 39296 36420 39300 36476
rect 39300 36420 39356 36476
rect 39356 36420 39360 36476
rect 39296 36416 39360 36420
rect 39376 36476 39440 36480
rect 39376 36420 39380 36476
rect 39380 36420 39436 36476
rect 39436 36420 39440 36476
rect 39376 36416 39440 36420
rect 39456 36476 39520 36480
rect 39456 36420 39460 36476
rect 39460 36420 39516 36476
rect 39516 36420 39520 36476
rect 39456 36416 39520 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 14216 35932 14280 35936
rect 14216 35876 14220 35932
rect 14220 35876 14276 35932
rect 14276 35876 14280 35932
rect 14216 35872 14280 35876
rect 14296 35932 14360 35936
rect 14296 35876 14300 35932
rect 14300 35876 14356 35932
rect 14356 35876 14360 35932
rect 14296 35872 14360 35876
rect 14376 35932 14440 35936
rect 14376 35876 14380 35932
rect 14380 35876 14436 35932
rect 14436 35876 14440 35932
rect 14376 35872 14440 35876
rect 14456 35932 14520 35936
rect 14456 35876 14460 35932
rect 14460 35876 14516 35932
rect 14516 35876 14520 35932
rect 14456 35872 14520 35876
rect 24216 35932 24280 35936
rect 24216 35876 24220 35932
rect 24220 35876 24276 35932
rect 24276 35876 24280 35932
rect 24216 35872 24280 35876
rect 24296 35932 24360 35936
rect 24296 35876 24300 35932
rect 24300 35876 24356 35932
rect 24356 35876 24360 35932
rect 24296 35872 24360 35876
rect 24376 35932 24440 35936
rect 24376 35876 24380 35932
rect 24380 35876 24436 35932
rect 24436 35876 24440 35932
rect 24376 35872 24440 35876
rect 24456 35932 24520 35936
rect 24456 35876 24460 35932
rect 24460 35876 24516 35932
rect 24516 35876 24520 35932
rect 24456 35872 24520 35876
rect 34216 35932 34280 35936
rect 34216 35876 34220 35932
rect 34220 35876 34276 35932
rect 34276 35876 34280 35932
rect 34216 35872 34280 35876
rect 34296 35932 34360 35936
rect 34296 35876 34300 35932
rect 34300 35876 34356 35932
rect 34356 35876 34360 35932
rect 34296 35872 34360 35876
rect 34376 35932 34440 35936
rect 34376 35876 34380 35932
rect 34380 35876 34436 35932
rect 34436 35876 34440 35932
rect 34376 35872 34440 35876
rect 34456 35932 34520 35936
rect 34456 35876 34460 35932
rect 34460 35876 34516 35932
rect 34516 35876 34520 35932
rect 34456 35872 34520 35876
rect 44216 35932 44280 35936
rect 44216 35876 44220 35932
rect 44220 35876 44276 35932
rect 44276 35876 44280 35932
rect 44216 35872 44280 35876
rect 44296 35932 44360 35936
rect 44296 35876 44300 35932
rect 44300 35876 44356 35932
rect 44356 35876 44360 35932
rect 44296 35872 44360 35876
rect 44376 35932 44440 35936
rect 44376 35876 44380 35932
rect 44380 35876 44436 35932
rect 44436 35876 44440 35932
rect 44376 35872 44440 35876
rect 44456 35932 44520 35936
rect 44456 35876 44460 35932
rect 44460 35876 44516 35932
rect 44516 35876 44520 35932
rect 44456 35872 44520 35876
rect 9216 35388 9280 35392
rect 9216 35332 9220 35388
rect 9220 35332 9276 35388
rect 9276 35332 9280 35388
rect 9216 35328 9280 35332
rect 9296 35388 9360 35392
rect 9296 35332 9300 35388
rect 9300 35332 9356 35388
rect 9356 35332 9360 35388
rect 9296 35328 9360 35332
rect 9376 35388 9440 35392
rect 9376 35332 9380 35388
rect 9380 35332 9436 35388
rect 9436 35332 9440 35388
rect 9376 35328 9440 35332
rect 9456 35388 9520 35392
rect 9456 35332 9460 35388
rect 9460 35332 9516 35388
rect 9516 35332 9520 35388
rect 9456 35328 9520 35332
rect 19216 35388 19280 35392
rect 19216 35332 19220 35388
rect 19220 35332 19276 35388
rect 19276 35332 19280 35388
rect 19216 35328 19280 35332
rect 19296 35388 19360 35392
rect 19296 35332 19300 35388
rect 19300 35332 19356 35388
rect 19356 35332 19360 35388
rect 19296 35328 19360 35332
rect 19376 35388 19440 35392
rect 19376 35332 19380 35388
rect 19380 35332 19436 35388
rect 19436 35332 19440 35388
rect 19376 35328 19440 35332
rect 19456 35388 19520 35392
rect 19456 35332 19460 35388
rect 19460 35332 19516 35388
rect 19516 35332 19520 35388
rect 19456 35328 19520 35332
rect 29216 35388 29280 35392
rect 29216 35332 29220 35388
rect 29220 35332 29276 35388
rect 29276 35332 29280 35388
rect 29216 35328 29280 35332
rect 29296 35388 29360 35392
rect 29296 35332 29300 35388
rect 29300 35332 29356 35388
rect 29356 35332 29360 35388
rect 29296 35328 29360 35332
rect 29376 35388 29440 35392
rect 29376 35332 29380 35388
rect 29380 35332 29436 35388
rect 29436 35332 29440 35388
rect 29376 35328 29440 35332
rect 29456 35388 29520 35392
rect 29456 35332 29460 35388
rect 29460 35332 29516 35388
rect 29516 35332 29520 35388
rect 29456 35328 29520 35332
rect 39216 35388 39280 35392
rect 39216 35332 39220 35388
rect 39220 35332 39276 35388
rect 39276 35332 39280 35388
rect 39216 35328 39280 35332
rect 39296 35388 39360 35392
rect 39296 35332 39300 35388
rect 39300 35332 39356 35388
rect 39356 35332 39360 35388
rect 39296 35328 39360 35332
rect 39376 35388 39440 35392
rect 39376 35332 39380 35388
rect 39380 35332 39436 35388
rect 39436 35332 39440 35388
rect 39376 35328 39440 35332
rect 39456 35388 39520 35392
rect 39456 35332 39460 35388
rect 39460 35332 39516 35388
rect 39516 35332 39520 35388
rect 39456 35328 39520 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 14216 34844 14280 34848
rect 14216 34788 14220 34844
rect 14220 34788 14276 34844
rect 14276 34788 14280 34844
rect 14216 34784 14280 34788
rect 14296 34844 14360 34848
rect 14296 34788 14300 34844
rect 14300 34788 14356 34844
rect 14356 34788 14360 34844
rect 14296 34784 14360 34788
rect 14376 34844 14440 34848
rect 14376 34788 14380 34844
rect 14380 34788 14436 34844
rect 14436 34788 14440 34844
rect 14376 34784 14440 34788
rect 14456 34844 14520 34848
rect 14456 34788 14460 34844
rect 14460 34788 14516 34844
rect 14516 34788 14520 34844
rect 14456 34784 14520 34788
rect 24216 34844 24280 34848
rect 24216 34788 24220 34844
rect 24220 34788 24276 34844
rect 24276 34788 24280 34844
rect 24216 34784 24280 34788
rect 24296 34844 24360 34848
rect 24296 34788 24300 34844
rect 24300 34788 24356 34844
rect 24356 34788 24360 34844
rect 24296 34784 24360 34788
rect 24376 34844 24440 34848
rect 24376 34788 24380 34844
rect 24380 34788 24436 34844
rect 24436 34788 24440 34844
rect 24376 34784 24440 34788
rect 24456 34844 24520 34848
rect 24456 34788 24460 34844
rect 24460 34788 24516 34844
rect 24516 34788 24520 34844
rect 24456 34784 24520 34788
rect 34216 34844 34280 34848
rect 34216 34788 34220 34844
rect 34220 34788 34276 34844
rect 34276 34788 34280 34844
rect 34216 34784 34280 34788
rect 34296 34844 34360 34848
rect 34296 34788 34300 34844
rect 34300 34788 34356 34844
rect 34356 34788 34360 34844
rect 34296 34784 34360 34788
rect 34376 34844 34440 34848
rect 34376 34788 34380 34844
rect 34380 34788 34436 34844
rect 34436 34788 34440 34844
rect 34376 34784 34440 34788
rect 34456 34844 34520 34848
rect 34456 34788 34460 34844
rect 34460 34788 34516 34844
rect 34516 34788 34520 34844
rect 34456 34784 34520 34788
rect 44216 34844 44280 34848
rect 44216 34788 44220 34844
rect 44220 34788 44276 34844
rect 44276 34788 44280 34844
rect 44216 34784 44280 34788
rect 44296 34844 44360 34848
rect 44296 34788 44300 34844
rect 44300 34788 44356 34844
rect 44356 34788 44360 34844
rect 44296 34784 44360 34788
rect 44376 34844 44440 34848
rect 44376 34788 44380 34844
rect 44380 34788 44436 34844
rect 44436 34788 44440 34844
rect 44376 34784 44440 34788
rect 44456 34844 44520 34848
rect 44456 34788 44460 34844
rect 44460 34788 44516 34844
rect 44516 34788 44520 34844
rect 44456 34784 44520 34788
rect 9216 34300 9280 34304
rect 9216 34244 9220 34300
rect 9220 34244 9276 34300
rect 9276 34244 9280 34300
rect 9216 34240 9280 34244
rect 9296 34300 9360 34304
rect 9296 34244 9300 34300
rect 9300 34244 9356 34300
rect 9356 34244 9360 34300
rect 9296 34240 9360 34244
rect 9376 34300 9440 34304
rect 9376 34244 9380 34300
rect 9380 34244 9436 34300
rect 9436 34244 9440 34300
rect 9376 34240 9440 34244
rect 9456 34300 9520 34304
rect 9456 34244 9460 34300
rect 9460 34244 9516 34300
rect 9516 34244 9520 34300
rect 9456 34240 9520 34244
rect 19216 34300 19280 34304
rect 19216 34244 19220 34300
rect 19220 34244 19276 34300
rect 19276 34244 19280 34300
rect 19216 34240 19280 34244
rect 19296 34300 19360 34304
rect 19296 34244 19300 34300
rect 19300 34244 19356 34300
rect 19356 34244 19360 34300
rect 19296 34240 19360 34244
rect 19376 34300 19440 34304
rect 19376 34244 19380 34300
rect 19380 34244 19436 34300
rect 19436 34244 19440 34300
rect 19376 34240 19440 34244
rect 19456 34300 19520 34304
rect 19456 34244 19460 34300
rect 19460 34244 19516 34300
rect 19516 34244 19520 34300
rect 19456 34240 19520 34244
rect 29216 34300 29280 34304
rect 29216 34244 29220 34300
rect 29220 34244 29276 34300
rect 29276 34244 29280 34300
rect 29216 34240 29280 34244
rect 29296 34300 29360 34304
rect 29296 34244 29300 34300
rect 29300 34244 29356 34300
rect 29356 34244 29360 34300
rect 29296 34240 29360 34244
rect 29376 34300 29440 34304
rect 29376 34244 29380 34300
rect 29380 34244 29436 34300
rect 29436 34244 29440 34300
rect 29376 34240 29440 34244
rect 29456 34300 29520 34304
rect 29456 34244 29460 34300
rect 29460 34244 29516 34300
rect 29516 34244 29520 34300
rect 29456 34240 29520 34244
rect 39216 34300 39280 34304
rect 39216 34244 39220 34300
rect 39220 34244 39276 34300
rect 39276 34244 39280 34300
rect 39216 34240 39280 34244
rect 39296 34300 39360 34304
rect 39296 34244 39300 34300
rect 39300 34244 39356 34300
rect 39356 34244 39360 34300
rect 39296 34240 39360 34244
rect 39376 34300 39440 34304
rect 39376 34244 39380 34300
rect 39380 34244 39436 34300
rect 39436 34244 39440 34300
rect 39376 34240 39440 34244
rect 39456 34300 39520 34304
rect 39456 34244 39460 34300
rect 39460 34244 39516 34300
rect 39516 34244 39520 34300
rect 39456 34240 39520 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 14216 33756 14280 33760
rect 14216 33700 14220 33756
rect 14220 33700 14276 33756
rect 14276 33700 14280 33756
rect 14216 33696 14280 33700
rect 14296 33756 14360 33760
rect 14296 33700 14300 33756
rect 14300 33700 14356 33756
rect 14356 33700 14360 33756
rect 14296 33696 14360 33700
rect 14376 33756 14440 33760
rect 14376 33700 14380 33756
rect 14380 33700 14436 33756
rect 14436 33700 14440 33756
rect 14376 33696 14440 33700
rect 14456 33756 14520 33760
rect 14456 33700 14460 33756
rect 14460 33700 14516 33756
rect 14516 33700 14520 33756
rect 14456 33696 14520 33700
rect 24216 33756 24280 33760
rect 24216 33700 24220 33756
rect 24220 33700 24276 33756
rect 24276 33700 24280 33756
rect 24216 33696 24280 33700
rect 24296 33756 24360 33760
rect 24296 33700 24300 33756
rect 24300 33700 24356 33756
rect 24356 33700 24360 33756
rect 24296 33696 24360 33700
rect 24376 33756 24440 33760
rect 24376 33700 24380 33756
rect 24380 33700 24436 33756
rect 24436 33700 24440 33756
rect 24376 33696 24440 33700
rect 24456 33756 24520 33760
rect 24456 33700 24460 33756
rect 24460 33700 24516 33756
rect 24516 33700 24520 33756
rect 24456 33696 24520 33700
rect 34216 33756 34280 33760
rect 34216 33700 34220 33756
rect 34220 33700 34276 33756
rect 34276 33700 34280 33756
rect 34216 33696 34280 33700
rect 34296 33756 34360 33760
rect 34296 33700 34300 33756
rect 34300 33700 34356 33756
rect 34356 33700 34360 33756
rect 34296 33696 34360 33700
rect 34376 33756 34440 33760
rect 34376 33700 34380 33756
rect 34380 33700 34436 33756
rect 34436 33700 34440 33756
rect 34376 33696 34440 33700
rect 34456 33756 34520 33760
rect 34456 33700 34460 33756
rect 34460 33700 34516 33756
rect 34516 33700 34520 33756
rect 34456 33696 34520 33700
rect 44216 33756 44280 33760
rect 44216 33700 44220 33756
rect 44220 33700 44276 33756
rect 44276 33700 44280 33756
rect 44216 33696 44280 33700
rect 44296 33756 44360 33760
rect 44296 33700 44300 33756
rect 44300 33700 44356 33756
rect 44356 33700 44360 33756
rect 44296 33696 44360 33700
rect 44376 33756 44440 33760
rect 44376 33700 44380 33756
rect 44380 33700 44436 33756
rect 44436 33700 44440 33756
rect 44376 33696 44440 33700
rect 44456 33756 44520 33760
rect 44456 33700 44460 33756
rect 44460 33700 44516 33756
rect 44516 33700 44520 33756
rect 44456 33696 44520 33700
rect 9216 33212 9280 33216
rect 9216 33156 9220 33212
rect 9220 33156 9276 33212
rect 9276 33156 9280 33212
rect 9216 33152 9280 33156
rect 9296 33212 9360 33216
rect 9296 33156 9300 33212
rect 9300 33156 9356 33212
rect 9356 33156 9360 33212
rect 9296 33152 9360 33156
rect 9376 33212 9440 33216
rect 9376 33156 9380 33212
rect 9380 33156 9436 33212
rect 9436 33156 9440 33212
rect 9376 33152 9440 33156
rect 9456 33212 9520 33216
rect 9456 33156 9460 33212
rect 9460 33156 9516 33212
rect 9516 33156 9520 33212
rect 9456 33152 9520 33156
rect 19216 33212 19280 33216
rect 19216 33156 19220 33212
rect 19220 33156 19276 33212
rect 19276 33156 19280 33212
rect 19216 33152 19280 33156
rect 19296 33212 19360 33216
rect 19296 33156 19300 33212
rect 19300 33156 19356 33212
rect 19356 33156 19360 33212
rect 19296 33152 19360 33156
rect 19376 33212 19440 33216
rect 19376 33156 19380 33212
rect 19380 33156 19436 33212
rect 19436 33156 19440 33212
rect 19376 33152 19440 33156
rect 19456 33212 19520 33216
rect 19456 33156 19460 33212
rect 19460 33156 19516 33212
rect 19516 33156 19520 33212
rect 19456 33152 19520 33156
rect 29216 33212 29280 33216
rect 29216 33156 29220 33212
rect 29220 33156 29276 33212
rect 29276 33156 29280 33212
rect 29216 33152 29280 33156
rect 29296 33212 29360 33216
rect 29296 33156 29300 33212
rect 29300 33156 29356 33212
rect 29356 33156 29360 33212
rect 29296 33152 29360 33156
rect 29376 33212 29440 33216
rect 29376 33156 29380 33212
rect 29380 33156 29436 33212
rect 29436 33156 29440 33212
rect 29376 33152 29440 33156
rect 29456 33212 29520 33216
rect 29456 33156 29460 33212
rect 29460 33156 29516 33212
rect 29516 33156 29520 33212
rect 29456 33152 29520 33156
rect 39216 33212 39280 33216
rect 39216 33156 39220 33212
rect 39220 33156 39276 33212
rect 39276 33156 39280 33212
rect 39216 33152 39280 33156
rect 39296 33212 39360 33216
rect 39296 33156 39300 33212
rect 39300 33156 39356 33212
rect 39356 33156 39360 33212
rect 39296 33152 39360 33156
rect 39376 33212 39440 33216
rect 39376 33156 39380 33212
rect 39380 33156 39436 33212
rect 39436 33156 39440 33212
rect 39376 33152 39440 33156
rect 39456 33212 39520 33216
rect 39456 33156 39460 33212
rect 39460 33156 39516 33212
rect 39516 33156 39520 33212
rect 39456 33152 39520 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 14216 32668 14280 32672
rect 14216 32612 14220 32668
rect 14220 32612 14276 32668
rect 14276 32612 14280 32668
rect 14216 32608 14280 32612
rect 14296 32668 14360 32672
rect 14296 32612 14300 32668
rect 14300 32612 14356 32668
rect 14356 32612 14360 32668
rect 14296 32608 14360 32612
rect 14376 32668 14440 32672
rect 14376 32612 14380 32668
rect 14380 32612 14436 32668
rect 14436 32612 14440 32668
rect 14376 32608 14440 32612
rect 14456 32668 14520 32672
rect 14456 32612 14460 32668
rect 14460 32612 14516 32668
rect 14516 32612 14520 32668
rect 14456 32608 14520 32612
rect 24216 32668 24280 32672
rect 24216 32612 24220 32668
rect 24220 32612 24276 32668
rect 24276 32612 24280 32668
rect 24216 32608 24280 32612
rect 24296 32668 24360 32672
rect 24296 32612 24300 32668
rect 24300 32612 24356 32668
rect 24356 32612 24360 32668
rect 24296 32608 24360 32612
rect 24376 32668 24440 32672
rect 24376 32612 24380 32668
rect 24380 32612 24436 32668
rect 24436 32612 24440 32668
rect 24376 32608 24440 32612
rect 24456 32668 24520 32672
rect 24456 32612 24460 32668
rect 24460 32612 24516 32668
rect 24516 32612 24520 32668
rect 24456 32608 24520 32612
rect 34216 32668 34280 32672
rect 34216 32612 34220 32668
rect 34220 32612 34276 32668
rect 34276 32612 34280 32668
rect 34216 32608 34280 32612
rect 34296 32668 34360 32672
rect 34296 32612 34300 32668
rect 34300 32612 34356 32668
rect 34356 32612 34360 32668
rect 34296 32608 34360 32612
rect 34376 32668 34440 32672
rect 34376 32612 34380 32668
rect 34380 32612 34436 32668
rect 34436 32612 34440 32668
rect 34376 32608 34440 32612
rect 34456 32668 34520 32672
rect 34456 32612 34460 32668
rect 34460 32612 34516 32668
rect 34516 32612 34520 32668
rect 34456 32608 34520 32612
rect 44216 32668 44280 32672
rect 44216 32612 44220 32668
rect 44220 32612 44276 32668
rect 44276 32612 44280 32668
rect 44216 32608 44280 32612
rect 44296 32668 44360 32672
rect 44296 32612 44300 32668
rect 44300 32612 44356 32668
rect 44356 32612 44360 32668
rect 44296 32608 44360 32612
rect 44376 32668 44440 32672
rect 44376 32612 44380 32668
rect 44380 32612 44436 32668
rect 44436 32612 44440 32668
rect 44376 32608 44440 32612
rect 44456 32668 44520 32672
rect 44456 32612 44460 32668
rect 44460 32612 44516 32668
rect 44516 32612 44520 32668
rect 44456 32608 44520 32612
rect 9216 32124 9280 32128
rect 9216 32068 9220 32124
rect 9220 32068 9276 32124
rect 9276 32068 9280 32124
rect 9216 32064 9280 32068
rect 9296 32124 9360 32128
rect 9296 32068 9300 32124
rect 9300 32068 9356 32124
rect 9356 32068 9360 32124
rect 9296 32064 9360 32068
rect 9376 32124 9440 32128
rect 9376 32068 9380 32124
rect 9380 32068 9436 32124
rect 9436 32068 9440 32124
rect 9376 32064 9440 32068
rect 9456 32124 9520 32128
rect 9456 32068 9460 32124
rect 9460 32068 9516 32124
rect 9516 32068 9520 32124
rect 9456 32064 9520 32068
rect 19216 32124 19280 32128
rect 19216 32068 19220 32124
rect 19220 32068 19276 32124
rect 19276 32068 19280 32124
rect 19216 32064 19280 32068
rect 19296 32124 19360 32128
rect 19296 32068 19300 32124
rect 19300 32068 19356 32124
rect 19356 32068 19360 32124
rect 19296 32064 19360 32068
rect 19376 32124 19440 32128
rect 19376 32068 19380 32124
rect 19380 32068 19436 32124
rect 19436 32068 19440 32124
rect 19376 32064 19440 32068
rect 19456 32124 19520 32128
rect 19456 32068 19460 32124
rect 19460 32068 19516 32124
rect 19516 32068 19520 32124
rect 19456 32064 19520 32068
rect 29216 32124 29280 32128
rect 29216 32068 29220 32124
rect 29220 32068 29276 32124
rect 29276 32068 29280 32124
rect 29216 32064 29280 32068
rect 29296 32124 29360 32128
rect 29296 32068 29300 32124
rect 29300 32068 29356 32124
rect 29356 32068 29360 32124
rect 29296 32064 29360 32068
rect 29376 32124 29440 32128
rect 29376 32068 29380 32124
rect 29380 32068 29436 32124
rect 29436 32068 29440 32124
rect 29376 32064 29440 32068
rect 29456 32124 29520 32128
rect 29456 32068 29460 32124
rect 29460 32068 29516 32124
rect 29516 32068 29520 32124
rect 29456 32064 29520 32068
rect 39216 32124 39280 32128
rect 39216 32068 39220 32124
rect 39220 32068 39276 32124
rect 39276 32068 39280 32124
rect 39216 32064 39280 32068
rect 39296 32124 39360 32128
rect 39296 32068 39300 32124
rect 39300 32068 39356 32124
rect 39356 32068 39360 32124
rect 39296 32064 39360 32068
rect 39376 32124 39440 32128
rect 39376 32068 39380 32124
rect 39380 32068 39436 32124
rect 39436 32068 39440 32124
rect 39376 32064 39440 32068
rect 39456 32124 39520 32128
rect 39456 32068 39460 32124
rect 39460 32068 39516 32124
rect 39516 32068 39520 32124
rect 39456 32064 39520 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 14216 31580 14280 31584
rect 14216 31524 14220 31580
rect 14220 31524 14276 31580
rect 14276 31524 14280 31580
rect 14216 31520 14280 31524
rect 14296 31580 14360 31584
rect 14296 31524 14300 31580
rect 14300 31524 14356 31580
rect 14356 31524 14360 31580
rect 14296 31520 14360 31524
rect 14376 31580 14440 31584
rect 14376 31524 14380 31580
rect 14380 31524 14436 31580
rect 14436 31524 14440 31580
rect 14376 31520 14440 31524
rect 14456 31580 14520 31584
rect 14456 31524 14460 31580
rect 14460 31524 14516 31580
rect 14516 31524 14520 31580
rect 14456 31520 14520 31524
rect 24216 31580 24280 31584
rect 24216 31524 24220 31580
rect 24220 31524 24276 31580
rect 24276 31524 24280 31580
rect 24216 31520 24280 31524
rect 24296 31580 24360 31584
rect 24296 31524 24300 31580
rect 24300 31524 24356 31580
rect 24356 31524 24360 31580
rect 24296 31520 24360 31524
rect 24376 31580 24440 31584
rect 24376 31524 24380 31580
rect 24380 31524 24436 31580
rect 24436 31524 24440 31580
rect 24376 31520 24440 31524
rect 24456 31580 24520 31584
rect 24456 31524 24460 31580
rect 24460 31524 24516 31580
rect 24516 31524 24520 31580
rect 24456 31520 24520 31524
rect 34216 31580 34280 31584
rect 34216 31524 34220 31580
rect 34220 31524 34276 31580
rect 34276 31524 34280 31580
rect 34216 31520 34280 31524
rect 34296 31580 34360 31584
rect 34296 31524 34300 31580
rect 34300 31524 34356 31580
rect 34356 31524 34360 31580
rect 34296 31520 34360 31524
rect 34376 31580 34440 31584
rect 34376 31524 34380 31580
rect 34380 31524 34436 31580
rect 34436 31524 34440 31580
rect 34376 31520 34440 31524
rect 34456 31580 34520 31584
rect 34456 31524 34460 31580
rect 34460 31524 34516 31580
rect 34516 31524 34520 31580
rect 34456 31520 34520 31524
rect 44216 31580 44280 31584
rect 44216 31524 44220 31580
rect 44220 31524 44276 31580
rect 44276 31524 44280 31580
rect 44216 31520 44280 31524
rect 44296 31580 44360 31584
rect 44296 31524 44300 31580
rect 44300 31524 44356 31580
rect 44356 31524 44360 31580
rect 44296 31520 44360 31524
rect 44376 31580 44440 31584
rect 44376 31524 44380 31580
rect 44380 31524 44436 31580
rect 44436 31524 44440 31580
rect 44376 31520 44440 31524
rect 44456 31580 44520 31584
rect 44456 31524 44460 31580
rect 44460 31524 44516 31580
rect 44516 31524 44520 31580
rect 44456 31520 44520 31524
rect 9216 31036 9280 31040
rect 9216 30980 9220 31036
rect 9220 30980 9276 31036
rect 9276 30980 9280 31036
rect 9216 30976 9280 30980
rect 9296 31036 9360 31040
rect 9296 30980 9300 31036
rect 9300 30980 9356 31036
rect 9356 30980 9360 31036
rect 9296 30976 9360 30980
rect 9376 31036 9440 31040
rect 9376 30980 9380 31036
rect 9380 30980 9436 31036
rect 9436 30980 9440 31036
rect 9376 30976 9440 30980
rect 9456 31036 9520 31040
rect 9456 30980 9460 31036
rect 9460 30980 9516 31036
rect 9516 30980 9520 31036
rect 9456 30976 9520 30980
rect 19216 31036 19280 31040
rect 19216 30980 19220 31036
rect 19220 30980 19276 31036
rect 19276 30980 19280 31036
rect 19216 30976 19280 30980
rect 19296 31036 19360 31040
rect 19296 30980 19300 31036
rect 19300 30980 19356 31036
rect 19356 30980 19360 31036
rect 19296 30976 19360 30980
rect 19376 31036 19440 31040
rect 19376 30980 19380 31036
rect 19380 30980 19436 31036
rect 19436 30980 19440 31036
rect 19376 30976 19440 30980
rect 19456 31036 19520 31040
rect 19456 30980 19460 31036
rect 19460 30980 19516 31036
rect 19516 30980 19520 31036
rect 19456 30976 19520 30980
rect 29216 31036 29280 31040
rect 29216 30980 29220 31036
rect 29220 30980 29276 31036
rect 29276 30980 29280 31036
rect 29216 30976 29280 30980
rect 29296 31036 29360 31040
rect 29296 30980 29300 31036
rect 29300 30980 29356 31036
rect 29356 30980 29360 31036
rect 29296 30976 29360 30980
rect 29376 31036 29440 31040
rect 29376 30980 29380 31036
rect 29380 30980 29436 31036
rect 29436 30980 29440 31036
rect 29376 30976 29440 30980
rect 29456 31036 29520 31040
rect 29456 30980 29460 31036
rect 29460 30980 29516 31036
rect 29516 30980 29520 31036
rect 29456 30976 29520 30980
rect 39216 31036 39280 31040
rect 39216 30980 39220 31036
rect 39220 30980 39276 31036
rect 39276 30980 39280 31036
rect 39216 30976 39280 30980
rect 39296 31036 39360 31040
rect 39296 30980 39300 31036
rect 39300 30980 39356 31036
rect 39356 30980 39360 31036
rect 39296 30976 39360 30980
rect 39376 31036 39440 31040
rect 39376 30980 39380 31036
rect 39380 30980 39436 31036
rect 39436 30980 39440 31036
rect 39376 30976 39440 30980
rect 39456 31036 39520 31040
rect 39456 30980 39460 31036
rect 39460 30980 39516 31036
rect 39516 30980 39520 31036
rect 39456 30976 39520 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 14216 30492 14280 30496
rect 14216 30436 14220 30492
rect 14220 30436 14276 30492
rect 14276 30436 14280 30492
rect 14216 30432 14280 30436
rect 14296 30492 14360 30496
rect 14296 30436 14300 30492
rect 14300 30436 14356 30492
rect 14356 30436 14360 30492
rect 14296 30432 14360 30436
rect 14376 30492 14440 30496
rect 14376 30436 14380 30492
rect 14380 30436 14436 30492
rect 14436 30436 14440 30492
rect 14376 30432 14440 30436
rect 14456 30492 14520 30496
rect 14456 30436 14460 30492
rect 14460 30436 14516 30492
rect 14516 30436 14520 30492
rect 14456 30432 14520 30436
rect 24216 30492 24280 30496
rect 24216 30436 24220 30492
rect 24220 30436 24276 30492
rect 24276 30436 24280 30492
rect 24216 30432 24280 30436
rect 24296 30492 24360 30496
rect 24296 30436 24300 30492
rect 24300 30436 24356 30492
rect 24356 30436 24360 30492
rect 24296 30432 24360 30436
rect 24376 30492 24440 30496
rect 24376 30436 24380 30492
rect 24380 30436 24436 30492
rect 24436 30436 24440 30492
rect 24376 30432 24440 30436
rect 24456 30492 24520 30496
rect 24456 30436 24460 30492
rect 24460 30436 24516 30492
rect 24516 30436 24520 30492
rect 24456 30432 24520 30436
rect 34216 30492 34280 30496
rect 34216 30436 34220 30492
rect 34220 30436 34276 30492
rect 34276 30436 34280 30492
rect 34216 30432 34280 30436
rect 34296 30492 34360 30496
rect 34296 30436 34300 30492
rect 34300 30436 34356 30492
rect 34356 30436 34360 30492
rect 34296 30432 34360 30436
rect 34376 30492 34440 30496
rect 34376 30436 34380 30492
rect 34380 30436 34436 30492
rect 34436 30436 34440 30492
rect 34376 30432 34440 30436
rect 34456 30492 34520 30496
rect 34456 30436 34460 30492
rect 34460 30436 34516 30492
rect 34516 30436 34520 30492
rect 34456 30432 34520 30436
rect 44216 30492 44280 30496
rect 44216 30436 44220 30492
rect 44220 30436 44276 30492
rect 44276 30436 44280 30492
rect 44216 30432 44280 30436
rect 44296 30492 44360 30496
rect 44296 30436 44300 30492
rect 44300 30436 44356 30492
rect 44356 30436 44360 30492
rect 44296 30432 44360 30436
rect 44376 30492 44440 30496
rect 44376 30436 44380 30492
rect 44380 30436 44436 30492
rect 44436 30436 44440 30492
rect 44376 30432 44440 30436
rect 44456 30492 44520 30496
rect 44456 30436 44460 30492
rect 44460 30436 44516 30492
rect 44516 30436 44520 30492
rect 44456 30432 44520 30436
rect 9216 29948 9280 29952
rect 9216 29892 9220 29948
rect 9220 29892 9276 29948
rect 9276 29892 9280 29948
rect 9216 29888 9280 29892
rect 9296 29948 9360 29952
rect 9296 29892 9300 29948
rect 9300 29892 9356 29948
rect 9356 29892 9360 29948
rect 9296 29888 9360 29892
rect 9376 29948 9440 29952
rect 9376 29892 9380 29948
rect 9380 29892 9436 29948
rect 9436 29892 9440 29948
rect 9376 29888 9440 29892
rect 9456 29948 9520 29952
rect 9456 29892 9460 29948
rect 9460 29892 9516 29948
rect 9516 29892 9520 29948
rect 9456 29888 9520 29892
rect 19216 29948 19280 29952
rect 19216 29892 19220 29948
rect 19220 29892 19276 29948
rect 19276 29892 19280 29948
rect 19216 29888 19280 29892
rect 19296 29948 19360 29952
rect 19296 29892 19300 29948
rect 19300 29892 19356 29948
rect 19356 29892 19360 29948
rect 19296 29888 19360 29892
rect 19376 29948 19440 29952
rect 19376 29892 19380 29948
rect 19380 29892 19436 29948
rect 19436 29892 19440 29948
rect 19376 29888 19440 29892
rect 19456 29948 19520 29952
rect 19456 29892 19460 29948
rect 19460 29892 19516 29948
rect 19516 29892 19520 29948
rect 19456 29888 19520 29892
rect 29216 29948 29280 29952
rect 29216 29892 29220 29948
rect 29220 29892 29276 29948
rect 29276 29892 29280 29948
rect 29216 29888 29280 29892
rect 29296 29948 29360 29952
rect 29296 29892 29300 29948
rect 29300 29892 29356 29948
rect 29356 29892 29360 29948
rect 29296 29888 29360 29892
rect 29376 29948 29440 29952
rect 29376 29892 29380 29948
rect 29380 29892 29436 29948
rect 29436 29892 29440 29948
rect 29376 29888 29440 29892
rect 29456 29948 29520 29952
rect 29456 29892 29460 29948
rect 29460 29892 29516 29948
rect 29516 29892 29520 29948
rect 29456 29888 29520 29892
rect 39216 29948 39280 29952
rect 39216 29892 39220 29948
rect 39220 29892 39276 29948
rect 39276 29892 39280 29948
rect 39216 29888 39280 29892
rect 39296 29948 39360 29952
rect 39296 29892 39300 29948
rect 39300 29892 39356 29948
rect 39356 29892 39360 29948
rect 39296 29888 39360 29892
rect 39376 29948 39440 29952
rect 39376 29892 39380 29948
rect 39380 29892 39436 29948
rect 39436 29892 39440 29948
rect 39376 29888 39440 29892
rect 39456 29948 39520 29952
rect 39456 29892 39460 29948
rect 39460 29892 39516 29948
rect 39516 29892 39520 29948
rect 39456 29888 39520 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 14216 29404 14280 29408
rect 14216 29348 14220 29404
rect 14220 29348 14276 29404
rect 14276 29348 14280 29404
rect 14216 29344 14280 29348
rect 14296 29404 14360 29408
rect 14296 29348 14300 29404
rect 14300 29348 14356 29404
rect 14356 29348 14360 29404
rect 14296 29344 14360 29348
rect 14376 29404 14440 29408
rect 14376 29348 14380 29404
rect 14380 29348 14436 29404
rect 14436 29348 14440 29404
rect 14376 29344 14440 29348
rect 14456 29404 14520 29408
rect 14456 29348 14460 29404
rect 14460 29348 14516 29404
rect 14516 29348 14520 29404
rect 14456 29344 14520 29348
rect 24216 29404 24280 29408
rect 24216 29348 24220 29404
rect 24220 29348 24276 29404
rect 24276 29348 24280 29404
rect 24216 29344 24280 29348
rect 24296 29404 24360 29408
rect 24296 29348 24300 29404
rect 24300 29348 24356 29404
rect 24356 29348 24360 29404
rect 24296 29344 24360 29348
rect 24376 29404 24440 29408
rect 24376 29348 24380 29404
rect 24380 29348 24436 29404
rect 24436 29348 24440 29404
rect 24376 29344 24440 29348
rect 24456 29404 24520 29408
rect 24456 29348 24460 29404
rect 24460 29348 24516 29404
rect 24516 29348 24520 29404
rect 24456 29344 24520 29348
rect 34216 29404 34280 29408
rect 34216 29348 34220 29404
rect 34220 29348 34276 29404
rect 34276 29348 34280 29404
rect 34216 29344 34280 29348
rect 34296 29404 34360 29408
rect 34296 29348 34300 29404
rect 34300 29348 34356 29404
rect 34356 29348 34360 29404
rect 34296 29344 34360 29348
rect 34376 29404 34440 29408
rect 34376 29348 34380 29404
rect 34380 29348 34436 29404
rect 34436 29348 34440 29404
rect 34376 29344 34440 29348
rect 34456 29404 34520 29408
rect 34456 29348 34460 29404
rect 34460 29348 34516 29404
rect 34516 29348 34520 29404
rect 34456 29344 34520 29348
rect 44216 29404 44280 29408
rect 44216 29348 44220 29404
rect 44220 29348 44276 29404
rect 44276 29348 44280 29404
rect 44216 29344 44280 29348
rect 44296 29404 44360 29408
rect 44296 29348 44300 29404
rect 44300 29348 44356 29404
rect 44356 29348 44360 29404
rect 44296 29344 44360 29348
rect 44376 29404 44440 29408
rect 44376 29348 44380 29404
rect 44380 29348 44436 29404
rect 44436 29348 44440 29404
rect 44376 29344 44440 29348
rect 44456 29404 44520 29408
rect 44456 29348 44460 29404
rect 44460 29348 44516 29404
rect 44516 29348 44520 29404
rect 44456 29344 44520 29348
rect 9216 28860 9280 28864
rect 9216 28804 9220 28860
rect 9220 28804 9276 28860
rect 9276 28804 9280 28860
rect 9216 28800 9280 28804
rect 9296 28860 9360 28864
rect 9296 28804 9300 28860
rect 9300 28804 9356 28860
rect 9356 28804 9360 28860
rect 9296 28800 9360 28804
rect 9376 28860 9440 28864
rect 9376 28804 9380 28860
rect 9380 28804 9436 28860
rect 9436 28804 9440 28860
rect 9376 28800 9440 28804
rect 9456 28860 9520 28864
rect 9456 28804 9460 28860
rect 9460 28804 9516 28860
rect 9516 28804 9520 28860
rect 9456 28800 9520 28804
rect 19216 28860 19280 28864
rect 19216 28804 19220 28860
rect 19220 28804 19276 28860
rect 19276 28804 19280 28860
rect 19216 28800 19280 28804
rect 19296 28860 19360 28864
rect 19296 28804 19300 28860
rect 19300 28804 19356 28860
rect 19356 28804 19360 28860
rect 19296 28800 19360 28804
rect 19376 28860 19440 28864
rect 19376 28804 19380 28860
rect 19380 28804 19436 28860
rect 19436 28804 19440 28860
rect 19376 28800 19440 28804
rect 19456 28860 19520 28864
rect 19456 28804 19460 28860
rect 19460 28804 19516 28860
rect 19516 28804 19520 28860
rect 19456 28800 19520 28804
rect 29216 28860 29280 28864
rect 29216 28804 29220 28860
rect 29220 28804 29276 28860
rect 29276 28804 29280 28860
rect 29216 28800 29280 28804
rect 29296 28860 29360 28864
rect 29296 28804 29300 28860
rect 29300 28804 29356 28860
rect 29356 28804 29360 28860
rect 29296 28800 29360 28804
rect 29376 28860 29440 28864
rect 29376 28804 29380 28860
rect 29380 28804 29436 28860
rect 29436 28804 29440 28860
rect 29376 28800 29440 28804
rect 29456 28860 29520 28864
rect 29456 28804 29460 28860
rect 29460 28804 29516 28860
rect 29516 28804 29520 28860
rect 29456 28800 29520 28804
rect 39216 28860 39280 28864
rect 39216 28804 39220 28860
rect 39220 28804 39276 28860
rect 39276 28804 39280 28860
rect 39216 28800 39280 28804
rect 39296 28860 39360 28864
rect 39296 28804 39300 28860
rect 39300 28804 39356 28860
rect 39356 28804 39360 28860
rect 39296 28800 39360 28804
rect 39376 28860 39440 28864
rect 39376 28804 39380 28860
rect 39380 28804 39436 28860
rect 39436 28804 39440 28860
rect 39376 28800 39440 28804
rect 39456 28860 39520 28864
rect 39456 28804 39460 28860
rect 39460 28804 39516 28860
rect 39516 28804 39520 28860
rect 39456 28800 39520 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 14216 28316 14280 28320
rect 14216 28260 14220 28316
rect 14220 28260 14276 28316
rect 14276 28260 14280 28316
rect 14216 28256 14280 28260
rect 14296 28316 14360 28320
rect 14296 28260 14300 28316
rect 14300 28260 14356 28316
rect 14356 28260 14360 28316
rect 14296 28256 14360 28260
rect 14376 28316 14440 28320
rect 14376 28260 14380 28316
rect 14380 28260 14436 28316
rect 14436 28260 14440 28316
rect 14376 28256 14440 28260
rect 14456 28316 14520 28320
rect 14456 28260 14460 28316
rect 14460 28260 14516 28316
rect 14516 28260 14520 28316
rect 14456 28256 14520 28260
rect 24216 28316 24280 28320
rect 24216 28260 24220 28316
rect 24220 28260 24276 28316
rect 24276 28260 24280 28316
rect 24216 28256 24280 28260
rect 24296 28316 24360 28320
rect 24296 28260 24300 28316
rect 24300 28260 24356 28316
rect 24356 28260 24360 28316
rect 24296 28256 24360 28260
rect 24376 28316 24440 28320
rect 24376 28260 24380 28316
rect 24380 28260 24436 28316
rect 24436 28260 24440 28316
rect 24376 28256 24440 28260
rect 24456 28316 24520 28320
rect 24456 28260 24460 28316
rect 24460 28260 24516 28316
rect 24516 28260 24520 28316
rect 24456 28256 24520 28260
rect 34216 28316 34280 28320
rect 34216 28260 34220 28316
rect 34220 28260 34276 28316
rect 34276 28260 34280 28316
rect 34216 28256 34280 28260
rect 34296 28316 34360 28320
rect 34296 28260 34300 28316
rect 34300 28260 34356 28316
rect 34356 28260 34360 28316
rect 34296 28256 34360 28260
rect 34376 28316 34440 28320
rect 34376 28260 34380 28316
rect 34380 28260 34436 28316
rect 34436 28260 34440 28316
rect 34376 28256 34440 28260
rect 34456 28316 34520 28320
rect 34456 28260 34460 28316
rect 34460 28260 34516 28316
rect 34516 28260 34520 28316
rect 34456 28256 34520 28260
rect 44216 28316 44280 28320
rect 44216 28260 44220 28316
rect 44220 28260 44276 28316
rect 44276 28260 44280 28316
rect 44216 28256 44280 28260
rect 44296 28316 44360 28320
rect 44296 28260 44300 28316
rect 44300 28260 44356 28316
rect 44356 28260 44360 28316
rect 44296 28256 44360 28260
rect 44376 28316 44440 28320
rect 44376 28260 44380 28316
rect 44380 28260 44436 28316
rect 44436 28260 44440 28316
rect 44376 28256 44440 28260
rect 44456 28316 44520 28320
rect 44456 28260 44460 28316
rect 44460 28260 44516 28316
rect 44516 28260 44520 28316
rect 44456 28256 44520 28260
rect 9216 27772 9280 27776
rect 9216 27716 9220 27772
rect 9220 27716 9276 27772
rect 9276 27716 9280 27772
rect 9216 27712 9280 27716
rect 9296 27772 9360 27776
rect 9296 27716 9300 27772
rect 9300 27716 9356 27772
rect 9356 27716 9360 27772
rect 9296 27712 9360 27716
rect 9376 27772 9440 27776
rect 9376 27716 9380 27772
rect 9380 27716 9436 27772
rect 9436 27716 9440 27772
rect 9376 27712 9440 27716
rect 9456 27772 9520 27776
rect 9456 27716 9460 27772
rect 9460 27716 9516 27772
rect 9516 27716 9520 27772
rect 9456 27712 9520 27716
rect 19216 27772 19280 27776
rect 19216 27716 19220 27772
rect 19220 27716 19276 27772
rect 19276 27716 19280 27772
rect 19216 27712 19280 27716
rect 19296 27772 19360 27776
rect 19296 27716 19300 27772
rect 19300 27716 19356 27772
rect 19356 27716 19360 27772
rect 19296 27712 19360 27716
rect 19376 27772 19440 27776
rect 19376 27716 19380 27772
rect 19380 27716 19436 27772
rect 19436 27716 19440 27772
rect 19376 27712 19440 27716
rect 19456 27772 19520 27776
rect 19456 27716 19460 27772
rect 19460 27716 19516 27772
rect 19516 27716 19520 27772
rect 19456 27712 19520 27716
rect 29216 27772 29280 27776
rect 29216 27716 29220 27772
rect 29220 27716 29276 27772
rect 29276 27716 29280 27772
rect 29216 27712 29280 27716
rect 29296 27772 29360 27776
rect 29296 27716 29300 27772
rect 29300 27716 29356 27772
rect 29356 27716 29360 27772
rect 29296 27712 29360 27716
rect 29376 27772 29440 27776
rect 29376 27716 29380 27772
rect 29380 27716 29436 27772
rect 29436 27716 29440 27772
rect 29376 27712 29440 27716
rect 29456 27772 29520 27776
rect 29456 27716 29460 27772
rect 29460 27716 29516 27772
rect 29516 27716 29520 27772
rect 29456 27712 29520 27716
rect 39216 27772 39280 27776
rect 39216 27716 39220 27772
rect 39220 27716 39276 27772
rect 39276 27716 39280 27772
rect 39216 27712 39280 27716
rect 39296 27772 39360 27776
rect 39296 27716 39300 27772
rect 39300 27716 39356 27772
rect 39356 27716 39360 27772
rect 39296 27712 39360 27716
rect 39376 27772 39440 27776
rect 39376 27716 39380 27772
rect 39380 27716 39436 27772
rect 39436 27716 39440 27772
rect 39376 27712 39440 27716
rect 39456 27772 39520 27776
rect 39456 27716 39460 27772
rect 39460 27716 39516 27772
rect 39516 27716 39520 27772
rect 39456 27712 39520 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 14216 27228 14280 27232
rect 14216 27172 14220 27228
rect 14220 27172 14276 27228
rect 14276 27172 14280 27228
rect 14216 27168 14280 27172
rect 14296 27228 14360 27232
rect 14296 27172 14300 27228
rect 14300 27172 14356 27228
rect 14356 27172 14360 27228
rect 14296 27168 14360 27172
rect 14376 27228 14440 27232
rect 14376 27172 14380 27228
rect 14380 27172 14436 27228
rect 14436 27172 14440 27228
rect 14376 27168 14440 27172
rect 14456 27228 14520 27232
rect 14456 27172 14460 27228
rect 14460 27172 14516 27228
rect 14516 27172 14520 27228
rect 14456 27168 14520 27172
rect 24216 27228 24280 27232
rect 24216 27172 24220 27228
rect 24220 27172 24276 27228
rect 24276 27172 24280 27228
rect 24216 27168 24280 27172
rect 24296 27228 24360 27232
rect 24296 27172 24300 27228
rect 24300 27172 24356 27228
rect 24356 27172 24360 27228
rect 24296 27168 24360 27172
rect 24376 27228 24440 27232
rect 24376 27172 24380 27228
rect 24380 27172 24436 27228
rect 24436 27172 24440 27228
rect 24376 27168 24440 27172
rect 24456 27228 24520 27232
rect 24456 27172 24460 27228
rect 24460 27172 24516 27228
rect 24516 27172 24520 27228
rect 24456 27168 24520 27172
rect 34216 27228 34280 27232
rect 34216 27172 34220 27228
rect 34220 27172 34276 27228
rect 34276 27172 34280 27228
rect 34216 27168 34280 27172
rect 34296 27228 34360 27232
rect 34296 27172 34300 27228
rect 34300 27172 34356 27228
rect 34356 27172 34360 27228
rect 34296 27168 34360 27172
rect 34376 27228 34440 27232
rect 34376 27172 34380 27228
rect 34380 27172 34436 27228
rect 34436 27172 34440 27228
rect 34376 27168 34440 27172
rect 34456 27228 34520 27232
rect 34456 27172 34460 27228
rect 34460 27172 34516 27228
rect 34516 27172 34520 27228
rect 34456 27168 34520 27172
rect 44216 27228 44280 27232
rect 44216 27172 44220 27228
rect 44220 27172 44276 27228
rect 44276 27172 44280 27228
rect 44216 27168 44280 27172
rect 44296 27228 44360 27232
rect 44296 27172 44300 27228
rect 44300 27172 44356 27228
rect 44356 27172 44360 27228
rect 44296 27168 44360 27172
rect 44376 27228 44440 27232
rect 44376 27172 44380 27228
rect 44380 27172 44436 27228
rect 44436 27172 44440 27228
rect 44376 27168 44440 27172
rect 44456 27228 44520 27232
rect 44456 27172 44460 27228
rect 44460 27172 44516 27228
rect 44516 27172 44520 27228
rect 44456 27168 44520 27172
rect 9216 26684 9280 26688
rect 9216 26628 9220 26684
rect 9220 26628 9276 26684
rect 9276 26628 9280 26684
rect 9216 26624 9280 26628
rect 9296 26684 9360 26688
rect 9296 26628 9300 26684
rect 9300 26628 9356 26684
rect 9356 26628 9360 26684
rect 9296 26624 9360 26628
rect 9376 26684 9440 26688
rect 9376 26628 9380 26684
rect 9380 26628 9436 26684
rect 9436 26628 9440 26684
rect 9376 26624 9440 26628
rect 9456 26684 9520 26688
rect 9456 26628 9460 26684
rect 9460 26628 9516 26684
rect 9516 26628 9520 26684
rect 9456 26624 9520 26628
rect 19216 26684 19280 26688
rect 19216 26628 19220 26684
rect 19220 26628 19276 26684
rect 19276 26628 19280 26684
rect 19216 26624 19280 26628
rect 19296 26684 19360 26688
rect 19296 26628 19300 26684
rect 19300 26628 19356 26684
rect 19356 26628 19360 26684
rect 19296 26624 19360 26628
rect 19376 26684 19440 26688
rect 19376 26628 19380 26684
rect 19380 26628 19436 26684
rect 19436 26628 19440 26684
rect 19376 26624 19440 26628
rect 19456 26684 19520 26688
rect 19456 26628 19460 26684
rect 19460 26628 19516 26684
rect 19516 26628 19520 26684
rect 19456 26624 19520 26628
rect 29216 26684 29280 26688
rect 29216 26628 29220 26684
rect 29220 26628 29276 26684
rect 29276 26628 29280 26684
rect 29216 26624 29280 26628
rect 29296 26684 29360 26688
rect 29296 26628 29300 26684
rect 29300 26628 29356 26684
rect 29356 26628 29360 26684
rect 29296 26624 29360 26628
rect 29376 26684 29440 26688
rect 29376 26628 29380 26684
rect 29380 26628 29436 26684
rect 29436 26628 29440 26684
rect 29376 26624 29440 26628
rect 29456 26684 29520 26688
rect 29456 26628 29460 26684
rect 29460 26628 29516 26684
rect 29516 26628 29520 26684
rect 29456 26624 29520 26628
rect 39216 26684 39280 26688
rect 39216 26628 39220 26684
rect 39220 26628 39276 26684
rect 39276 26628 39280 26684
rect 39216 26624 39280 26628
rect 39296 26684 39360 26688
rect 39296 26628 39300 26684
rect 39300 26628 39356 26684
rect 39356 26628 39360 26684
rect 39296 26624 39360 26628
rect 39376 26684 39440 26688
rect 39376 26628 39380 26684
rect 39380 26628 39436 26684
rect 39436 26628 39440 26684
rect 39376 26624 39440 26628
rect 39456 26684 39520 26688
rect 39456 26628 39460 26684
rect 39460 26628 39516 26684
rect 39516 26628 39520 26684
rect 39456 26624 39520 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 14216 26140 14280 26144
rect 14216 26084 14220 26140
rect 14220 26084 14276 26140
rect 14276 26084 14280 26140
rect 14216 26080 14280 26084
rect 14296 26140 14360 26144
rect 14296 26084 14300 26140
rect 14300 26084 14356 26140
rect 14356 26084 14360 26140
rect 14296 26080 14360 26084
rect 14376 26140 14440 26144
rect 14376 26084 14380 26140
rect 14380 26084 14436 26140
rect 14436 26084 14440 26140
rect 14376 26080 14440 26084
rect 14456 26140 14520 26144
rect 14456 26084 14460 26140
rect 14460 26084 14516 26140
rect 14516 26084 14520 26140
rect 14456 26080 14520 26084
rect 24216 26140 24280 26144
rect 24216 26084 24220 26140
rect 24220 26084 24276 26140
rect 24276 26084 24280 26140
rect 24216 26080 24280 26084
rect 24296 26140 24360 26144
rect 24296 26084 24300 26140
rect 24300 26084 24356 26140
rect 24356 26084 24360 26140
rect 24296 26080 24360 26084
rect 24376 26140 24440 26144
rect 24376 26084 24380 26140
rect 24380 26084 24436 26140
rect 24436 26084 24440 26140
rect 24376 26080 24440 26084
rect 24456 26140 24520 26144
rect 24456 26084 24460 26140
rect 24460 26084 24516 26140
rect 24516 26084 24520 26140
rect 24456 26080 24520 26084
rect 34216 26140 34280 26144
rect 34216 26084 34220 26140
rect 34220 26084 34276 26140
rect 34276 26084 34280 26140
rect 34216 26080 34280 26084
rect 34296 26140 34360 26144
rect 34296 26084 34300 26140
rect 34300 26084 34356 26140
rect 34356 26084 34360 26140
rect 34296 26080 34360 26084
rect 34376 26140 34440 26144
rect 34376 26084 34380 26140
rect 34380 26084 34436 26140
rect 34436 26084 34440 26140
rect 34376 26080 34440 26084
rect 34456 26140 34520 26144
rect 34456 26084 34460 26140
rect 34460 26084 34516 26140
rect 34516 26084 34520 26140
rect 34456 26080 34520 26084
rect 44216 26140 44280 26144
rect 44216 26084 44220 26140
rect 44220 26084 44276 26140
rect 44276 26084 44280 26140
rect 44216 26080 44280 26084
rect 44296 26140 44360 26144
rect 44296 26084 44300 26140
rect 44300 26084 44356 26140
rect 44356 26084 44360 26140
rect 44296 26080 44360 26084
rect 44376 26140 44440 26144
rect 44376 26084 44380 26140
rect 44380 26084 44436 26140
rect 44436 26084 44440 26140
rect 44376 26080 44440 26084
rect 44456 26140 44520 26144
rect 44456 26084 44460 26140
rect 44460 26084 44516 26140
rect 44516 26084 44520 26140
rect 44456 26080 44520 26084
rect 9216 25596 9280 25600
rect 9216 25540 9220 25596
rect 9220 25540 9276 25596
rect 9276 25540 9280 25596
rect 9216 25536 9280 25540
rect 9296 25596 9360 25600
rect 9296 25540 9300 25596
rect 9300 25540 9356 25596
rect 9356 25540 9360 25596
rect 9296 25536 9360 25540
rect 9376 25596 9440 25600
rect 9376 25540 9380 25596
rect 9380 25540 9436 25596
rect 9436 25540 9440 25596
rect 9376 25536 9440 25540
rect 9456 25596 9520 25600
rect 9456 25540 9460 25596
rect 9460 25540 9516 25596
rect 9516 25540 9520 25596
rect 9456 25536 9520 25540
rect 19216 25596 19280 25600
rect 19216 25540 19220 25596
rect 19220 25540 19276 25596
rect 19276 25540 19280 25596
rect 19216 25536 19280 25540
rect 19296 25596 19360 25600
rect 19296 25540 19300 25596
rect 19300 25540 19356 25596
rect 19356 25540 19360 25596
rect 19296 25536 19360 25540
rect 19376 25596 19440 25600
rect 19376 25540 19380 25596
rect 19380 25540 19436 25596
rect 19436 25540 19440 25596
rect 19376 25536 19440 25540
rect 19456 25596 19520 25600
rect 19456 25540 19460 25596
rect 19460 25540 19516 25596
rect 19516 25540 19520 25596
rect 19456 25536 19520 25540
rect 29216 25596 29280 25600
rect 29216 25540 29220 25596
rect 29220 25540 29276 25596
rect 29276 25540 29280 25596
rect 29216 25536 29280 25540
rect 29296 25596 29360 25600
rect 29296 25540 29300 25596
rect 29300 25540 29356 25596
rect 29356 25540 29360 25596
rect 29296 25536 29360 25540
rect 29376 25596 29440 25600
rect 29376 25540 29380 25596
rect 29380 25540 29436 25596
rect 29436 25540 29440 25596
rect 29376 25536 29440 25540
rect 29456 25596 29520 25600
rect 29456 25540 29460 25596
rect 29460 25540 29516 25596
rect 29516 25540 29520 25596
rect 29456 25536 29520 25540
rect 39216 25596 39280 25600
rect 39216 25540 39220 25596
rect 39220 25540 39276 25596
rect 39276 25540 39280 25596
rect 39216 25536 39280 25540
rect 39296 25596 39360 25600
rect 39296 25540 39300 25596
rect 39300 25540 39356 25596
rect 39356 25540 39360 25596
rect 39296 25536 39360 25540
rect 39376 25596 39440 25600
rect 39376 25540 39380 25596
rect 39380 25540 39436 25596
rect 39436 25540 39440 25596
rect 39376 25536 39440 25540
rect 39456 25596 39520 25600
rect 39456 25540 39460 25596
rect 39460 25540 39516 25596
rect 39516 25540 39520 25596
rect 39456 25536 39520 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 14216 25052 14280 25056
rect 14216 24996 14220 25052
rect 14220 24996 14276 25052
rect 14276 24996 14280 25052
rect 14216 24992 14280 24996
rect 14296 25052 14360 25056
rect 14296 24996 14300 25052
rect 14300 24996 14356 25052
rect 14356 24996 14360 25052
rect 14296 24992 14360 24996
rect 14376 25052 14440 25056
rect 14376 24996 14380 25052
rect 14380 24996 14436 25052
rect 14436 24996 14440 25052
rect 14376 24992 14440 24996
rect 14456 25052 14520 25056
rect 14456 24996 14460 25052
rect 14460 24996 14516 25052
rect 14516 24996 14520 25052
rect 14456 24992 14520 24996
rect 24216 25052 24280 25056
rect 24216 24996 24220 25052
rect 24220 24996 24276 25052
rect 24276 24996 24280 25052
rect 24216 24992 24280 24996
rect 24296 25052 24360 25056
rect 24296 24996 24300 25052
rect 24300 24996 24356 25052
rect 24356 24996 24360 25052
rect 24296 24992 24360 24996
rect 24376 25052 24440 25056
rect 24376 24996 24380 25052
rect 24380 24996 24436 25052
rect 24436 24996 24440 25052
rect 24376 24992 24440 24996
rect 24456 25052 24520 25056
rect 24456 24996 24460 25052
rect 24460 24996 24516 25052
rect 24516 24996 24520 25052
rect 24456 24992 24520 24996
rect 34216 25052 34280 25056
rect 34216 24996 34220 25052
rect 34220 24996 34276 25052
rect 34276 24996 34280 25052
rect 34216 24992 34280 24996
rect 34296 25052 34360 25056
rect 34296 24996 34300 25052
rect 34300 24996 34356 25052
rect 34356 24996 34360 25052
rect 34296 24992 34360 24996
rect 34376 25052 34440 25056
rect 34376 24996 34380 25052
rect 34380 24996 34436 25052
rect 34436 24996 34440 25052
rect 34376 24992 34440 24996
rect 34456 25052 34520 25056
rect 34456 24996 34460 25052
rect 34460 24996 34516 25052
rect 34516 24996 34520 25052
rect 34456 24992 34520 24996
rect 44216 25052 44280 25056
rect 44216 24996 44220 25052
rect 44220 24996 44276 25052
rect 44276 24996 44280 25052
rect 44216 24992 44280 24996
rect 44296 25052 44360 25056
rect 44296 24996 44300 25052
rect 44300 24996 44356 25052
rect 44356 24996 44360 25052
rect 44296 24992 44360 24996
rect 44376 25052 44440 25056
rect 44376 24996 44380 25052
rect 44380 24996 44436 25052
rect 44436 24996 44440 25052
rect 44376 24992 44440 24996
rect 44456 25052 44520 25056
rect 44456 24996 44460 25052
rect 44460 24996 44516 25052
rect 44516 24996 44520 25052
rect 44456 24992 44520 24996
rect 9216 24508 9280 24512
rect 9216 24452 9220 24508
rect 9220 24452 9276 24508
rect 9276 24452 9280 24508
rect 9216 24448 9280 24452
rect 9296 24508 9360 24512
rect 9296 24452 9300 24508
rect 9300 24452 9356 24508
rect 9356 24452 9360 24508
rect 9296 24448 9360 24452
rect 9376 24508 9440 24512
rect 9376 24452 9380 24508
rect 9380 24452 9436 24508
rect 9436 24452 9440 24508
rect 9376 24448 9440 24452
rect 9456 24508 9520 24512
rect 9456 24452 9460 24508
rect 9460 24452 9516 24508
rect 9516 24452 9520 24508
rect 9456 24448 9520 24452
rect 19216 24508 19280 24512
rect 19216 24452 19220 24508
rect 19220 24452 19276 24508
rect 19276 24452 19280 24508
rect 19216 24448 19280 24452
rect 19296 24508 19360 24512
rect 19296 24452 19300 24508
rect 19300 24452 19356 24508
rect 19356 24452 19360 24508
rect 19296 24448 19360 24452
rect 19376 24508 19440 24512
rect 19376 24452 19380 24508
rect 19380 24452 19436 24508
rect 19436 24452 19440 24508
rect 19376 24448 19440 24452
rect 19456 24508 19520 24512
rect 19456 24452 19460 24508
rect 19460 24452 19516 24508
rect 19516 24452 19520 24508
rect 19456 24448 19520 24452
rect 29216 24508 29280 24512
rect 29216 24452 29220 24508
rect 29220 24452 29276 24508
rect 29276 24452 29280 24508
rect 29216 24448 29280 24452
rect 29296 24508 29360 24512
rect 29296 24452 29300 24508
rect 29300 24452 29356 24508
rect 29356 24452 29360 24508
rect 29296 24448 29360 24452
rect 29376 24508 29440 24512
rect 29376 24452 29380 24508
rect 29380 24452 29436 24508
rect 29436 24452 29440 24508
rect 29376 24448 29440 24452
rect 29456 24508 29520 24512
rect 29456 24452 29460 24508
rect 29460 24452 29516 24508
rect 29516 24452 29520 24508
rect 29456 24448 29520 24452
rect 39216 24508 39280 24512
rect 39216 24452 39220 24508
rect 39220 24452 39276 24508
rect 39276 24452 39280 24508
rect 39216 24448 39280 24452
rect 39296 24508 39360 24512
rect 39296 24452 39300 24508
rect 39300 24452 39356 24508
rect 39356 24452 39360 24508
rect 39296 24448 39360 24452
rect 39376 24508 39440 24512
rect 39376 24452 39380 24508
rect 39380 24452 39436 24508
rect 39436 24452 39440 24508
rect 39376 24448 39440 24452
rect 39456 24508 39520 24512
rect 39456 24452 39460 24508
rect 39460 24452 39516 24508
rect 39516 24452 39520 24508
rect 39456 24448 39520 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 14216 23964 14280 23968
rect 14216 23908 14220 23964
rect 14220 23908 14276 23964
rect 14276 23908 14280 23964
rect 14216 23904 14280 23908
rect 14296 23964 14360 23968
rect 14296 23908 14300 23964
rect 14300 23908 14356 23964
rect 14356 23908 14360 23964
rect 14296 23904 14360 23908
rect 14376 23964 14440 23968
rect 14376 23908 14380 23964
rect 14380 23908 14436 23964
rect 14436 23908 14440 23964
rect 14376 23904 14440 23908
rect 14456 23964 14520 23968
rect 14456 23908 14460 23964
rect 14460 23908 14516 23964
rect 14516 23908 14520 23964
rect 14456 23904 14520 23908
rect 24216 23964 24280 23968
rect 24216 23908 24220 23964
rect 24220 23908 24276 23964
rect 24276 23908 24280 23964
rect 24216 23904 24280 23908
rect 24296 23964 24360 23968
rect 24296 23908 24300 23964
rect 24300 23908 24356 23964
rect 24356 23908 24360 23964
rect 24296 23904 24360 23908
rect 24376 23964 24440 23968
rect 24376 23908 24380 23964
rect 24380 23908 24436 23964
rect 24436 23908 24440 23964
rect 24376 23904 24440 23908
rect 24456 23964 24520 23968
rect 24456 23908 24460 23964
rect 24460 23908 24516 23964
rect 24516 23908 24520 23964
rect 24456 23904 24520 23908
rect 34216 23964 34280 23968
rect 34216 23908 34220 23964
rect 34220 23908 34276 23964
rect 34276 23908 34280 23964
rect 34216 23904 34280 23908
rect 34296 23964 34360 23968
rect 34296 23908 34300 23964
rect 34300 23908 34356 23964
rect 34356 23908 34360 23964
rect 34296 23904 34360 23908
rect 34376 23964 34440 23968
rect 34376 23908 34380 23964
rect 34380 23908 34436 23964
rect 34436 23908 34440 23964
rect 34376 23904 34440 23908
rect 34456 23964 34520 23968
rect 34456 23908 34460 23964
rect 34460 23908 34516 23964
rect 34516 23908 34520 23964
rect 34456 23904 34520 23908
rect 44216 23964 44280 23968
rect 44216 23908 44220 23964
rect 44220 23908 44276 23964
rect 44276 23908 44280 23964
rect 44216 23904 44280 23908
rect 44296 23964 44360 23968
rect 44296 23908 44300 23964
rect 44300 23908 44356 23964
rect 44356 23908 44360 23964
rect 44296 23904 44360 23908
rect 44376 23964 44440 23968
rect 44376 23908 44380 23964
rect 44380 23908 44436 23964
rect 44436 23908 44440 23964
rect 44376 23904 44440 23908
rect 44456 23964 44520 23968
rect 44456 23908 44460 23964
rect 44460 23908 44516 23964
rect 44516 23908 44520 23964
rect 44456 23904 44520 23908
rect 9216 23420 9280 23424
rect 9216 23364 9220 23420
rect 9220 23364 9276 23420
rect 9276 23364 9280 23420
rect 9216 23360 9280 23364
rect 9296 23420 9360 23424
rect 9296 23364 9300 23420
rect 9300 23364 9356 23420
rect 9356 23364 9360 23420
rect 9296 23360 9360 23364
rect 9376 23420 9440 23424
rect 9376 23364 9380 23420
rect 9380 23364 9436 23420
rect 9436 23364 9440 23420
rect 9376 23360 9440 23364
rect 9456 23420 9520 23424
rect 9456 23364 9460 23420
rect 9460 23364 9516 23420
rect 9516 23364 9520 23420
rect 9456 23360 9520 23364
rect 19216 23420 19280 23424
rect 19216 23364 19220 23420
rect 19220 23364 19276 23420
rect 19276 23364 19280 23420
rect 19216 23360 19280 23364
rect 19296 23420 19360 23424
rect 19296 23364 19300 23420
rect 19300 23364 19356 23420
rect 19356 23364 19360 23420
rect 19296 23360 19360 23364
rect 19376 23420 19440 23424
rect 19376 23364 19380 23420
rect 19380 23364 19436 23420
rect 19436 23364 19440 23420
rect 19376 23360 19440 23364
rect 19456 23420 19520 23424
rect 19456 23364 19460 23420
rect 19460 23364 19516 23420
rect 19516 23364 19520 23420
rect 19456 23360 19520 23364
rect 29216 23420 29280 23424
rect 29216 23364 29220 23420
rect 29220 23364 29276 23420
rect 29276 23364 29280 23420
rect 29216 23360 29280 23364
rect 29296 23420 29360 23424
rect 29296 23364 29300 23420
rect 29300 23364 29356 23420
rect 29356 23364 29360 23420
rect 29296 23360 29360 23364
rect 29376 23420 29440 23424
rect 29376 23364 29380 23420
rect 29380 23364 29436 23420
rect 29436 23364 29440 23420
rect 29376 23360 29440 23364
rect 29456 23420 29520 23424
rect 29456 23364 29460 23420
rect 29460 23364 29516 23420
rect 29516 23364 29520 23420
rect 29456 23360 29520 23364
rect 39216 23420 39280 23424
rect 39216 23364 39220 23420
rect 39220 23364 39276 23420
rect 39276 23364 39280 23420
rect 39216 23360 39280 23364
rect 39296 23420 39360 23424
rect 39296 23364 39300 23420
rect 39300 23364 39356 23420
rect 39356 23364 39360 23420
rect 39296 23360 39360 23364
rect 39376 23420 39440 23424
rect 39376 23364 39380 23420
rect 39380 23364 39436 23420
rect 39436 23364 39440 23420
rect 39376 23360 39440 23364
rect 39456 23420 39520 23424
rect 39456 23364 39460 23420
rect 39460 23364 39516 23420
rect 39516 23364 39520 23420
rect 39456 23360 39520 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 14216 22876 14280 22880
rect 14216 22820 14220 22876
rect 14220 22820 14276 22876
rect 14276 22820 14280 22876
rect 14216 22816 14280 22820
rect 14296 22876 14360 22880
rect 14296 22820 14300 22876
rect 14300 22820 14356 22876
rect 14356 22820 14360 22876
rect 14296 22816 14360 22820
rect 14376 22876 14440 22880
rect 14376 22820 14380 22876
rect 14380 22820 14436 22876
rect 14436 22820 14440 22876
rect 14376 22816 14440 22820
rect 14456 22876 14520 22880
rect 14456 22820 14460 22876
rect 14460 22820 14516 22876
rect 14516 22820 14520 22876
rect 14456 22816 14520 22820
rect 24216 22876 24280 22880
rect 24216 22820 24220 22876
rect 24220 22820 24276 22876
rect 24276 22820 24280 22876
rect 24216 22816 24280 22820
rect 24296 22876 24360 22880
rect 24296 22820 24300 22876
rect 24300 22820 24356 22876
rect 24356 22820 24360 22876
rect 24296 22816 24360 22820
rect 24376 22876 24440 22880
rect 24376 22820 24380 22876
rect 24380 22820 24436 22876
rect 24436 22820 24440 22876
rect 24376 22816 24440 22820
rect 24456 22876 24520 22880
rect 24456 22820 24460 22876
rect 24460 22820 24516 22876
rect 24516 22820 24520 22876
rect 24456 22816 24520 22820
rect 34216 22876 34280 22880
rect 34216 22820 34220 22876
rect 34220 22820 34276 22876
rect 34276 22820 34280 22876
rect 34216 22816 34280 22820
rect 34296 22876 34360 22880
rect 34296 22820 34300 22876
rect 34300 22820 34356 22876
rect 34356 22820 34360 22876
rect 34296 22816 34360 22820
rect 34376 22876 34440 22880
rect 34376 22820 34380 22876
rect 34380 22820 34436 22876
rect 34436 22820 34440 22876
rect 34376 22816 34440 22820
rect 34456 22876 34520 22880
rect 34456 22820 34460 22876
rect 34460 22820 34516 22876
rect 34516 22820 34520 22876
rect 34456 22816 34520 22820
rect 44216 22876 44280 22880
rect 44216 22820 44220 22876
rect 44220 22820 44276 22876
rect 44276 22820 44280 22876
rect 44216 22816 44280 22820
rect 44296 22876 44360 22880
rect 44296 22820 44300 22876
rect 44300 22820 44356 22876
rect 44356 22820 44360 22876
rect 44296 22816 44360 22820
rect 44376 22876 44440 22880
rect 44376 22820 44380 22876
rect 44380 22820 44436 22876
rect 44436 22820 44440 22876
rect 44376 22816 44440 22820
rect 44456 22876 44520 22880
rect 44456 22820 44460 22876
rect 44460 22820 44516 22876
rect 44516 22820 44520 22876
rect 44456 22816 44520 22820
rect 9216 22332 9280 22336
rect 9216 22276 9220 22332
rect 9220 22276 9276 22332
rect 9276 22276 9280 22332
rect 9216 22272 9280 22276
rect 9296 22332 9360 22336
rect 9296 22276 9300 22332
rect 9300 22276 9356 22332
rect 9356 22276 9360 22332
rect 9296 22272 9360 22276
rect 9376 22332 9440 22336
rect 9376 22276 9380 22332
rect 9380 22276 9436 22332
rect 9436 22276 9440 22332
rect 9376 22272 9440 22276
rect 9456 22332 9520 22336
rect 9456 22276 9460 22332
rect 9460 22276 9516 22332
rect 9516 22276 9520 22332
rect 9456 22272 9520 22276
rect 19216 22332 19280 22336
rect 19216 22276 19220 22332
rect 19220 22276 19276 22332
rect 19276 22276 19280 22332
rect 19216 22272 19280 22276
rect 19296 22332 19360 22336
rect 19296 22276 19300 22332
rect 19300 22276 19356 22332
rect 19356 22276 19360 22332
rect 19296 22272 19360 22276
rect 19376 22332 19440 22336
rect 19376 22276 19380 22332
rect 19380 22276 19436 22332
rect 19436 22276 19440 22332
rect 19376 22272 19440 22276
rect 19456 22332 19520 22336
rect 19456 22276 19460 22332
rect 19460 22276 19516 22332
rect 19516 22276 19520 22332
rect 19456 22272 19520 22276
rect 29216 22332 29280 22336
rect 29216 22276 29220 22332
rect 29220 22276 29276 22332
rect 29276 22276 29280 22332
rect 29216 22272 29280 22276
rect 29296 22332 29360 22336
rect 29296 22276 29300 22332
rect 29300 22276 29356 22332
rect 29356 22276 29360 22332
rect 29296 22272 29360 22276
rect 29376 22332 29440 22336
rect 29376 22276 29380 22332
rect 29380 22276 29436 22332
rect 29436 22276 29440 22332
rect 29376 22272 29440 22276
rect 29456 22332 29520 22336
rect 29456 22276 29460 22332
rect 29460 22276 29516 22332
rect 29516 22276 29520 22332
rect 29456 22272 29520 22276
rect 39216 22332 39280 22336
rect 39216 22276 39220 22332
rect 39220 22276 39276 22332
rect 39276 22276 39280 22332
rect 39216 22272 39280 22276
rect 39296 22332 39360 22336
rect 39296 22276 39300 22332
rect 39300 22276 39356 22332
rect 39356 22276 39360 22332
rect 39296 22272 39360 22276
rect 39376 22332 39440 22336
rect 39376 22276 39380 22332
rect 39380 22276 39436 22332
rect 39436 22276 39440 22332
rect 39376 22272 39440 22276
rect 39456 22332 39520 22336
rect 39456 22276 39460 22332
rect 39460 22276 39516 22332
rect 39516 22276 39520 22332
rect 39456 22272 39520 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 14216 21788 14280 21792
rect 14216 21732 14220 21788
rect 14220 21732 14276 21788
rect 14276 21732 14280 21788
rect 14216 21728 14280 21732
rect 14296 21788 14360 21792
rect 14296 21732 14300 21788
rect 14300 21732 14356 21788
rect 14356 21732 14360 21788
rect 14296 21728 14360 21732
rect 14376 21788 14440 21792
rect 14376 21732 14380 21788
rect 14380 21732 14436 21788
rect 14436 21732 14440 21788
rect 14376 21728 14440 21732
rect 14456 21788 14520 21792
rect 14456 21732 14460 21788
rect 14460 21732 14516 21788
rect 14516 21732 14520 21788
rect 14456 21728 14520 21732
rect 24216 21788 24280 21792
rect 24216 21732 24220 21788
rect 24220 21732 24276 21788
rect 24276 21732 24280 21788
rect 24216 21728 24280 21732
rect 24296 21788 24360 21792
rect 24296 21732 24300 21788
rect 24300 21732 24356 21788
rect 24356 21732 24360 21788
rect 24296 21728 24360 21732
rect 24376 21788 24440 21792
rect 24376 21732 24380 21788
rect 24380 21732 24436 21788
rect 24436 21732 24440 21788
rect 24376 21728 24440 21732
rect 24456 21788 24520 21792
rect 24456 21732 24460 21788
rect 24460 21732 24516 21788
rect 24516 21732 24520 21788
rect 24456 21728 24520 21732
rect 34216 21788 34280 21792
rect 34216 21732 34220 21788
rect 34220 21732 34276 21788
rect 34276 21732 34280 21788
rect 34216 21728 34280 21732
rect 34296 21788 34360 21792
rect 34296 21732 34300 21788
rect 34300 21732 34356 21788
rect 34356 21732 34360 21788
rect 34296 21728 34360 21732
rect 34376 21788 34440 21792
rect 34376 21732 34380 21788
rect 34380 21732 34436 21788
rect 34436 21732 34440 21788
rect 34376 21728 34440 21732
rect 34456 21788 34520 21792
rect 34456 21732 34460 21788
rect 34460 21732 34516 21788
rect 34516 21732 34520 21788
rect 34456 21728 34520 21732
rect 44216 21788 44280 21792
rect 44216 21732 44220 21788
rect 44220 21732 44276 21788
rect 44276 21732 44280 21788
rect 44216 21728 44280 21732
rect 44296 21788 44360 21792
rect 44296 21732 44300 21788
rect 44300 21732 44356 21788
rect 44356 21732 44360 21788
rect 44296 21728 44360 21732
rect 44376 21788 44440 21792
rect 44376 21732 44380 21788
rect 44380 21732 44436 21788
rect 44436 21732 44440 21788
rect 44376 21728 44440 21732
rect 44456 21788 44520 21792
rect 44456 21732 44460 21788
rect 44460 21732 44516 21788
rect 44516 21732 44520 21788
rect 44456 21728 44520 21732
rect 9216 21244 9280 21248
rect 9216 21188 9220 21244
rect 9220 21188 9276 21244
rect 9276 21188 9280 21244
rect 9216 21184 9280 21188
rect 9296 21244 9360 21248
rect 9296 21188 9300 21244
rect 9300 21188 9356 21244
rect 9356 21188 9360 21244
rect 9296 21184 9360 21188
rect 9376 21244 9440 21248
rect 9376 21188 9380 21244
rect 9380 21188 9436 21244
rect 9436 21188 9440 21244
rect 9376 21184 9440 21188
rect 9456 21244 9520 21248
rect 9456 21188 9460 21244
rect 9460 21188 9516 21244
rect 9516 21188 9520 21244
rect 9456 21184 9520 21188
rect 19216 21244 19280 21248
rect 19216 21188 19220 21244
rect 19220 21188 19276 21244
rect 19276 21188 19280 21244
rect 19216 21184 19280 21188
rect 19296 21244 19360 21248
rect 19296 21188 19300 21244
rect 19300 21188 19356 21244
rect 19356 21188 19360 21244
rect 19296 21184 19360 21188
rect 19376 21244 19440 21248
rect 19376 21188 19380 21244
rect 19380 21188 19436 21244
rect 19436 21188 19440 21244
rect 19376 21184 19440 21188
rect 19456 21244 19520 21248
rect 19456 21188 19460 21244
rect 19460 21188 19516 21244
rect 19516 21188 19520 21244
rect 19456 21184 19520 21188
rect 29216 21244 29280 21248
rect 29216 21188 29220 21244
rect 29220 21188 29276 21244
rect 29276 21188 29280 21244
rect 29216 21184 29280 21188
rect 29296 21244 29360 21248
rect 29296 21188 29300 21244
rect 29300 21188 29356 21244
rect 29356 21188 29360 21244
rect 29296 21184 29360 21188
rect 29376 21244 29440 21248
rect 29376 21188 29380 21244
rect 29380 21188 29436 21244
rect 29436 21188 29440 21244
rect 29376 21184 29440 21188
rect 29456 21244 29520 21248
rect 29456 21188 29460 21244
rect 29460 21188 29516 21244
rect 29516 21188 29520 21244
rect 29456 21184 29520 21188
rect 39216 21244 39280 21248
rect 39216 21188 39220 21244
rect 39220 21188 39276 21244
rect 39276 21188 39280 21244
rect 39216 21184 39280 21188
rect 39296 21244 39360 21248
rect 39296 21188 39300 21244
rect 39300 21188 39356 21244
rect 39356 21188 39360 21244
rect 39296 21184 39360 21188
rect 39376 21244 39440 21248
rect 39376 21188 39380 21244
rect 39380 21188 39436 21244
rect 39436 21188 39440 21244
rect 39376 21184 39440 21188
rect 39456 21244 39520 21248
rect 39456 21188 39460 21244
rect 39460 21188 39516 21244
rect 39516 21188 39520 21244
rect 39456 21184 39520 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 14216 20700 14280 20704
rect 14216 20644 14220 20700
rect 14220 20644 14276 20700
rect 14276 20644 14280 20700
rect 14216 20640 14280 20644
rect 14296 20700 14360 20704
rect 14296 20644 14300 20700
rect 14300 20644 14356 20700
rect 14356 20644 14360 20700
rect 14296 20640 14360 20644
rect 14376 20700 14440 20704
rect 14376 20644 14380 20700
rect 14380 20644 14436 20700
rect 14436 20644 14440 20700
rect 14376 20640 14440 20644
rect 14456 20700 14520 20704
rect 14456 20644 14460 20700
rect 14460 20644 14516 20700
rect 14516 20644 14520 20700
rect 14456 20640 14520 20644
rect 24216 20700 24280 20704
rect 24216 20644 24220 20700
rect 24220 20644 24276 20700
rect 24276 20644 24280 20700
rect 24216 20640 24280 20644
rect 24296 20700 24360 20704
rect 24296 20644 24300 20700
rect 24300 20644 24356 20700
rect 24356 20644 24360 20700
rect 24296 20640 24360 20644
rect 24376 20700 24440 20704
rect 24376 20644 24380 20700
rect 24380 20644 24436 20700
rect 24436 20644 24440 20700
rect 24376 20640 24440 20644
rect 24456 20700 24520 20704
rect 24456 20644 24460 20700
rect 24460 20644 24516 20700
rect 24516 20644 24520 20700
rect 24456 20640 24520 20644
rect 34216 20700 34280 20704
rect 34216 20644 34220 20700
rect 34220 20644 34276 20700
rect 34276 20644 34280 20700
rect 34216 20640 34280 20644
rect 34296 20700 34360 20704
rect 34296 20644 34300 20700
rect 34300 20644 34356 20700
rect 34356 20644 34360 20700
rect 34296 20640 34360 20644
rect 34376 20700 34440 20704
rect 34376 20644 34380 20700
rect 34380 20644 34436 20700
rect 34436 20644 34440 20700
rect 34376 20640 34440 20644
rect 34456 20700 34520 20704
rect 34456 20644 34460 20700
rect 34460 20644 34516 20700
rect 34516 20644 34520 20700
rect 34456 20640 34520 20644
rect 44216 20700 44280 20704
rect 44216 20644 44220 20700
rect 44220 20644 44276 20700
rect 44276 20644 44280 20700
rect 44216 20640 44280 20644
rect 44296 20700 44360 20704
rect 44296 20644 44300 20700
rect 44300 20644 44356 20700
rect 44356 20644 44360 20700
rect 44296 20640 44360 20644
rect 44376 20700 44440 20704
rect 44376 20644 44380 20700
rect 44380 20644 44436 20700
rect 44436 20644 44440 20700
rect 44376 20640 44440 20644
rect 44456 20700 44520 20704
rect 44456 20644 44460 20700
rect 44460 20644 44516 20700
rect 44516 20644 44520 20700
rect 44456 20640 44520 20644
rect 9216 20156 9280 20160
rect 9216 20100 9220 20156
rect 9220 20100 9276 20156
rect 9276 20100 9280 20156
rect 9216 20096 9280 20100
rect 9296 20156 9360 20160
rect 9296 20100 9300 20156
rect 9300 20100 9356 20156
rect 9356 20100 9360 20156
rect 9296 20096 9360 20100
rect 9376 20156 9440 20160
rect 9376 20100 9380 20156
rect 9380 20100 9436 20156
rect 9436 20100 9440 20156
rect 9376 20096 9440 20100
rect 9456 20156 9520 20160
rect 9456 20100 9460 20156
rect 9460 20100 9516 20156
rect 9516 20100 9520 20156
rect 9456 20096 9520 20100
rect 19216 20156 19280 20160
rect 19216 20100 19220 20156
rect 19220 20100 19276 20156
rect 19276 20100 19280 20156
rect 19216 20096 19280 20100
rect 19296 20156 19360 20160
rect 19296 20100 19300 20156
rect 19300 20100 19356 20156
rect 19356 20100 19360 20156
rect 19296 20096 19360 20100
rect 19376 20156 19440 20160
rect 19376 20100 19380 20156
rect 19380 20100 19436 20156
rect 19436 20100 19440 20156
rect 19376 20096 19440 20100
rect 19456 20156 19520 20160
rect 19456 20100 19460 20156
rect 19460 20100 19516 20156
rect 19516 20100 19520 20156
rect 19456 20096 19520 20100
rect 29216 20156 29280 20160
rect 29216 20100 29220 20156
rect 29220 20100 29276 20156
rect 29276 20100 29280 20156
rect 29216 20096 29280 20100
rect 29296 20156 29360 20160
rect 29296 20100 29300 20156
rect 29300 20100 29356 20156
rect 29356 20100 29360 20156
rect 29296 20096 29360 20100
rect 29376 20156 29440 20160
rect 29376 20100 29380 20156
rect 29380 20100 29436 20156
rect 29436 20100 29440 20156
rect 29376 20096 29440 20100
rect 29456 20156 29520 20160
rect 29456 20100 29460 20156
rect 29460 20100 29516 20156
rect 29516 20100 29520 20156
rect 29456 20096 29520 20100
rect 39216 20156 39280 20160
rect 39216 20100 39220 20156
rect 39220 20100 39276 20156
rect 39276 20100 39280 20156
rect 39216 20096 39280 20100
rect 39296 20156 39360 20160
rect 39296 20100 39300 20156
rect 39300 20100 39356 20156
rect 39356 20100 39360 20156
rect 39296 20096 39360 20100
rect 39376 20156 39440 20160
rect 39376 20100 39380 20156
rect 39380 20100 39436 20156
rect 39436 20100 39440 20156
rect 39376 20096 39440 20100
rect 39456 20156 39520 20160
rect 39456 20100 39460 20156
rect 39460 20100 39516 20156
rect 39516 20100 39520 20156
rect 39456 20096 39520 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 14216 19612 14280 19616
rect 14216 19556 14220 19612
rect 14220 19556 14276 19612
rect 14276 19556 14280 19612
rect 14216 19552 14280 19556
rect 14296 19612 14360 19616
rect 14296 19556 14300 19612
rect 14300 19556 14356 19612
rect 14356 19556 14360 19612
rect 14296 19552 14360 19556
rect 14376 19612 14440 19616
rect 14376 19556 14380 19612
rect 14380 19556 14436 19612
rect 14436 19556 14440 19612
rect 14376 19552 14440 19556
rect 14456 19612 14520 19616
rect 14456 19556 14460 19612
rect 14460 19556 14516 19612
rect 14516 19556 14520 19612
rect 14456 19552 14520 19556
rect 24216 19612 24280 19616
rect 24216 19556 24220 19612
rect 24220 19556 24276 19612
rect 24276 19556 24280 19612
rect 24216 19552 24280 19556
rect 24296 19612 24360 19616
rect 24296 19556 24300 19612
rect 24300 19556 24356 19612
rect 24356 19556 24360 19612
rect 24296 19552 24360 19556
rect 24376 19612 24440 19616
rect 24376 19556 24380 19612
rect 24380 19556 24436 19612
rect 24436 19556 24440 19612
rect 24376 19552 24440 19556
rect 24456 19612 24520 19616
rect 24456 19556 24460 19612
rect 24460 19556 24516 19612
rect 24516 19556 24520 19612
rect 24456 19552 24520 19556
rect 34216 19612 34280 19616
rect 34216 19556 34220 19612
rect 34220 19556 34276 19612
rect 34276 19556 34280 19612
rect 34216 19552 34280 19556
rect 34296 19612 34360 19616
rect 34296 19556 34300 19612
rect 34300 19556 34356 19612
rect 34356 19556 34360 19612
rect 34296 19552 34360 19556
rect 34376 19612 34440 19616
rect 34376 19556 34380 19612
rect 34380 19556 34436 19612
rect 34436 19556 34440 19612
rect 34376 19552 34440 19556
rect 34456 19612 34520 19616
rect 34456 19556 34460 19612
rect 34460 19556 34516 19612
rect 34516 19556 34520 19612
rect 34456 19552 34520 19556
rect 44216 19612 44280 19616
rect 44216 19556 44220 19612
rect 44220 19556 44276 19612
rect 44276 19556 44280 19612
rect 44216 19552 44280 19556
rect 44296 19612 44360 19616
rect 44296 19556 44300 19612
rect 44300 19556 44356 19612
rect 44356 19556 44360 19612
rect 44296 19552 44360 19556
rect 44376 19612 44440 19616
rect 44376 19556 44380 19612
rect 44380 19556 44436 19612
rect 44436 19556 44440 19612
rect 44376 19552 44440 19556
rect 44456 19612 44520 19616
rect 44456 19556 44460 19612
rect 44460 19556 44516 19612
rect 44516 19556 44520 19612
rect 44456 19552 44520 19556
rect 9216 19068 9280 19072
rect 9216 19012 9220 19068
rect 9220 19012 9276 19068
rect 9276 19012 9280 19068
rect 9216 19008 9280 19012
rect 9296 19068 9360 19072
rect 9296 19012 9300 19068
rect 9300 19012 9356 19068
rect 9356 19012 9360 19068
rect 9296 19008 9360 19012
rect 9376 19068 9440 19072
rect 9376 19012 9380 19068
rect 9380 19012 9436 19068
rect 9436 19012 9440 19068
rect 9376 19008 9440 19012
rect 9456 19068 9520 19072
rect 9456 19012 9460 19068
rect 9460 19012 9516 19068
rect 9516 19012 9520 19068
rect 9456 19008 9520 19012
rect 39216 19068 39280 19072
rect 39216 19012 39220 19068
rect 39220 19012 39276 19068
rect 39276 19012 39280 19068
rect 39216 19008 39280 19012
rect 39296 19068 39360 19072
rect 39296 19012 39300 19068
rect 39300 19012 39356 19068
rect 39356 19012 39360 19068
rect 39296 19008 39360 19012
rect 39376 19068 39440 19072
rect 39376 19012 39380 19068
rect 39380 19012 39436 19068
rect 39436 19012 39440 19068
rect 39376 19008 39440 19012
rect 39456 19068 39520 19072
rect 39456 19012 39460 19068
rect 39460 19012 39516 19068
rect 39516 19012 39520 19068
rect 39456 19008 39520 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 14216 18524 14280 18528
rect 14216 18468 14220 18524
rect 14220 18468 14276 18524
rect 14276 18468 14280 18524
rect 14216 18464 14280 18468
rect 14296 18524 14360 18528
rect 14296 18468 14300 18524
rect 14300 18468 14356 18524
rect 14356 18468 14360 18524
rect 14296 18464 14360 18468
rect 14376 18524 14440 18528
rect 14376 18468 14380 18524
rect 14380 18468 14436 18524
rect 14436 18468 14440 18524
rect 14376 18464 14440 18468
rect 14456 18524 14520 18528
rect 14456 18468 14460 18524
rect 14460 18468 14516 18524
rect 14516 18468 14520 18524
rect 14456 18464 14520 18468
rect 44216 18524 44280 18528
rect 44216 18468 44220 18524
rect 44220 18468 44276 18524
rect 44276 18468 44280 18524
rect 44216 18464 44280 18468
rect 44296 18524 44360 18528
rect 44296 18468 44300 18524
rect 44300 18468 44356 18524
rect 44356 18468 44360 18524
rect 44296 18464 44360 18468
rect 44376 18524 44440 18528
rect 44376 18468 44380 18524
rect 44380 18468 44436 18524
rect 44436 18468 44440 18524
rect 44376 18464 44440 18468
rect 44456 18524 44520 18528
rect 44456 18468 44460 18524
rect 44460 18468 44516 18524
rect 44516 18468 44520 18524
rect 44456 18464 44520 18468
rect 9216 17980 9280 17984
rect 9216 17924 9220 17980
rect 9220 17924 9276 17980
rect 9276 17924 9280 17980
rect 9216 17920 9280 17924
rect 9296 17980 9360 17984
rect 9296 17924 9300 17980
rect 9300 17924 9356 17980
rect 9356 17924 9360 17980
rect 9296 17920 9360 17924
rect 9376 17980 9440 17984
rect 9376 17924 9380 17980
rect 9380 17924 9436 17980
rect 9436 17924 9440 17980
rect 9376 17920 9440 17924
rect 9456 17980 9520 17984
rect 9456 17924 9460 17980
rect 9460 17924 9516 17980
rect 9516 17924 9520 17980
rect 9456 17920 9520 17924
rect 39216 17980 39280 17984
rect 39216 17924 39220 17980
rect 39220 17924 39276 17980
rect 39276 17924 39280 17980
rect 39216 17920 39280 17924
rect 39296 17980 39360 17984
rect 39296 17924 39300 17980
rect 39300 17924 39356 17980
rect 39356 17924 39360 17980
rect 39296 17920 39360 17924
rect 39376 17980 39440 17984
rect 39376 17924 39380 17980
rect 39380 17924 39436 17980
rect 39436 17924 39440 17980
rect 39376 17920 39440 17924
rect 39456 17980 39520 17984
rect 39456 17924 39460 17980
rect 39460 17924 39516 17980
rect 39516 17924 39520 17980
rect 39456 17920 39520 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 14216 17436 14280 17440
rect 14216 17380 14220 17436
rect 14220 17380 14276 17436
rect 14276 17380 14280 17436
rect 14216 17376 14280 17380
rect 14296 17436 14360 17440
rect 14296 17380 14300 17436
rect 14300 17380 14356 17436
rect 14356 17380 14360 17436
rect 14296 17376 14360 17380
rect 14376 17436 14440 17440
rect 14376 17380 14380 17436
rect 14380 17380 14436 17436
rect 14436 17380 14440 17436
rect 14376 17376 14440 17380
rect 14456 17436 14520 17440
rect 14456 17380 14460 17436
rect 14460 17380 14516 17436
rect 14516 17380 14520 17436
rect 14456 17376 14520 17380
rect 44216 17436 44280 17440
rect 44216 17380 44220 17436
rect 44220 17380 44276 17436
rect 44276 17380 44280 17436
rect 44216 17376 44280 17380
rect 44296 17436 44360 17440
rect 44296 17380 44300 17436
rect 44300 17380 44356 17436
rect 44356 17380 44360 17436
rect 44296 17376 44360 17380
rect 44376 17436 44440 17440
rect 44376 17380 44380 17436
rect 44380 17380 44436 17436
rect 44436 17380 44440 17436
rect 44376 17376 44440 17380
rect 44456 17436 44520 17440
rect 44456 17380 44460 17436
rect 44460 17380 44516 17436
rect 44516 17380 44520 17436
rect 44456 17376 44520 17380
rect 9216 16892 9280 16896
rect 9216 16836 9220 16892
rect 9220 16836 9276 16892
rect 9276 16836 9280 16892
rect 9216 16832 9280 16836
rect 9296 16892 9360 16896
rect 9296 16836 9300 16892
rect 9300 16836 9356 16892
rect 9356 16836 9360 16892
rect 9296 16832 9360 16836
rect 9376 16892 9440 16896
rect 9376 16836 9380 16892
rect 9380 16836 9436 16892
rect 9436 16836 9440 16892
rect 9376 16832 9440 16836
rect 9456 16892 9520 16896
rect 9456 16836 9460 16892
rect 9460 16836 9516 16892
rect 9516 16836 9520 16892
rect 9456 16832 9520 16836
rect 39216 16892 39280 16896
rect 39216 16836 39220 16892
rect 39220 16836 39276 16892
rect 39276 16836 39280 16892
rect 39216 16832 39280 16836
rect 39296 16892 39360 16896
rect 39296 16836 39300 16892
rect 39300 16836 39356 16892
rect 39356 16836 39360 16892
rect 39296 16832 39360 16836
rect 39376 16892 39440 16896
rect 39376 16836 39380 16892
rect 39380 16836 39436 16892
rect 39436 16836 39440 16892
rect 39376 16832 39440 16836
rect 39456 16892 39520 16896
rect 39456 16836 39460 16892
rect 39460 16836 39516 16892
rect 39516 16836 39520 16892
rect 39456 16832 39520 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 14216 16348 14280 16352
rect 14216 16292 14220 16348
rect 14220 16292 14276 16348
rect 14276 16292 14280 16348
rect 14216 16288 14280 16292
rect 14296 16348 14360 16352
rect 14296 16292 14300 16348
rect 14300 16292 14356 16348
rect 14356 16292 14360 16348
rect 14296 16288 14360 16292
rect 14376 16348 14440 16352
rect 14376 16292 14380 16348
rect 14380 16292 14436 16348
rect 14436 16292 14440 16348
rect 14376 16288 14440 16292
rect 14456 16348 14520 16352
rect 14456 16292 14460 16348
rect 14460 16292 14516 16348
rect 14516 16292 14520 16348
rect 14456 16288 14520 16292
rect 29216 16054 29520 16438
rect 44216 16348 44280 16352
rect 44216 16292 44220 16348
rect 44220 16292 44276 16348
rect 44276 16292 44280 16348
rect 44216 16288 44280 16292
rect 44296 16348 44360 16352
rect 44296 16292 44300 16348
rect 44300 16292 44356 16348
rect 44356 16292 44360 16348
rect 44296 16288 44360 16292
rect 44376 16348 44440 16352
rect 44376 16292 44380 16348
rect 44380 16292 44436 16348
rect 44436 16292 44440 16348
rect 44376 16288 44440 16292
rect 44456 16348 44520 16352
rect 44456 16292 44460 16348
rect 44460 16292 44516 16348
rect 44516 16292 44520 16348
rect 44456 16288 44520 16292
rect 9216 15804 9280 15808
rect 9216 15748 9220 15804
rect 9220 15748 9276 15804
rect 9276 15748 9280 15804
rect 9216 15744 9280 15748
rect 9296 15804 9360 15808
rect 9296 15748 9300 15804
rect 9300 15748 9356 15804
rect 9356 15748 9360 15804
rect 9296 15744 9360 15748
rect 9376 15804 9440 15808
rect 9376 15748 9380 15804
rect 9380 15748 9436 15804
rect 9436 15748 9440 15804
rect 9376 15744 9440 15748
rect 9456 15804 9520 15808
rect 9456 15748 9460 15804
rect 9460 15748 9516 15804
rect 9516 15748 9520 15804
rect 9456 15744 9520 15748
rect 39216 15804 39280 15808
rect 39216 15748 39220 15804
rect 39220 15748 39276 15804
rect 39276 15748 39280 15804
rect 39216 15744 39280 15748
rect 39296 15804 39360 15808
rect 39296 15748 39300 15804
rect 39300 15748 39356 15804
rect 39356 15748 39360 15804
rect 39296 15744 39360 15748
rect 39376 15804 39440 15808
rect 39376 15748 39380 15804
rect 39380 15748 39436 15804
rect 39436 15748 39440 15804
rect 39376 15744 39440 15748
rect 39456 15804 39520 15808
rect 39456 15748 39460 15804
rect 39460 15748 39516 15804
rect 39516 15748 39520 15804
rect 39456 15744 39520 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 14216 15260 14280 15264
rect 14216 15204 14220 15260
rect 14220 15204 14276 15260
rect 14276 15204 14280 15260
rect 14216 15200 14280 15204
rect 14296 15260 14360 15264
rect 14296 15204 14300 15260
rect 14300 15204 14356 15260
rect 14356 15204 14360 15260
rect 14296 15200 14360 15204
rect 14376 15260 14440 15264
rect 14376 15204 14380 15260
rect 14380 15204 14436 15260
rect 14436 15204 14440 15260
rect 14376 15200 14440 15204
rect 14456 15260 14520 15264
rect 14456 15204 14460 15260
rect 14460 15204 14516 15260
rect 14516 15204 14520 15260
rect 14456 15200 14520 15204
rect 24216 15254 24520 15638
rect 44216 15260 44280 15264
rect 44216 15204 44220 15260
rect 44220 15204 44276 15260
rect 44276 15204 44280 15260
rect 44216 15200 44280 15204
rect 44296 15260 44360 15264
rect 44296 15204 44300 15260
rect 44300 15204 44356 15260
rect 44356 15204 44360 15260
rect 44296 15200 44360 15204
rect 44376 15260 44440 15264
rect 44376 15204 44380 15260
rect 44380 15204 44436 15260
rect 44436 15204 44440 15260
rect 44376 15200 44440 15204
rect 44456 15260 44520 15264
rect 44456 15204 44460 15260
rect 44460 15204 44516 15260
rect 44516 15204 44520 15260
rect 44456 15200 44520 15204
rect 9216 14716 9280 14720
rect 9216 14660 9220 14716
rect 9220 14660 9276 14716
rect 9276 14660 9280 14716
rect 9216 14656 9280 14660
rect 9296 14716 9360 14720
rect 9296 14660 9300 14716
rect 9300 14660 9356 14716
rect 9356 14660 9360 14716
rect 9296 14656 9360 14660
rect 9376 14716 9440 14720
rect 9376 14660 9380 14716
rect 9380 14660 9436 14716
rect 9436 14660 9440 14716
rect 9376 14656 9440 14660
rect 9456 14716 9520 14720
rect 9456 14660 9460 14716
rect 9460 14660 9516 14716
rect 9516 14660 9520 14716
rect 9456 14656 9520 14660
rect 39216 14716 39280 14720
rect 39216 14660 39220 14716
rect 39220 14660 39276 14716
rect 39276 14660 39280 14716
rect 39216 14656 39280 14660
rect 39296 14716 39360 14720
rect 39296 14660 39300 14716
rect 39300 14660 39356 14716
rect 39356 14660 39360 14716
rect 39296 14656 39360 14660
rect 39376 14716 39440 14720
rect 39376 14660 39380 14716
rect 39380 14660 39436 14716
rect 39436 14660 39440 14716
rect 39376 14656 39440 14660
rect 39456 14716 39520 14720
rect 39456 14660 39460 14716
rect 39460 14660 39516 14716
rect 39516 14660 39520 14716
rect 39456 14656 39520 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 14216 14172 14280 14176
rect 14216 14116 14220 14172
rect 14220 14116 14276 14172
rect 14276 14116 14280 14172
rect 14216 14112 14280 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 44216 14172 44280 14176
rect 44216 14116 44220 14172
rect 44220 14116 44276 14172
rect 44276 14116 44280 14172
rect 44216 14112 44280 14116
rect 44296 14172 44360 14176
rect 44296 14116 44300 14172
rect 44300 14116 44356 14172
rect 44356 14116 44360 14172
rect 44296 14112 44360 14116
rect 44376 14172 44440 14176
rect 44376 14116 44380 14172
rect 44380 14116 44436 14172
rect 44436 14116 44440 14172
rect 44376 14112 44440 14116
rect 44456 14172 44520 14176
rect 44456 14116 44460 14172
rect 44460 14116 44516 14172
rect 44516 14116 44520 14172
rect 44456 14112 44520 14116
rect 9216 13628 9280 13632
rect 9216 13572 9220 13628
rect 9220 13572 9276 13628
rect 9276 13572 9280 13628
rect 9216 13568 9280 13572
rect 9296 13628 9360 13632
rect 9296 13572 9300 13628
rect 9300 13572 9356 13628
rect 9356 13572 9360 13628
rect 9296 13568 9360 13572
rect 9376 13628 9440 13632
rect 9376 13572 9380 13628
rect 9380 13572 9436 13628
rect 9436 13572 9440 13628
rect 9376 13568 9440 13572
rect 9456 13628 9520 13632
rect 9456 13572 9460 13628
rect 9460 13572 9516 13628
rect 9516 13572 9520 13628
rect 9456 13568 9520 13572
rect 39216 13628 39280 13632
rect 39216 13572 39220 13628
rect 39220 13572 39276 13628
rect 39276 13572 39280 13628
rect 39216 13568 39280 13572
rect 39296 13628 39360 13632
rect 39296 13572 39300 13628
rect 39300 13572 39356 13628
rect 39356 13572 39360 13628
rect 39296 13568 39360 13572
rect 39376 13628 39440 13632
rect 39376 13572 39380 13628
rect 39380 13572 39436 13628
rect 39436 13572 39440 13628
rect 39376 13568 39440 13572
rect 39456 13628 39520 13632
rect 39456 13572 39460 13628
rect 39460 13572 39516 13628
rect 39516 13572 39520 13628
rect 39456 13568 39520 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 14216 13084 14280 13088
rect 14216 13028 14220 13084
rect 14220 13028 14276 13084
rect 14276 13028 14280 13084
rect 14216 13024 14280 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 44216 13084 44280 13088
rect 44216 13028 44220 13084
rect 44220 13028 44276 13084
rect 44276 13028 44280 13084
rect 44216 13024 44280 13028
rect 44296 13084 44360 13088
rect 44296 13028 44300 13084
rect 44300 13028 44356 13084
rect 44356 13028 44360 13084
rect 44296 13024 44360 13028
rect 44376 13084 44440 13088
rect 44376 13028 44380 13084
rect 44380 13028 44436 13084
rect 44436 13028 44440 13084
rect 44376 13024 44440 13028
rect 44456 13084 44520 13088
rect 44456 13028 44460 13084
rect 44460 13028 44516 13084
rect 44516 13028 44520 13084
rect 44456 13024 44520 13028
rect 9216 12540 9280 12544
rect 9216 12484 9220 12540
rect 9220 12484 9276 12540
rect 9276 12484 9280 12540
rect 9216 12480 9280 12484
rect 9296 12540 9360 12544
rect 9296 12484 9300 12540
rect 9300 12484 9356 12540
rect 9356 12484 9360 12540
rect 9296 12480 9360 12484
rect 9376 12540 9440 12544
rect 9376 12484 9380 12540
rect 9380 12484 9436 12540
rect 9436 12484 9440 12540
rect 9376 12480 9440 12484
rect 9456 12540 9520 12544
rect 9456 12484 9460 12540
rect 9460 12484 9516 12540
rect 9516 12484 9520 12540
rect 9456 12480 9520 12484
rect 39216 12540 39280 12544
rect 39216 12484 39220 12540
rect 39220 12484 39276 12540
rect 39276 12484 39280 12540
rect 39216 12480 39280 12484
rect 39296 12540 39360 12544
rect 39296 12484 39300 12540
rect 39300 12484 39356 12540
rect 39356 12484 39360 12540
rect 39296 12480 39360 12484
rect 39376 12540 39440 12544
rect 39376 12484 39380 12540
rect 39380 12484 39436 12540
rect 39436 12484 39440 12540
rect 39376 12480 39440 12484
rect 39456 12540 39520 12544
rect 39456 12484 39460 12540
rect 39460 12484 39516 12540
rect 39516 12484 39520 12540
rect 39456 12480 39520 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 14216 11996 14280 12000
rect 14216 11940 14220 11996
rect 14220 11940 14276 11996
rect 14276 11940 14280 11996
rect 14216 11936 14280 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 44216 11996 44280 12000
rect 44216 11940 44220 11996
rect 44220 11940 44276 11996
rect 44276 11940 44280 11996
rect 44216 11936 44280 11940
rect 44296 11996 44360 12000
rect 44296 11940 44300 11996
rect 44300 11940 44356 11996
rect 44356 11940 44360 11996
rect 44296 11936 44360 11940
rect 44376 11996 44440 12000
rect 44376 11940 44380 11996
rect 44380 11940 44436 11996
rect 44436 11940 44440 11996
rect 44376 11936 44440 11940
rect 44456 11996 44520 12000
rect 44456 11940 44460 11996
rect 44460 11940 44516 11996
rect 44516 11940 44520 11996
rect 44456 11936 44520 11940
rect 24216 11603 24520 11907
rect 34216 11603 34520 11907
rect 9216 11452 9280 11456
rect 9216 11396 9220 11452
rect 9220 11396 9276 11452
rect 9276 11396 9280 11452
rect 9216 11392 9280 11396
rect 9296 11452 9360 11456
rect 9296 11396 9300 11452
rect 9300 11396 9356 11452
rect 9356 11396 9360 11452
rect 9296 11392 9360 11396
rect 9376 11452 9440 11456
rect 9376 11396 9380 11452
rect 9380 11396 9436 11452
rect 9436 11396 9440 11452
rect 9376 11392 9440 11396
rect 9456 11452 9520 11456
rect 9456 11396 9460 11452
rect 9460 11396 9516 11452
rect 9516 11396 9520 11452
rect 9456 11392 9520 11396
rect 39216 11452 39280 11456
rect 39216 11396 39220 11452
rect 39220 11396 39276 11452
rect 39276 11396 39280 11452
rect 39216 11392 39280 11396
rect 39296 11452 39360 11456
rect 39296 11396 39300 11452
rect 39300 11396 39356 11452
rect 39356 11396 39360 11452
rect 39296 11392 39360 11396
rect 39376 11452 39440 11456
rect 39376 11396 39380 11452
rect 39380 11396 39436 11452
rect 39436 11396 39440 11452
rect 39376 11392 39440 11396
rect 39456 11452 39520 11456
rect 39456 11396 39460 11452
rect 39460 11396 39516 11452
rect 39516 11396 39520 11452
rect 39456 11392 39520 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 14216 10908 14280 10912
rect 14216 10852 14220 10908
rect 14220 10852 14276 10908
rect 14276 10852 14280 10908
rect 14216 10848 14280 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 44216 10908 44280 10912
rect 44216 10852 44220 10908
rect 44220 10852 44276 10908
rect 44276 10852 44280 10908
rect 44216 10848 44280 10852
rect 44296 10908 44360 10912
rect 44296 10852 44300 10908
rect 44300 10852 44356 10908
rect 44356 10852 44360 10908
rect 44296 10848 44360 10852
rect 44376 10908 44440 10912
rect 44376 10852 44380 10908
rect 44380 10852 44436 10908
rect 44436 10852 44440 10908
rect 44376 10848 44440 10852
rect 44456 10908 44520 10912
rect 44456 10852 44460 10908
rect 44460 10852 44516 10908
rect 44516 10852 44520 10908
rect 44456 10848 44520 10852
rect 9216 10364 9280 10368
rect 9216 10308 9220 10364
rect 9220 10308 9276 10364
rect 9276 10308 9280 10364
rect 9216 10304 9280 10308
rect 9296 10364 9360 10368
rect 9296 10308 9300 10364
rect 9300 10308 9356 10364
rect 9356 10308 9360 10364
rect 9296 10304 9360 10308
rect 9376 10364 9440 10368
rect 9376 10308 9380 10364
rect 9380 10308 9436 10364
rect 9436 10308 9440 10364
rect 9376 10304 9440 10308
rect 9456 10364 9520 10368
rect 9456 10308 9460 10364
rect 9460 10308 9516 10364
rect 9516 10308 9520 10364
rect 9456 10304 9520 10308
rect 29216 10329 29520 10633
rect 39216 10364 39280 10368
rect 39216 10308 39220 10364
rect 39220 10308 39276 10364
rect 39276 10308 39280 10364
rect 39216 10304 39280 10308
rect 39296 10364 39360 10368
rect 39296 10308 39300 10364
rect 39300 10308 39356 10364
rect 39356 10308 39360 10364
rect 39296 10304 39360 10308
rect 39376 10364 39440 10368
rect 39376 10308 39380 10364
rect 39380 10308 39436 10364
rect 39436 10308 39440 10364
rect 39376 10304 39440 10308
rect 39456 10364 39520 10368
rect 39456 10308 39460 10364
rect 39460 10308 39516 10364
rect 39516 10308 39520 10364
rect 39456 10304 39520 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 14216 9820 14280 9824
rect 14216 9764 14220 9820
rect 14220 9764 14276 9820
rect 14276 9764 14280 9820
rect 14216 9760 14280 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 44216 9820 44280 9824
rect 44216 9764 44220 9820
rect 44220 9764 44276 9820
rect 44276 9764 44280 9820
rect 44216 9760 44280 9764
rect 44296 9820 44360 9824
rect 44296 9764 44300 9820
rect 44300 9764 44356 9820
rect 44356 9764 44360 9820
rect 44296 9760 44360 9764
rect 44376 9820 44440 9824
rect 44376 9764 44380 9820
rect 44380 9764 44436 9820
rect 44436 9764 44440 9820
rect 44376 9760 44440 9764
rect 44456 9820 44520 9824
rect 44456 9764 44460 9820
rect 44460 9764 44516 9820
rect 44516 9764 44520 9820
rect 44456 9760 44520 9764
rect 9216 9276 9280 9280
rect 9216 9220 9220 9276
rect 9220 9220 9276 9276
rect 9276 9220 9280 9276
rect 9216 9216 9280 9220
rect 9296 9276 9360 9280
rect 9296 9220 9300 9276
rect 9300 9220 9356 9276
rect 9356 9220 9360 9276
rect 9296 9216 9360 9220
rect 9376 9276 9440 9280
rect 9376 9220 9380 9276
rect 9380 9220 9436 9276
rect 9436 9220 9440 9276
rect 9376 9216 9440 9220
rect 9456 9276 9520 9280
rect 9456 9220 9460 9276
rect 9460 9220 9516 9276
rect 9516 9220 9520 9276
rect 9456 9216 9520 9220
rect 24216 9054 24520 9358
rect 34216 9054 34520 9358
rect 39216 9276 39280 9280
rect 39216 9220 39220 9276
rect 39220 9220 39276 9276
rect 39276 9220 39280 9276
rect 39216 9216 39280 9220
rect 39296 9276 39360 9280
rect 39296 9220 39300 9276
rect 39300 9220 39356 9276
rect 39356 9220 39360 9276
rect 39296 9216 39360 9220
rect 39376 9276 39440 9280
rect 39376 9220 39380 9276
rect 39380 9220 39436 9276
rect 39436 9220 39440 9276
rect 39376 9216 39440 9220
rect 39456 9276 39520 9280
rect 39456 9220 39460 9276
rect 39460 9220 39516 9276
rect 39516 9220 39520 9276
rect 39456 9216 39520 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 14216 8732 14280 8736
rect 14216 8676 14220 8732
rect 14220 8676 14276 8732
rect 14276 8676 14280 8732
rect 14216 8672 14280 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 44216 8732 44280 8736
rect 44216 8676 44220 8732
rect 44220 8676 44276 8732
rect 44276 8676 44280 8732
rect 44216 8672 44280 8676
rect 44296 8732 44360 8736
rect 44296 8676 44300 8732
rect 44300 8676 44356 8732
rect 44356 8676 44360 8732
rect 44296 8672 44360 8676
rect 44376 8732 44440 8736
rect 44376 8676 44380 8732
rect 44380 8676 44436 8732
rect 44436 8676 44440 8732
rect 44376 8672 44440 8676
rect 44456 8732 44520 8736
rect 44456 8676 44460 8732
rect 44460 8676 44516 8732
rect 44516 8676 44520 8732
rect 44456 8672 44520 8676
rect 9216 8188 9280 8192
rect 9216 8132 9220 8188
rect 9220 8132 9276 8188
rect 9276 8132 9280 8188
rect 9216 8128 9280 8132
rect 9296 8188 9360 8192
rect 9296 8132 9300 8188
rect 9300 8132 9356 8188
rect 9356 8132 9360 8188
rect 9296 8128 9360 8132
rect 9376 8188 9440 8192
rect 9376 8132 9380 8188
rect 9380 8132 9436 8188
rect 9436 8132 9440 8188
rect 9376 8128 9440 8132
rect 9456 8188 9520 8192
rect 9456 8132 9460 8188
rect 9460 8132 9516 8188
rect 9516 8132 9520 8188
rect 9456 8128 9520 8132
rect 39216 8188 39280 8192
rect 39216 8132 39220 8188
rect 39220 8132 39276 8188
rect 39276 8132 39280 8188
rect 39216 8128 39280 8132
rect 39296 8188 39360 8192
rect 39296 8132 39300 8188
rect 39300 8132 39356 8188
rect 39356 8132 39360 8188
rect 39296 8128 39360 8132
rect 39376 8188 39440 8192
rect 39376 8132 39380 8188
rect 39380 8132 39436 8188
rect 39436 8132 39440 8188
rect 39376 8128 39440 8132
rect 39456 8188 39520 8192
rect 39456 8132 39460 8188
rect 39460 8132 39516 8188
rect 39516 8132 39520 8188
rect 39456 8128 39520 8132
rect 29216 7779 29520 8083
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 14216 7644 14280 7648
rect 14216 7588 14220 7644
rect 14220 7588 14276 7644
rect 14276 7588 14280 7644
rect 14216 7584 14280 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 44216 7644 44280 7648
rect 44216 7588 44220 7644
rect 44220 7588 44276 7644
rect 44276 7588 44280 7644
rect 44216 7584 44280 7588
rect 44296 7644 44360 7648
rect 44296 7588 44300 7644
rect 44300 7588 44356 7644
rect 44356 7588 44360 7644
rect 44296 7584 44360 7588
rect 44376 7644 44440 7648
rect 44376 7588 44380 7644
rect 44380 7588 44436 7644
rect 44436 7588 44440 7644
rect 44376 7584 44440 7588
rect 44456 7644 44520 7648
rect 44456 7588 44460 7644
rect 44460 7588 44516 7644
rect 44516 7588 44520 7644
rect 44456 7584 44520 7588
rect 9216 7100 9280 7104
rect 9216 7044 9220 7100
rect 9220 7044 9276 7100
rect 9276 7044 9280 7100
rect 9216 7040 9280 7044
rect 9296 7100 9360 7104
rect 9296 7044 9300 7100
rect 9300 7044 9356 7100
rect 9356 7044 9360 7100
rect 9296 7040 9360 7044
rect 9376 7100 9440 7104
rect 9376 7044 9380 7100
rect 9380 7044 9436 7100
rect 9436 7044 9440 7100
rect 9376 7040 9440 7044
rect 9456 7100 9520 7104
rect 9456 7044 9460 7100
rect 9460 7044 9516 7100
rect 9516 7044 9520 7100
rect 9456 7040 9520 7044
rect 39216 7100 39280 7104
rect 39216 7044 39220 7100
rect 39220 7044 39276 7100
rect 39276 7044 39280 7100
rect 39216 7040 39280 7044
rect 39296 7100 39360 7104
rect 39296 7044 39300 7100
rect 39300 7044 39356 7100
rect 39356 7044 39360 7100
rect 39296 7040 39360 7044
rect 39376 7100 39440 7104
rect 39376 7044 39380 7100
rect 39380 7044 39436 7100
rect 39436 7044 39440 7100
rect 39376 7040 39440 7044
rect 39456 7100 39520 7104
rect 39456 7044 39460 7100
rect 39460 7044 39516 7100
rect 39516 7044 39520 7100
rect 39456 7040 39520 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 14216 6556 14280 6560
rect 14216 6500 14220 6556
rect 14220 6500 14276 6556
rect 14276 6500 14280 6556
rect 14216 6496 14280 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 24216 6505 24520 6809
rect 34216 6505 34520 6809
rect 44216 6556 44280 6560
rect 44216 6500 44220 6556
rect 44220 6500 44276 6556
rect 44276 6500 44280 6556
rect 44216 6496 44280 6500
rect 44296 6556 44360 6560
rect 44296 6500 44300 6556
rect 44300 6500 44356 6556
rect 44356 6500 44360 6556
rect 44296 6496 44360 6500
rect 44376 6556 44440 6560
rect 44376 6500 44380 6556
rect 44380 6500 44436 6556
rect 44436 6500 44440 6556
rect 44376 6496 44440 6500
rect 44456 6556 44520 6560
rect 44456 6500 44460 6556
rect 44460 6500 44516 6556
rect 44516 6500 44520 6556
rect 44456 6496 44520 6500
rect 9216 6012 9280 6016
rect 9216 5956 9220 6012
rect 9220 5956 9276 6012
rect 9276 5956 9280 6012
rect 9216 5952 9280 5956
rect 9296 6012 9360 6016
rect 9296 5956 9300 6012
rect 9300 5956 9356 6012
rect 9356 5956 9360 6012
rect 9296 5952 9360 5956
rect 9376 6012 9440 6016
rect 9376 5956 9380 6012
rect 9380 5956 9436 6012
rect 9436 5956 9440 6012
rect 9376 5952 9440 5956
rect 9456 6012 9520 6016
rect 9456 5956 9460 6012
rect 9460 5956 9516 6012
rect 9516 5956 9520 6012
rect 9456 5952 9520 5956
rect 39216 6012 39280 6016
rect 39216 5956 39220 6012
rect 39220 5956 39276 6012
rect 39276 5956 39280 6012
rect 39216 5952 39280 5956
rect 39296 6012 39360 6016
rect 39296 5956 39300 6012
rect 39300 5956 39356 6012
rect 39356 5956 39360 6012
rect 39296 5952 39360 5956
rect 39376 6012 39440 6016
rect 39376 5956 39380 6012
rect 39380 5956 39436 6012
rect 39436 5956 39440 6012
rect 39376 5952 39440 5956
rect 39456 6012 39520 6016
rect 39456 5956 39460 6012
rect 39460 5956 39516 6012
rect 39516 5956 39520 6012
rect 39456 5952 39520 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 14216 5468 14280 5472
rect 14216 5412 14220 5468
rect 14220 5412 14276 5468
rect 14276 5412 14280 5468
rect 14216 5408 14280 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 44216 5468 44280 5472
rect 44216 5412 44220 5468
rect 44220 5412 44276 5468
rect 44276 5412 44280 5468
rect 44216 5408 44280 5412
rect 44296 5468 44360 5472
rect 44296 5412 44300 5468
rect 44300 5412 44356 5468
rect 44356 5412 44360 5468
rect 44296 5408 44360 5412
rect 44376 5468 44440 5472
rect 44376 5412 44380 5468
rect 44380 5412 44436 5468
rect 44436 5412 44440 5468
rect 44376 5408 44440 5412
rect 44456 5468 44520 5472
rect 44456 5412 44460 5468
rect 44460 5412 44516 5468
rect 44516 5412 44520 5468
rect 44456 5408 44520 5412
rect 9216 4924 9280 4928
rect 9216 4868 9220 4924
rect 9220 4868 9276 4924
rect 9276 4868 9280 4924
rect 9216 4864 9280 4868
rect 9296 4924 9360 4928
rect 9296 4868 9300 4924
rect 9300 4868 9356 4924
rect 9356 4868 9360 4924
rect 9296 4864 9360 4868
rect 9376 4924 9440 4928
rect 9376 4868 9380 4924
rect 9380 4868 9436 4924
rect 9436 4868 9440 4924
rect 9376 4864 9440 4868
rect 9456 4924 9520 4928
rect 9456 4868 9460 4924
rect 9460 4868 9516 4924
rect 9516 4868 9520 4924
rect 9456 4864 9520 4868
rect 39216 4924 39280 4928
rect 39216 4868 39220 4924
rect 39220 4868 39276 4924
rect 39276 4868 39280 4924
rect 39216 4864 39280 4868
rect 39296 4924 39360 4928
rect 39296 4868 39300 4924
rect 39300 4868 39356 4924
rect 39356 4868 39360 4924
rect 39296 4864 39360 4868
rect 39376 4924 39440 4928
rect 39376 4868 39380 4924
rect 39380 4868 39436 4924
rect 39436 4868 39440 4924
rect 39376 4864 39440 4868
rect 39456 4924 39520 4928
rect 39456 4868 39460 4924
rect 39460 4868 39516 4924
rect 39516 4868 39520 4924
rect 39456 4864 39520 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 14216 4380 14280 4384
rect 14216 4324 14220 4380
rect 14220 4324 14276 4380
rect 14276 4324 14280 4380
rect 14216 4320 14280 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 44216 4380 44280 4384
rect 44216 4324 44220 4380
rect 44220 4324 44276 4380
rect 44276 4324 44280 4380
rect 44216 4320 44280 4324
rect 44296 4380 44360 4384
rect 44296 4324 44300 4380
rect 44300 4324 44356 4380
rect 44356 4324 44360 4380
rect 44296 4320 44360 4324
rect 44376 4380 44440 4384
rect 44376 4324 44380 4380
rect 44380 4324 44436 4380
rect 44436 4324 44440 4380
rect 44376 4320 44440 4324
rect 44456 4380 44520 4384
rect 44456 4324 44460 4380
rect 44460 4324 44516 4380
rect 44516 4324 44520 4380
rect 44456 4320 44520 4324
rect 9216 3836 9280 3840
rect 9216 3780 9220 3836
rect 9220 3780 9276 3836
rect 9276 3780 9280 3836
rect 9216 3776 9280 3780
rect 9296 3836 9360 3840
rect 9296 3780 9300 3836
rect 9300 3780 9356 3836
rect 9356 3780 9360 3836
rect 9296 3776 9360 3780
rect 9376 3836 9440 3840
rect 9376 3780 9380 3836
rect 9380 3780 9436 3836
rect 9436 3780 9440 3836
rect 9376 3776 9440 3780
rect 9456 3836 9520 3840
rect 9456 3780 9460 3836
rect 9460 3780 9516 3836
rect 9516 3780 9520 3836
rect 9456 3776 9520 3780
rect 39216 3836 39280 3840
rect 39216 3780 39220 3836
rect 39220 3780 39276 3836
rect 39276 3780 39280 3836
rect 39216 3776 39280 3780
rect 39296 3836 39360 3840
rect 39296 3780 39300 3836
rect 39300 3780 39356 3836
rect 39356 3780 39360 3836
rect 39296 3776 39360 3780
rect 39376 3836 39440 3840
rect 39376 3780 39380 3836
rect 39380 3780 39436 3836
rect 39436 3780 39440 3836
rect 39376 3776 39440 3780
rect 39456 3836 39520 3840
rect 39456 3780 39460 3836
rect 39460 3780 39516 3836
rect 39516 3780 39520 3836
rect 39456 3776 39520 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 14216 3292 14280 3296
rect 14216 3236 14220 3292
rect 14220 3236 14276 3292
rect 14276 3236 14280 3292
rect 14216 3232 14280 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 44216 3292 44280 3296
rect 44216 3236 44220 3292
rect 44220 3236 44276 3292
rect 44276 3236 44280 3292
rect 44216 3232 44280 3236
rect 44296 3292 44360 3296
rect 44296 3236 44300 3292
rect 44300 3236 44356 3292
rect 44356 3236 44360 3292
rect 44296 3232 44360 3236
rect 44376 3292 44440 3296
rect 44376 3236 44380 3292
rect 44380 3236 44436 3292
rect 44436 3236 44440 3292
rect 44376 3232 44440 3236
rect 44456 3292 44520 3296
rect 44456 3236 44460 3292
rect 44460 3236 44516 3292
rect 44516 3236 44520 3292
rect 44456 3232 44520 3236
rect 24216 2838 24520 3222
rect 9216 2748 9280 2752
rect 9216 2692 9220 2748
rect 9220 2692 9276 2748
rect 9276 2692 9280 2748
rect 9216 2688 9280 2692
rect 9296 2748 9360 2752
rect 9296 2692 9300 2748
rect 9300 2692 9356 2748
rect 9356 2692 9360 2748
rect 9296 2688 9360 2692
rect 9376 2748 9440 2752
rect 9376 2692 9380 2748
rect 9380 2692 9436 2748
rect 9436 2692 9440 2748
rect 9376 2688 9440 2692
rect 9456 2748 9520 2752
rect 9456 2692 9460 2748
rect 9460 2692 9516 2748
rect 9516 2692 9520 2748
rect 9456 2688 9520 2692
rect 39216 2748 39280 2752
rect 39216 2692 39220 2748
rect 39220 2692 39276 2748
rect 39276 2692 39280 2748
rect 39216 2688 39280 2692
rect 39296 2748 39360 2752
rect 39296 2692 39300 2748
rect 39300 2692 39356 2748
rect 39356 2692 39360 2748
rect 39296 2688 39360 2692
rect 39376 2748 39440 2752
rect 39376 2692 39380 2748
rect 39380 2692 39436 2748
rect 39436 2692 39440 2748
rect 39376 2688 39440 2692
rect 39456 2748 39520 2752
rect 39456 2692 39460 2748
rect 39460 2692 39516 2748
rect 39516 2692 39520 2748
rect 39456 2688 39520 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 14216 2204 14280 2208
rect 14216 2148 14220 2204
rect 14220 2148 14276 2204
rect 14276 2148 14280 2204
rect 14216 2144 14280 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 29216 2206 29520 2430
rect 44216 2204 44280 2208
rect 44216 2148 44220 2204
rect 44220 2148 44276 2204
rect 44276 2148 44280 2204
rect 44216 2144 44280 2148
rect 44296 2204 44360 2208
rect 44296 2148 44300 2204
rect 44300 2148 44356 2204
rect 44356 2148 44360 2204
rect 44296 2144 44360 2148
rect 44376 2204 44440 2208
rect 44376 2148 44380 2204
rect 44380 2148 44436 2204
rect 44436 2148 44440 2204
rect 44376 2144 44440 2148
rect 44456 2204 44520 2208
rect 44456 2148 44460 2204
rect 44460 2148 44516 2204
rect 44516 2148 44520 2204
rect 44456 2144 44520 2148
<< metal4 >>
rect 4208 46816 4528 47376
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 9208 47360 9528 47376
rect 9208 47296 9216 47360
rect 9280 47296 9296 47360
rect 9360 47296 9376 47360
rect 9440 47296 9456 47360
rect 9520 47296 9528 47360
rect 9208 46272 9528 47296
rect 9208 46208 9216 46272
rect 9280 46208 9296 46272
rect 9360 46208 9376 46272
rect 9440 46208 9456 46272
rect 9520 46208 9528 46272
rect 9208 45184 9528 46208
rect 9208 45120 9216 45184
rect 9280 45120 9296 45184
rect 9360 45120 9376 45184
rect 9440 45120 9456 45184
rect 9520 45120 9528 45184
rect 9208 44096 9528 45120
rect 9208 44032 9216 44096
rect 9280 44032 9296 44096
rect 9360 44032 9376 44096
rect 9440 44032 9456 44096
rect 9520 44032 9528 44096
rect 9208 43008 9528 44032
rect 9208 42944 9216 43008
rect 9280 42944 9296 43008
rect 9360 42944 9376 43008
rect 9440 42944 9456 43008
rect 9520 42944 9528 43008
rect 9208 41920 9528 42944
rect 9208 41856 9216 41920
rect 9280 41856 9296 41920
rect 9360 41856 9376 41920
rect 9440 41856 9456 41920
rect 9520 41856 9528 41920
rect 9208 40832 9528 41856
rect 9208 40768 9216 40832
rect 9280 40768 9296 40832
rect 9360 40768 9376 40832
rect 9440 40768 9456 40832
rect 9520 40768 9528 40832
rect 9208 39744 9528 40768
rect 9208 39680 9216 39744
rect 9280 39680 9296 39744
rect 9360 39680 9376 39744
rect 9440 39680 9456 39744
rect 9520 39680 9528 39744
rect 9208 38656 9528 39680
rect 9208 38592 9216 38656
rect 9280 38592 9296 38656
rect 9360 38592 9376 38656
rect 9440 38592 9456 38656
rect 9520 38592 9528 38656
rect 9208 37568 9528 38592
rect 9208 37504 9216 37568
rect 9280 37504 9296 37568
rect 9360 37504 9376 37568
rect 9440 37504 9456 37568
rect 9520 37504 9528 37568
rect 9208 36480 9528 37504
rect 9208 36416 9216 36480
rect 9280 36416 9296 36480
rect 9360 36416 9376 36480
rect 9440 36416 9456 36480
rect 9520 36416 9528 36480
rect 9208 35392 9528 36416
rect 9208 35328 9216 35392
rect 9280 35328 9296 35392
rect 9360 35328 9376 35392
rect 9440 35328 9456 35392
rect 9520 35328 9528 35392
rect 9208 34304 9528 35328
rect 9208 34240 9216 34304
rect 9280 34240 9296 34304
rect 9360 34240 9376 34304
rect 9440 34240 9456 34304
rect 9520 34240 9528 34304
rect 9208 33216 9528 34240
rect 9208 33152 9216 33216
rect 9280 33152 9296 33216
rect 9360 33152 9376 33216
rect 9440 33152 9456 33216
rect 9520 33152 9528 33216
rect 9208 32128 9528 33152
rect 9208 32064 9216 32128
rect 9280 32064 9296 32128
rect 9360 32064 9376 32128
rect 9440 32064 9456 32128
rect 9520 32064 9528 32128
rect 9208 31040 9528 32064
rect 9208 30976 9216 31040
rect 9280 30976 9296 31040
rect 9360 30976 9376 31040
rect 9440 30976 9456 31040
rect 9520 30976 9528 31040
rect 9208 29952 9528 30976
rect 9208 29888 9216 29952
rect 9280 29888 9296 29952
rect 9360 29888 9376 29952
rect 9440 29888 9456 29952
rect 9520 29888 9528 29952
rect 9208 28864 9528 29888
rect 9208 28800 9216 28864
rect 9280 28800 9296 28864
rect 9360 28800 9376 28864
rect 9440 28800 9456 28864
rect 9520 28800 9528 28864
rect 9208 27776 9528 28800
rect 9208 27712 9216 27776
rect 9280 27712 9296 27776
rect 9360 27712 9376 27776
rect 9440 27712 9456 27776
rect 9520 27712 9528 27776
rect 9208 26688 9528 27712
rect 9208 26624 9216 26688
rect 9280 26624 9296 26688
rect 9360 26624 9376 26688
rect 9440 26624 9456 26688
rect 9520 26624 9528 26688
rect 9208 25600 9528 26624
rect 9208 25536 9216 25600
rect 9280 25536 9296 25600
rect 9360 25536 9376 25600
rect 9440 25536 9456 25600
rect 9520 25536 9528 25600
rect 9208 24512 9528 25536
rect 9208 24448 9216 24512
rect 9280 24448 9296 24512
rect 9360 24448 9376 24512
rect 9440 24448 9456 24512
rect 9520 24448 9528 24512
rect 9208 23424 9528 24448
rect 9208 23360 9216 23424
rect 9280 23360 9296 23424
rect 9360 23360 9376 23424
rect 9440 23360 9456 23424
rect 9520 23360 9528 23424
rect 9208 22336 9528 23360
rect 9208 22272 9216 22336
rect 9280 22272 9296 22336
rect 9360 22272 9376 22336
rect 9440 22272 9456 22336
rect 9520 22272 9528 22336
rect 9208 21248 9528 22272
rect 9208 21184 9216 21248
rect 9280 21184 9296 21248
rect 9360 21184 9376 21248
rect 9440 21184 9456 21248
rect 9520 21184 9528 21248
rect 9208 20160 9528 21184
rect 9208 20096 9216 20160
rect 9280 20096 9296 20160
rect 9360 20096 9376 20160
rect 9440 20096 9456 20160
rect 9520 20096 9528 20160
rect 9208 19072 9528 20096
rect 9208 19008 9216 19072
rect 9280 19008 9296 19072
rect 9360 19008 9376 19072
rect 9440 19008 9456 19072
rect 9520 19008 9528 19072
rect 9208 17984 9528 19008
rect 9208 17920 9216 17984
rect 9280 17920 9296 17984
rect 9360 17920 9376 17984
rect 9440 17920 9456 17984
rect 9520 17920 9528 17984
rect 9208 16896 9528 17920
rect 9208 16832 9216 16896
rect 9280 16832 9296 16896
rect 9360 16832 9376 16896
rect 9440 16832 9456 16896
rect 9520 16832 9528 16896
rect 9208 15808 9528 16832
rect 9208 15744 9216 15808
rect 9280 15744 9296 15808
rect 9360 15744 9376 15808
rect 9440 15744 9456 15808
rect 9520 15744 9528 15808
rect 9208 14720 9528 15744
rect 9208 14656 9216 14720
rect 9280 14656 9296 14720
rect 9360 14656 9376 14720
rect 9440 14656 9456 14720
rect 9520 14656 9528 14720
rect 9208 13632 9528 14656
rect 9208 13568 9216 13632
rect 9280 13568 9296 13632
rect 9360 13568 9376 13632
rect 9440 13568 9456 13632
rect 9520 13568 9528 13632
rect 9208 12544 9528 13568
rect 9208 12480 9216 12544
rect 9280 12480 9296 12544
rect 9360 12480 9376 12544
rect 9440 12480 9456 12544
rect 9520 12480 9528 12544
rect 9208 11456 9528 12480
rect 9208 11392 9216 11456
rect 9280 11392 9296 11456
rect 9360 11392 9376 11456
rect 9440 11392 9456 11456
rect 9520 11392 9528 11456
rect 9208 10368 9528 11392
rect 9208 10304 9216 10368
rect 9280 10304 9296 10368
rect 9360 10304 9376 10368
rect 9440 10304 9456 10368
rect 9520 10304 9528 10368
rect 9208 9280 9528 10304
rect 9208 9216 9216 9280
rect 9280 9216 9296 9280
rect 9360 9216 9376 9280
rect 9440 9216 9456 9280
rect 9520 9216 9528 9280
rect 9208 8192 9528 9216
rect 9208 8128 9216 8192
rect 9280 8128 9296 8192
rect 9360 8128 9376 8192
rect 9440 8128 9456 8192
rect 9520 8128 9528 8192
rect 9208 7104 9528 8128
rect 9208 7040 9216 7104
rect 9280 7040 9296 7104
rect 9360 7040 9376 7104
rect 9440 7040 9456 7104
rect 9520 7040 9528 7104
rect 9208 6016 9528 7040
rect 9208 5952 9216 6016
rect 9280 5952 9296 6016
rect 9360 5952 9376 6016
rect 9440 5952 9456 6016
rect 9520 5952 9528 6016
rect 9208 4928 9528 5952
rect 9208 4864 9216 4928
rect 9280 4864 9296 4928
rect 9360 4864 9376 4928
rect 9440 4864 9456 4928
rect 9520 4864 9528 4928
rect 9208 3840 9528 4864
rect 9208 3776 9216 3840
rect 9280 3776 9296 3840
rect 9360 3776 9376 3840
rect 9440 3776 9456 3840
rect 9520 3776 9528 3840
rect 9208 2752 9528 3776
rect 9208 2688 9216 2752
rect 9280 2688 9296 2752
rect 9360 2688 9376 2752
rect 9440 2688 9456 2752
rect 9520 2688 9528 2752
rect 9208 2128 9528 2688
rect 14208 46816 14528 47376
rect 14208 46752 14216 46816
rect 14280 46752 14296 46816
rect 14360 46752 14376 46816
rect 14440 46752 14456 46816
rect 14520 46752 14528 46816
rect 14208 45728 14528 46752
rect 14208 45664 14216 45728
rect 14280 45664 14296 45728
rect 14360 45664 14376 45728
rect 14440 45664 14456 45728
rect 14520 45664 14528 45728
rect 14208 44640 14528 45664
rect 14208 44576 14216 44640
rect 14280 44576 14296 44640
rect 14360 44576 14376 44640
rect 14440 44576 14456 44640
rect 14520 44576 14528 44640
rect 14208 43552 14528 44576
rect 14208 43488 14216 43552
rect 14280 43488 14296 43552
rect 14360 43488 14376 43552
rect 14440 43488 14456 43552
rect 14520 43488 14528 43552
rect 14208 42464 14528 43488
rect 14208 42400 14216 42464
rect 14280 42400 14296 42464
rect 14360 42400 14376 42464
rect 14440 42400 14456 42464
rect 14520 42400 14528 42464
rect 14208 41376 14528 42400
rect 14208 41312 14216 41376
rect 14280 41312 14296 41376
rect 14360 41312 14376 41376
rect 14440 41312 14456 41376
rect 14520 41312 14528 41376
rect 14208 40288 14528 41312
rect 14208 40224 14216 40288
rect 14280 40224 14296 40288
rect 14360 40224 14376 40288
rect 14440 40224 14456 40288
rect 14520 40224 14528 40288
rect 14208 39200 14528 40224
rect 14208 39136 14216 39200
rect 14280 39136 14296 39200
rect 14360 39136 14376 39200
rect 14440 39136 14456 39200
rect 14520 39136 14528 39200
rect 14208 38112 14528 39136
rect 14208 38048 14216 38112
rect 14280 38048 14296 38112
rect 14360 38048 14376 38112
rect 14440 38048 14456 38112
rect 14520 38048 14528 38112
rect 14208 37024 14528 38048
rect 14208 36960 14216 37024
rect 14280 36960 14296 37024
rect 14360 36960 14376 37024
rect 14440 36960 14456 37024
rect 14520 36960 14528 37024
rect 14208 35936 14528 36960
rect 14208 35872 14216 35936
rect 14280 35872 14296 35936
rect 14360 35872 14376 35936
rect 14440 35872 14456 35936
rect 14520 35872 14528 35936
rect 14208 34848 14528 35872
rect 14208 34784 14216 34848
rect 14280 34784 14296 34848
rect 14360 34784 14376 34848
rect 14440 34784 14456 34848
rect 14520 34784 14528 34848
rect 14208 33760 14528 34784
rect 14208 33696 14216 33760
rect 14280 33696 14296 33760
rect 14360 33696 14376 33760
rect 14440 33696 14456 33760
rect 14520 33696 14528 33760
rect 14208 32672 14528 33696
rect 14208 32608 14216 32672
rect 14280 32608 14296 32672
rect 14360 32608 14376 32672
rect 14440 32608 14456 32672
rect 14520 32608 14528 32672
rect 14208 31584 14528 32608
rect 14208 31520 14216 31584
rect 14280 31520 14296 31584
rect 14360 31520 14376 31584
rect 14440 31520 14456 31584
rect 14520 31520 14528 31584
rect 14208 30496 14528 31520
rect 14208 30432 14216 30496
rect 14280 30432 14296 30496
rect 14360 30432 14376 30496
rect 14440 30432 14456 30496
rect 14520 30432 14528 30496
rect 14208 29408 14528 30432
rect 14208 29344 14216 29408
rect 14280 29344 14296 29408
rect 14360 29344 14376 29408
rect 14440 29344 14456 29408
rect 14520 29344 14528 29408
rect 14208 28320 14528 29344
rect 14208 28256 14216 28320
rect 14280 28256 14296 28320
rect 14360 28256 14376 28320
rect 14440 28256 14456 28320
rect 14520 28256 14528 28320
rect 14208 27232 14528 28256
rect 14208 27168 14216 27232
rect 14280 27168 14296 27232
rect 14360 27168 14376 27232
rect 14440 27168 14456 27232
rect 14520 27168 14528 27232
rect 14208 26144 14528 27168
rect 14208 26080 14216 26144
rect 14280 26080 14296 26144
rect 14360 26080 14376 26144
rect 14440 26080 14456 26144
rect 14520 26080 14528 26144
rect 14208 25056 14528 26080
rect 14208 24992 14216 25056
rect 14280 24992 14296 25056
rect 14360 24992 14376 25056
rect 14440 24992 14456 25056
rect 14520 24992 14528 25056
rect 14208 23968 14528 24992
rect 14208 23904 14216 23968
rect 14280 23904 14296 23968
rect 14360 23904 14376 23968
rect 14440 23904 14456 23968
rect 14520 23904 14528 23968
rect 14208 22880 14528 23904
rect 14208 22816 14216 22880
rect 14280 22816 14296 22880
rect 14360 22816 14376 22880
rect 14440 22816 14456 22880
rect 14520 22816 14528 22880
rect 14208 21792 14528 22816
rect 14208 21728 14216 21792
rect 14280 21728 14296 21792
rect 14360 21728 14376 21792
rect 14440 21728 14456 21792
rect 14520 21728 14528 21792
rect 14208 20704 14528 21728
rect 14208 20640 14216 20704
rect 14280 20640 14296 20704
rect 14360 20640 14376 20704
rect 14440 20640 14456 20704
rect 14520 20640 14528 20704
rect 14208 19616 14528 20640
rect 14208 19552 14216 19616
rect 14280 19552 14296 19616
rect 14360 19552 14376 19616
rect 14440 19552 14456 19616
rect 14520 19552 14528 19616
rect 14208 18528 14528 19552
rect 14208 18464 14216 18528
rect 14280 18464 14296 18528
rect 14360 18464 14376 18528
rect 14440 18464 14456 18528
rect 14520 18464 14528 18528
rect 14208 17440 14528 18464
rect 14208 17376 14216 17440
rect 14280 17376 14296 17440
rect 14360 17376 14376 17440
rect 14440 17376 14456 17440
rect 14520 17376 14528 17440
rect 14208 16352 14528 17376
rect 14208 16288 14216 16352
rect 14280 16288 14296 16352
rect 14360 16288 14376 16352
rect 14440 16288 14456 16352
rect 14520 16288 14528 16352
rect 14208 15264 14528 16288
rect 14208 15200 14216 15264
rect 14280 15200 14296 15264
rect 14360 15200 14376 15264
rect 14440 15200 14456 15264
rect 14520 15200 14528 15264
rect 14208 14176 14528 15200
rect 14208 14112 14216 14176
rect 14280 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14528 14176
rect 14208 13088 14528 14112
rect 14208 13024 14216 13088
rect 14280 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14528 13088
rect 14208 12000 14528 13024
rect 14208 11936 14216 12000
rect 14280 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14528 12000
rect 14208 10912 14528 11936
rect 14208 10848 14216 10912
rect 14280 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14528 10912
rect 14208 9824 14528 10848
rect 14208 9760 14216 9824
rect 14280 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14528 9824
rect 14208 8736 14528 9760
rect 14208 8672 14216 8736
rect 14280 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14528 8736
rect 14208 7648 14528 8672
rect 14208 7584 14216 7648
rect 14280 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14528 7648
rect 14208 6560 14528 7584
rect 14208 6496 14216 6560
rect 14280 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14528 6560
rect 14208 5472 14528 6496
rect 14208 5408 14216 5472
rect 14280 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14528 5472
rect 14208 4384 14528 5408
rect 14208 4320 14216 4384
rect 14280 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14528 4384
rect 14208 3296 14528 4320
rect 14208 3232 14216 3296
rect 14280 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14528 3296
rect 14208 2208 14528 3232
rect 14208 2144 14216 2208
rect 14280 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14528 2208
rect 19208 47360 19528 47376
rect 19208 47296 19216 47360
rect 19280 47296 19296 47360
rect 19360 47296 19376 47360
rect 19440 47296 19456 47360
rect 19520 47296 19528 47360
rect 19208 46272 19528 47296
rect 19208 46208 19216 46272
rect 19280 46208 19296 46272
rect 19360 46208 19376 46272
rect 19440 46208 19456 46272
rect 19520 46208 19528 46272
rect 19208 45184 19528 46208
rect 19208 45120 19216 45184
rect 19280 45120 19296 45184
rect 19360 45120 19376 45184
rect 19440 45120 19456 45184
rect 19520 45120 19528 45184
rect 19208 44096 19528 45120
rect 19208 44032 19216 44096
rect 19280 44032 19296 44096
rect 19360 44032 19376 44096
rect 19440 44032 19456 44096
rect 19520 44032 19528 44096
rect 19208 43008 19528 44032
rect 19208 42944 19216 43008
rect 19280 42944 19296 43008
rect 19360 42944 19376 43008
rect 19440 42944 19456 43008
rect 19520 42944 19528 43008
rect 19208 41920 19528 42944
rect 19208 41856 19216 41920
rect 19280 41856 19296 41920
rect 19360 41856 19376 41920
rect 19440 41856 19456 41920
rect 19520 41856 19528 41920
rect 19208 40832 19528 41856
rect 19208 40768 19216 40832
rect 19280 40768 19296 40832
rect 19360 40768 19376 40832
rect 19440 40768 19456 40832
rect 19520 40768 19528 40832
rect 19208 39744 19528 40768
rect 19208 39680 19216 39744
rect 19280 39680 19296 39744
rect 19360 39680 19376 39744
rect 19440 39680 19456 39744
rect 19520 39680 19528 39744
rect 19208 38656 19528 39680
rect 19208 38592 19216 38656
rect 19280 38592 19296 38656
rect 19360 38592 19376 38656
rect 19440 38592 19456 38656
rect 19520 38592 19528 38656
rect 19208 37568 19528 38592
rect 19208 37504 19216 37568
rect 19280 37504 19296 37568
rect 19360 37504 19376 37568
rect 19440 37504 19456 37568
rect 19520 37504 19528 37568
rect 19208 36480 19528 37504
rect 19208 36416 19216 36480
rect 19280 36416 19296 36480
rect 19360 36416 19376 36480
rect 19440 36416 19456 36480
rect 19520 36416 19528 36480
rect 19208 35392 19528 36416
rect 19208 35328 19216 35392
rect 19280 35328 19296 35392
rect 19360 35328 19376 35392
rect 19440 35328 19456 35392
rect 19520 35328 19528 35392
rect 19208 34304 19528 35328
rect 19208 34240 19216 34304
rect 19280 34240 19296 34304
rect 19360 34240 19376 34304
rect 19440 34240 19456 34304
rect 19520 34240 19528 34304
rect 19208 33216 19528 34240
rect 19208 33152 19216 33216
rect 19280 33152 19296 33216
rect 19360 33152 19376 33216
rect 19440 33152 19456 33216
rect 19520 33152 19528 33216
rect 19208 32128 19528 33152
rect 19208 32064 19216 32128
rect 19280 32064 19296 32128
rect 19360 32064 19376 32128
rect 19440 32064 19456 32128
rect 19520 32064 19528 32128
rect 19208 31040 19528 32064
rect 19208 30976 19216 31040
rect 19280 30976 19296 31040
rect 19360 30976 19376 31040
rect 19440 30976 19456 31040
rect 19520 30976 19528 31040
rect 19208 29952 19528 30976
rect 19208 29888 19216 29952
rect 19280 29888 19296 29952
rect 19360 29888 19376 29952
rect 19440 29888 19456 29952
rect 19520 29888 19528 29952
rect 19208 28864 19528 29888
rect 19208 28800 19216 28864
rect 19280 28800 19296 28864
rect 19360 28800 19376 28864
rect 19440 28800 19456 28864
rect 19520 28800 19528 28864
rect 19208 27776 19528 28800
rect 19208 27712 19216 27776
rect 19280 27712 19296 27776
rect 19360 27712 19376 27776
rect 19440 27712 19456 27776
rect 19520 27712 19528 27776
rect 19208 26688 19528 27712
rect 19208 26624 19216 26688
rect 19280 26624 19296 26688
rect 19360 26624 19376 26688
rect 19440 26624 19456 26688
rect 19520 26624 19528 26688
rect 19208 25600 19528 26624
rect 19208 25536 19216 25600
rect 19280 25536 19296 25600
rect 19360 25536 19376 25600
rect 19440 25536 19456 25600
rect 19520 25536 19528 25600
rect 19208 24512 19528 25536
rect 19208 24448 19216 24512
rect 19280 24448 19296 24512
rect 19360 24448 19376 24512
rect 19440 24448 19456 24512
rect 19520 24448 19528 24512
rect 19208 23424 19528 24448
rect 19208 23360 19216 23424
rect 19280 23360 19296 23424
rect 19360 23360 19376 23424
rect 19440 23360 19456 23424
rect 19520 23360 19528 23424
rect 19208 22336 19528 23360
rect 19208 22272 19216 22336
rect 19280 22272 19296 22336
rect 19360 22272 19376 22336
rect 19440 22272 19456 22336
rect 19520 22272 19528 22336
rect 19208 21248 19528 22272
rect 19208 21184 19216 21248
rect 19280 21184 19296 21248
rect 19360 21184 19376 21248
rect 19440 21184 19456 21248
rect 19520 21184 19528 21248
rect 19208 20160 19528 21184
rect 19208 20096 19216 20160
rect 19280 20096 19296 20160
rect 19360 20096 19376 20160
rect 19440 20096 19456 20160
rect 19520 20096 19528 20160
rect 19208 2176 19528 20096
rect 24208 46816 24528 47376
rect 24208 46752 24216 46816
rect 24280 46752 24296 46816
rect 24360 46752 24376 46816
rect 24440 46752 24456 46816
rect 24520 46752 24528 46816
rect 24208 45728 24528 46752
rect 24208 45664 24216 45728
rect 24280 45664 24296 45728
rect 24360 45664 24376 45728
rect 24440 45664 24456 45728
rect 24520 45664 24528 45728
rect 24208 44640 24528 45664
rect 24208 44576 24216 44640
rect 24280 44576 24296 44640
rect 24360 44576 24376 44640
rect 24440 44576 24456 44640
rect 24520 44576 24528 44640
rect 24208 43552 24528 44576
rect 24208 43488 24216 43552
rect 24280 43488 24296 43552
rect 24360 43488 24376 43552
rect 24440 43488 24456 43552
rect 24520 43488 24528 43552
rect 24208 42464 24528 43488
rect 24208 42400 24216 42464
rect 24280 42400 24296 42464
rect 24360 42400 24376 42464
rect 24440 42400 24456 42464
rect 24520 42400 24528 42464
rect 24208 41376 24528 42400
rect 24208 41312 24216 41376
rect 24280 41312 24296 41376
rect 24360 41312 24376 41376
rect 24440 41312 24456 41376
rect 24520 41312 24528 41376
rect 24208 40288 24528 41312
rect 24208 40224 24216 40288
rect 24280 40224 24296 40288
rect 24360 40224 24376 40288
rect 24440 40224 24456 40288
rect 24520 40224 24528 40288
rect 24208 39200 24528 40224
rect 24208 39136 24216 39200
rect 24280 39136 24296 39200
rect 24360 39136 24376 39200
rect 24440 39136 24456 39200
rect 24520 39136 24528 39200
rect 24208 38112 24528 39136
rect 24208 38048 24216 38112
rect 24280 38048 24296 38112
rect 24360 38048 24376 38112
rect 24440 38048 24456 38112
rect 24520 38048 24528 38112
rect 24208 37024 24528 38048
rect 24208 36960 24216 37024
rect 24280 36960 24296 37024
rect 24360 36960 24376 37024
rect 24440 36960 24456 37024
rect 24520 36960 24528 37024
rect 24208 35936 24528 36960
rect 24208 35872 24216 35936
rect 24280 35872 24296 35936
rect 24360 35872 24376 35936
rect 24440 35872 24456 35936
rect 24520 35872 24528 35936
rect 24208 34848 24528 35872
rect 24208 34784 24216 34848
rect 24280 34784 24296 34848
rect 24360 34784 24376 34848
rect 24440 34784 24456 34848
rect 24520 34784 24528 34848
rect 24208 33760 24528 34784
rect 24208 33696 24216 33760
rect 24280 33696 24296 33760
rect 24360 33696 24376 33760
rect 24440 33696 24456 33760
rect 24520 33696 24528 33760
rect 24208 32672 24528 33696
rect 24208 32608 24216 32672
rect 24280 32608 24296 32672
rect 24360 32608 24376 32672
rect 24440 32608 24456 32672
rect 24520 32608 24528 32672
rect 24208 31584 24528 32608
rect 24208 31520 24216 31584
rect 24280 31520 24296 31584
rect 24360 31520 24376 31584
rect 24440 31520 24456 31584
rect 24520 31520 24528 31584
rect 24208 30496 24528 31520
rect 24208 30432 24216 30496
rect 24280 30432 24296 30496
rect 24360 30432 24376 30496
rect 24440 30432 24456 30496
rect 24520 30432 24528 30496
rect 24208 29408 24528 30432
rect 24208 29344 24216 29408
rect 24280 29344 24296 29408
rect 24360 29344 24376 29408
rect 24440 29344 24456 29408
rect 24520 29344 24528 29408
rect 24208 28320 24528 29344
rect 24208 28256 24216 28320
rect 24280 28256 24296 28320
rect 24360 28256 24376 28320
rect 24440 28256 24456 28320
rect 24520 28256 24528 28320
rect 24208 27232 24528 28256
rect 24208 27168 24216 27232
rect 24280 27168 24296 27232
rect 24360 27168 24376 27232
rect 24440 27168 24456 27232
rect 24520 27168 24528 27232
rect 24208 26144 24528 27168
rect 24208 26080 24216 26144
rect 24280 26080 24296 26144
rect 24360 26080 24376 26144
rect 24440 26080 24456 26144
rect 24520 26080 24528 26144
rect 24208 25056 24528 26080
rect 24208 24992 24216 25056
rect 24280 24992 24296 25056
rect 24360 24992 24376 25056
rect 24440 24992 24456 25056
rect 24520 24992 24528 25056
rect 24208 23968 24528 24992
rect 24208 23904 24216 23968
rect 24280 23904 24296 23968
rect 24360 23904 24376 23968
rect 24440 23904 24456 23968
rect 24520 23904 24528 23968
rect 24208 22880 24528 23904
rect 24208 22816 24216 22880
rect 24280 22816 24296 22880
rect 24360 22816 24376 22880
rect 24440 22816 24456 22880
rect 24520 22816 24528 22880
rect 24208 21792 24528 22816
rect 24208 21728 24216 21792
rect 24280 21728 24296 21792
rect 24360 21728 24376 21792
rect 24440 21728 24456 21792
rect 24520 21728 24528 21792
rect 24208 20704 24528 21728
rect 24208 20640 24216 20704
rect 24280 20640 24296 20704
rect 24360 20640 24376 20704
rect 24440 20640 24456 20704
rect 24520 20640 24528 20704
rect 24208 19616 24528 20640
rect 24208 19552 24216 19616
rect 24280 19552 24296 19616
rect 24360 19552 24376 19616
rect 24440 19552 24456 19616
rect 24520 19552 24528 19616
rect 24208 15638 24528 19552
rect 24208 15254 24216 15638
rect 24520 15254 24528 15638
rect 24208 11907 24528 15254
rect 24208 11603 24216 11907
rect 24520 11603 24528 11907
rect 24208 9358 24528 11603
rect 24208 9054 24216 9358
rect 24520 9054 24528 9358
rect 24208 6809 24528 9054
rect 24208 6505 24216 6809
rect 24520 6505 24528 6809
rect 24208 3222 24528 6505
rect 24208 2838 24216 3222
rect 24520 2838 24528 3222
rect 24208 2176 24528 2838
rect 29208 47360 29528 47376
rect 29208 47296 29216 47360
rect 29280 47296 29296 47360
rect 29360 47296 29376 47360
rect 29440 47296 29456 47360
rect 29520 47296 29528 47360
rect 29208 46272 29528 47296
rect 29208 46208 29216 46272
rect 29280 46208 29296 46272
rect 29360 46208 29376 46272
rect 29440 46208 29456 46272
rect 29520 46208 29528 46272
rect 29208 45184 29528 46208
rect 29208 45120 29216 45184
rect 29280 45120 29296 45184
rect 29360 45120 29376 45184
rect 29440 45120 29456 45184
rect 29520 45120 29528 45184
rect 29208 44096 29528 45120
rect 29208 44032 29216 44096
rect 29280 44032 29296 44096
rect 29360 44032 29376 44096
rect 29440 44032 29456 44096
rect 29520 44032 29528 44096
rect 29208 43008 29528 44032
rect 29208 42944 29216 43008
rect 29280 42944 29296 43008
rect 29360 42944 29376 43008
rect 29440 42944 29456 43008
rect 29520 42944 29528 43008
rect 29208 41920 29528 42944
rect 29208 41856 29216 41920
rect 29280 41856 29296 41920
rect 29360 41856 29376 41920
rect 29440 41856 29456 41920
rect 29520 41856 29528 41920
rect 29208 40832 29528 41856
rect 29208 40768 29216 40832
rect 29280 40768 29296 40832
rect 29360 40768 29376 40832
rect 29440 40768 29456 40832
rect 29520 40768 29528 40832
rect 29208 39744 29528 40768
rect 29208 39680 29216 39744
rect 29280 39680 29296 39744
rect 29360 39680 29376 39744
rect 29440 39680 29456 39744
rect 29520 39680 29528 39744
rect 29208 38656 29528 39680
rect 29208 38592 29216 38656
rect 29280 38592 29296 38656
rect 29360 38592 29376 38656
rect 29440 38592 29456 38656
rect 29520 38592 29528 38656
rect 29208 37568 29528 38592
rect 29208 37504 29216 37568
rect 29280 37504 29296 37568
rect 29360 37504 29376 37568
rect 29440 37504 29456 37568
rect 29520 37504 29528 37568
rect 29208 36480 29528 37504
rect 29208 36416 29216 36480
rect 29280 36416 29296 36480
rect 29360 36416 29376 36480
rect 29440 36416 29456 36480
rect 29520 36416 29528 36480
rect 29208 35392 29528 36416
rect 29208 35328 29216 35392
rect 29280 35328 29296 35392
rect 29360 35328 29376 35392
rect 29440 35328 29456 35392
rect 29520 35328 29528 35392
rect 29208 34304 29528 35328
rect 29208 34240 29216 34304
rect 29280 34240 29296 34304
rect 29360 34240 29376 34304
rect 29440 34240 29456 34304
rect 29520 34240 29528 34304
rect 29208 33216 29528 34240
rect 29208 33152 29216 33216
rect 29280 33152 29296 33216
rect 29360 33152 29376 33216
rect 29440 33152 29456 33216
rect 29520 33152 29528 33216
rect 29208 32128 29528 33152
rect 29208 32064 29216 32128
rect 29280 32064 29296 32128
rect 29360 32064 29376 32128
rect 29440 32064 29456 32128
rect 29520 32064 29528 32128
rect 29208 31040 29528 32064
rect 29208 30976 29216 31040
rect 29280 30976 29296 31040
rect 29360 30976 29376 31040
rect 29440 30976 29456 31040
rect 29520 30976 29528 31040
rect 29208 29952 29528 30976
rect 29208 29888 29216 29952
rect 29280 29888 29296 29952
rect 29360 29888 29376 29952
rect 29440 29888 29456 29952
rect 29520 29888 29528 29952
rect 29208 28864 29528 29888
rect 29208 28800 29216 28864
rect 29280 28800 29296 28864
rect 29360 28800 29376 28864
rect 29440 28800 29456 28864
rect 29520 28800 29528 28864
rect 29208 27776 29528 28800
rect 29208 27712 29216 27776
rect 29280 27712 29296 27776
rect 29360 27712 29376 27776
rect 29440 27712 29456 27776
rect 29520 27712 29528 27776
rect 29208 26688 29528 27712
rect 29208 26624 29216 26688
rect 29280 26624 29296 26688
rect 29360 26624 29376 26688
rect 29440 26624 29456 26688
rect 29520 26624 29528 26688
rect 29208 25600 29528 26624
rect 29208 25536 29216 25600
rect 29280 25536 29296 25600
rect 29360 25536 29376 25600
rect 29440 25536 29456 25600
rect 29520 25536 29528 25600
rect 29208 24512 29528 25536
rect 29208 24448 29216 24512
rect 29280 24448 29296 24512
rect 29360 24448 29376 24512
rect 29440 24448 29456 24512
rect 29520 24448 29528 24512
rect 29208 23424 29528 24448
rect 29208 23360 29216 23424
rect 29280 23360 29296 23424
rect 29360 23360 29376 23424
rect 29440 23360 29456 23424
rect 29520 23360 29528 23424
rect 29208 22336 29528 23360
rect 29208 22272 29216 22336
rect 29280 22272 29296 22336
rect 29360 22272 29376 22336
rect 29440 22272 29456 22336
rect 29520 22272 29528 22336
rect 29208 21248 29528 22272
rect 29208 21184 29216 21248
rect 29280 21184 29296 21248
rect 29360 21184 29376 21248
rect 29440 21184 29456 21248
rect 29520 21184 29528 21248
rect 29208 20160 29528 21184
rect 29208 20096 29216 20160
rect 29280 20096 29296 20160
rect 29360 20096 29376 20160
rect 29440 20096 29456 20160
rect 29520 20096 29528 20160
rect 29208 16438 29528 20096
rect 29208 16054 29216 16438
rect 29520 16054 29528 16438
rect 29208 10633 29528 16054
rect 29208 10329 29216 10633
rect 29520 10329 29528 10633
rect 29208 8083 29528 10329
rect 29208 7779 29216 8083
rect 29520 7779 29528 8083
rect 29208 2430 29528 7779
rect 29208 2206 29216 2430
rect 29520 2206 29528 2430
rect 29208 2176 29528 2206
rect 34208 46816 34528 47376
rect 34208 46752 34216 46816
rect 34280 46752 34296 46816
rect 34360 46752 34376 46816
rect 34440 46752 34456 46816
rect 34520 46752 34528 46816
rect 34208 45728 34528 46752
rect 34208 45664 34216 45728
rect 34280 45664 34296 45728
rect 34360 45664 34376 45728
rect 34440 45664 34456 45728
rect 34520 45664 34528 45728
rect 34208 44640 34528 45664
rect 34208 44576 34216 44640
rect 34280 44576 34296 44640
rect 34360 44576 34376 44640
rect 34440 44576 34456 44640
rect 34520 44576 34528 44640
rect 34208 43552 34528 44576
rect 34208 43488 34216 43552
rect 34280 43488 34296 43552
rect 34360 43488 34376 43552
rect 34440 43488 34456 43552
rect 34520 43488 34528 43552
rect 34208 42464 34528 43488
rect 34208 42400 34216 42464
rect 34280 42400 34296 42464
rect 34360 42400 34376 42464
rect 34440 42400 34456 42464
rect 34520 42400 34528 42464
rect 34208 41376 34528 42400
rect 34208 41312 34216 41376
rect 34280 41312 34296 41376
rect 34360 41312 34376 41376
rect 34440 41312 34456 41376
rect 34520 41312 34528 41376
rect 34208 40288 34528 41312
rect 34208 40224 34216 40288
rect 34280 40224 34296 40288
rect 34360 40224 34376 40288
rect 34440 40224 34456 40288
rect 34520 40224 34528 40288
rect 34208 39200 34528 40224
rect 34208 39136 34216 39200
rect 34280 39136 34296 39200
rect 34360 39136 34376 39200
rect 34440 39136 34456 39200
rect 34520 39136 34528 39200
rect 34208 38112 34528 39136
rect 34208 38048 34216 38112
rect 34280 38048 34296 38112
rect 34360 38048 34376 38112
rect 34440 38048 34456 38112
rect 34520 38048 34528 38112
rect 34208 37024 34528 38048
rect 34208 36960 34216 37024
rect 34280 36960 34296 37024
rect 34360 36960 34376 37024
rect 34440 36960 34456 37024
rect 34520 36960 34528 37024
rect 34208 35936 34528 36960
rect 34208 35872 34216 35936
rect 34280 35872 34296 35936
rect 34360 35872 34376 35936
rect 34440 35872 34456 35936
rect 34520 35872 34528 35936
rect 34208 34848 34528 35872
rect 34208 34784 34216 34848
rect 34280 34784 34296 34848
rect 34360 34784 34376 34848
rect 34440 34784 34456 34848
rect 34520 34784 34528 34848
rect 34208 33760 34528 34784
rect 34208 33696 34216 33760
rect 34280 33696 34296 33760
rect 34360 33696 34376 33760
rect 34440 33696 34456 33760
rect 34520 33696 34528 33760
rect 34208 32672 34528 33696
rect 34208 32608 34216 32672
rect 34280 32608 34296 32672
rect 34360 32608 34376 32672
rect 34440 32608 34456 32672
rect 34520 32608 34528 32672
rect 34208 31584 34528 32608
rect 34208 31520 34216 31584
rect 34280 31520 34296 31584
rect 34360 31520 34376 31584
rect 34440 31520 34456 31584
rect 34520 31520 34528 31584
rect 34208 30496 34528 31520
rect 34208 30432 34216 30496
rect 34280 30432 34296 30496
rect 34360 30432 34376 30496
rect 34440 30432 34456 30496
rect 34520 30432 34528 30496
rect 34208 29408 34528 30432
rect 34208 29344 34216 29408
rect 34280 29344 34296 29408
rect 34360 29344 34376 29408
rect 34440 29344 34456 29408
rect 34520 29344 34528 29408
rect 34208 28320 34528 29344
rect 34208 28256 34216 28320
rect 34280 28256 34296 28320
rect 34360 28256 34376 28320
rect 34440 28256 34456 28320
rect 34520 28256 34528 28320
rect 34208 27232 34528 28256
rect 34208 27168 34216 27232
rect 34280 27168 34296 27232
rect 34360 27168 34376 27232
rect 34440 27168 34456 27232
rect 34520 27168 34528 27232
rect 34208 26144 34528 27168
rect 34208 26080 34216 26144
rect 34280 26080 34296 26144
rect 34360 26080 34376 26144
rect 34440 26080 34456 26144
rect 34520 26080 34528 26144
rect 34208 25056 34528 26080
rect 34208 24992 34216 25056
rect 34280 24992 34296 25056
rect 34360 24992 34376 25056
rect 34440 24992 34456 25056
rect 34520 24992 34528 25056
rect 34208 23968 34528 24992
rect 34208 23904 34216 23968
rect 34280 23904 34296 23968
rect 34360 23904 34376 23968
rect 34440 23904 34456 23968
rect 34520 23904 34528 23968
rect 34208 22880 34528 23904
rect 34208 22816 34216 22880
rect 34280 22816 34296 22880
rect 34360 22816 34376 22880
rect 34440 22816 34456 22880
rect 34520 22816 34528 22880
rect 34208 21792 34528 22816
rect 34208 21728 34216 21792
rect 34280 21728 34296 21792
rect 34360 21728 34376 21792
rect 34440 21728 34456 21792
rect 34520 21728 34528 21792
rect 34208 20704 34528 21728
rect 34208 20640 34216 20704
rect 34280 20640 34296 20704
rect 34360 20640 34376 20704
rect 34440 20640 34456 20704
rect 34520 20640 34528 20704
rect 34208 19616 34528 20640
rect 34208 19552 34216 19616
rect 34280 19552 34296 19616
rect 34360 19552 34376 19616
rect 34440 19552 34456 19616
rect 34520 19552 34528 19616
rect 34208 11907 34528 19552
rect 34208 11603 34216 11907
rect 34520 11603 34528 11907
rect 34208 9358 34528 11603
rect 34208 9054 34216 9358
rect 34520 9054 34528 9358
rect 34208 6809 34528 9054
rect 34208 6505 34216 6809
rect 34520 6505 34528 6809
rect 34208 2176 34528 6505
rect 39208 47360 39528 47376
rect 39208 47296 39216 47360
rect 39280 47296 39296 47360
rect 39360 47296 39376 47360
rect 39440 47296 39456 47360
rect 39520 47296 39528 47360
rect 39208 46272 39528 47296
rect 39208 46208 39216 46272
rect 39280 46208 39296 46272
rect 39360 46208 39376 46272
rect 39440 46208 39456 46272
rect 39520 46208 39528 46272
rect 39208 45184 39528 46208
rect 39208 45120 39216 45184
rect 39280 45120 39296 45184
rect 39360 45120 39376 45184
rect 39440 45120 39456 45184
rect 39520 45120 39528 45184
rect 39208 44096 39528 45120
rect 39208 44032 39216 44096
rect 39280 44032 39296 44096
rect 39360 44032 39376 44096
rect 39440 44032 39456 44096
rect 39520 44032 39528 44096
rect 39208 43008 39528 44032
rect 39208 42944 39216 43008
rect 39280 42944 39296 43008
rect 39360 42944 39376 43008
rect 39440 42944 39456 43008
rect 39520 42944 39528 43008
rect 39208 41920 39528 42944
rect 39208 41856 39216 41920
rect 39280 41856 39296 41920
rect 39360 41856 39376 41920
rect 39440 41856 39456 41920
rect 39520 41856 39528 41920
rect 39208 40832 39528 41856
rect 39208 40768 39216 40832
rect 39280 40768 39296 40832
rect 39360 40768 39376 40832
rect 39440 40768 39456 40832
rect 39520 40768 39528 40832
rect 39208 39744 39528 40768
rect 39208 39680 39216 39744
rect 39280 39680 39296 39744
rect 39360 39680 39376 39744
rect 39440 39680 39456 39744
rect 39520 39680 39528 39744
rect 39208 38656 39528 39680
rect 39208 38592 39216 38656
rect 39280 38592 39296 38656
rect 39360 38592 39376 38656
rect 39440 38592 39456 38656
rect 39520 38592 39528 38656
rect 39208 37568 39528 38592
rect 39208 37504 39216 37568
rect 39280 37504 39296 37568
rect 39360 37504 39376 37568
rect 39440 37504 39456 37568
rect 39520 37504 39528 37568
rect 39208 36480 39528 37504
rect 39208 36416 39216 36480
rect 39280 36416 39296 36480
rect 39360 36416 39376 36480
rect 39440 36416 39456 36480
rect 39520 36416 39528 36480
rect 39208 35392 39528 36416
rect 39208 35328 39216 35392
rect 39280 35328 39296 35392
rect 39360 35328 39376 35392
rect 39440 35328 39456 35392
rect 39520 35328 39528 35392
rect 39208 34304 39528 35328
rect 39208 34240 39216 34304
rect 39280 34240 39296 34304
rect 39360 34240 39376 34304
rect 39440 34240 39456 34304
rect 39520 34240 39528 34304
rect 39208 33216 39528 34240
rect 39208 33152 39216 33216
rect 39280 33152 39296 33216
rect 39360 33152 39376 33216
rect 39440 33152 39456 33216
rect 39520 33152 39528 33216
rect 39208 32128 39528 33152
rect 39208 32064 39216 32128
rect 39280 32064 39296 32128
rect 39360 32064 39376 32128
rect 39440 32064 39456 32128
rect 39520 32064 39528 32128
rect 39208 31040 39528 32064
rect 39208 30976 39216 31040
rect 39280 30976 39296 31040
rect 39360 30976 39376 31040
rect 39440 30976 39456 31040
rect 39520 30976 39528 31040
rect 39208 29952 39528 30976
rect 39208 29888 39216 29952
rect 39280 29888 39296 29952
rect 39360 29888 39376 29952
rect 39440 29888 39456 29952
rect 39520 29888 39528 29952
rect 39208 28864 39528 29888
rect 39208 28800 39216 28864
rect 39280 28800 39296 28864
rect 39360 28800 39376 28864
rect 39440 28800 39456 28864
rect 39520 28800 39528 28864
rect 39208 27776 39528 28800
rect 39208 27712 39216 27776
rect 39280 27712 39296 27776
rect 39360 27712 39376 27776
rect 39440 27712 39456 27776
rect 39520 27712 39528 27776
rect 39208 26688 39528 27712
rect 39208 26624 39216 26688
rect 39280 26624 39296 26688
rect 39360 26624 39376 26688
rect 39440 26624 39456 26688
rect 39520 26624 39528 26688
rect 39208 25600 39528 26624
rect 39208 25536 39216 25600
rect 39280 25536 39296 25600
rect 39360 25536 39376 25600
rect 39440 25536 39456 25600
rect 39520 25536 39528 25600
rect 39208 24512 39528 25536
rect 39208 24448 39216 24512
rect 39280 24448 39296 24512
rect 39360 24448 39376 24512
rect 39440 24448 39456 24512
rect 39520 24448 39528 24512
rect 39208 23424 39528 24448
rect 39208 23360 39216 23424
rect 39280 23360 39296 23424
rect 39360 23360 39376 23424
rect 39440 23360 39456 23424
rect 39520 23360 39528 23424
rect 39208 22336 39528 23360
rect 39208 22272 39216 22336
rect 39280 22272 39296 22336
rect 39360 22272 39376 22336
rect 39440 22272 39456 22336
rect 39520 22272 39528 22336
rect 39208 21248 39528 22272
rect 39208 21184 39216 21248
rect 39280 21184 39296 21248
rect 39360 21184 39376 21248
rect 39440 21184 39456 21248
rect 39520 21184 39528 21248
rect 39208 20160 39528 21184
rect 39208 20096 39216 20160
rect 39280 20096 39296 20160
rect 39360 20096 39376 20160
rect 39440 20096 39456 20160
rect 39520 20096 39528 20160
rect 39208 19072 39528 20096
rect 39208 19008 39216 19072
rect 39280 19008 39296 19072
rect 39360 19008 39376 19072
rect 39440 19008 39456 19072
rect 39520 19008 39528 19072
rect 39208 17984 39528 19008
rect 39208 17920 39216 17984
rect 39280 17920 39296 17984
rect 39360 17920 39376 17984
rect 39440 17920 39456 17984
rect 39520 17920 39528 17984
rect 39208 16896 39528 17920
rect 39208 16832 39216 16896
rect 39280 16832 39296 16896
rect 39360 16832 39376 16896
rect 39440 16832 39456 16896
rect 39520 16832 39528 16896
rect 39208 15808 39528 16832
rect 39208 15744 39216 15808
rect 39280 15744 39296 15808
rect 39360 15744 39376 15808
rect 39440 15744 39456 15808
rect 39520 15744 39528 15808
rect 39208 14720 39528 15744
rect 39208 14656 39216 14720
rect 39280 14656 39296 14720
rect 39360 14656 39376 14720
rect 39440 14656 39456 14720
rect 39520 14656 39528 14720
rect 39208 13632 39528 14656
rect 39208 13568 39216 13632
rect 39280 13568 39296 13632
rect 39360 13568 39376 13632
rect 39440 13568 39456 13632
rect 39520 13568 39528 13632
rect 39208 12544 39528 13568
rect 39208 12480 39216 12544
rect 39280 12480 39296 12544
rect 39360 12480 39376 12544
rect 39440 12480 39456 12544
rect 39520 12480 39528 12544
rect 39208 11456 39528 12480
rect 39208 11392 39216 11456
rect 39280 11392 39296 11456
rect 39360 11392 39376 11456
rect 39440 11392 39456 11456
rect 39520 11392 39528 11456
rect 39208 10368 39528 11392
rect 39208 10304 39216 10368
rect 39280 10304 39296 10368
rect 39360 10304 39376 10368
rect 39440 10304 39456 10368
rect 39520 10304 39528 10368
rect 39208 9280 39528 10304
rect 39208 9216 39216 9280
rect 39280 9216 39296 9280
rect 39360 9216 39376 9280
rect 39440 9216 39456 9280
rect 39520 9216 39528 9280
rect 39208 8192 39528 9216
rect 39208 8128 39216 8192
rect 39280 8128 39296 8192
rect 39360 8128 39376 8192
rect 39440 8128 39456 8192
rect 39520 8128 39528 8192
rect 39208 7104 39528 8128
rect 39208 7040 39216 7104
rect 39280 7040 39296 7104
rect 39360 7040 39376 7104
rect 39440 7040 39456 7104
rect 39520 7040 39528 7104
rect 39208 6016 39528 7040
rect 39208 5952 39216 6016
rect 39280 5952 39296 6016
rect 39360 5952 39376 6016
rect 39440 5952 39456 6016
rect 39520 5952 39528 6016
rect 39208 4928 39528 5952
rect 39208 4864 39216 4928
rect 39280 4864 39296 4928
rect 39360 4864 39376 4928
rect 39440 4864 39456 4928
rect 39520 4864 39528 4928
rect 39208 3840 39528 4864
rect 39208 3776 39216 3840
rect 39280 3776 39296 3840
rect 39360 3776 39376 3840
rect 39440 3776 39456 3840
rect 39520 3776 39528 3840
rect 39208 2752 39528 3776
rect 39208 2688 39216 2752
rect 39280 2688 39296 2752
rect 39360 2688 39376 2752
rect 39440 2688 39456 2752
rect 39520 2688 39528 2752
rect 14208 2128 14528 2144
rect 39208 2128 39528 2688
rect 44208 46816 44528 47376
rect 44208 46752 44216 46816
rect 44280 46752 44296 46816
rect 44360 46752 44376 46816
rect 44440 46752 44456 46816
rect 44520 46752 44528 46816
rect 44208 45728 44528 46752
rect 44208 45664 44216 45728
rect 44280 45664 44296 45728
rect 44360 45664 44376 45728
rect 44440 45664 44456 45728
rect 44520 45664 44528 45728
rect 44208 44640 44528 45664
rect 44208 44576 44216 44640
rect 44280 44576 44296 44640
rect 44360 44576 44376 44640
rect 44440 44576 44456 44640
rect 44520 44576 44528 44640
rect 44208 43552 44528 44576
rect 44208 43488 44216 43552
rect 44280 43488 44296 43552
rect 44360 43488 44376 43552
rect 44440 43488 44456 43552
rect 44520 43488 44528 43552
rect 44208 42464 44528 43488
rect 44208 42400 44216 42464
rect 44280 42400 44296 42464
rect 44360 42400 44376 42464
rect 44440 42400 44456 42464
rect 44520 42400 44528 42464
rect 44208 41376 44528 42400
rect 44208 41312 44216 41376
rect 44280 41312 44296 41376
rect 44360 41312 44376 41376
rect 44440 41312 44456 41376
rect 44520 41312 44528 41376
rect 44208 40288 44528 41312
rect 44208 40224 44216 40288
rect 44280 40224 44296 40288
rect 44360 40224 44376 40288
rect 44440 40224 44456 40288
rect 44520 40224 44528 40288
rect 44208 39200 44528 40224
rect 44208 39136 44216 39200
rect 44280 39136 44296 39200
rect 44360 39136 44376 39200
rect 44440 39136 44456 39200
rect 44520 39136 44528 39200
rect 44208 38112 44528 39136
rect 44208 38048 44216 38112
rect 44280 38048 44296 38112
rect 44360 38048 44376 38112
rect 44440 38048 44456 38112
rect 44520 38048 44528 38112
rect 44208 37024 44528 38048
rect 44208 36960 44216 37024
rect 44280 36960 44296 37024
rect 44360 36960 44376 37024
rect 44440 36960 44456 37024
rect 44520 36960 44528 37024
rect 44208 35936 44528 36960
rect 44208 35872 44216 35936
rect 44280 35872 44296 35936
rect 44360 35872 44376 35936
rect 44440 35872 44456 35936
rect 44520 35872 44528 35936
rect 44208 34848 44528 35872
rect 44208 34784 44216 34848
rect 44280 34784 44296 34848
rect 44360 34784 44376 34848
rect 44440 34784 44456 34848
rect 44520 34784 44528 34848
rect 44208 33760 44528 34784
rect 44208 33696 44216 33760
rect 44280 33696 44296 33760
rect 44360 33696 44376 33760
rect 44440 33696 44456 33760
rect 44520 33696 44528 33760
rect 44208 32672 44528 33696
rect 44208 32608 44216 32672
rect 44280 32608 44296 32672
rect 44360 32608 44376 32672
rect 44440 32608 44456 32672
rect 44520 32608 44528 32672
rect 44208 31584 44528 32608
rect 44208 31520 44216 31584
rect 44280 31520 44296 31584
rect 44360 31520 44376 31584
rect 44440 31520 44456 31584
rect 44520 31520 44528 31584
rect 44208 30496 44528 31520
rect 44208 30432 44216 30496
rect 44280 30432 44296 30496
rect 44360 30432 44376 30496
rect 44440 30432 44456 30496
rect 44520 30432 44528 30496
rect 44208 29408 44528 30432
rect 44208 29344 44216 29408
rect 44280 29344 44296 29408
rect 44360 29344 44376 29408
rect 44440 29344 44456 29408
rect 44520 29344 44528 29408
rect 44208 28320 44528 29344
rect 44208 28256 44216 28320
rect 44280 28256 44296 28320
rect 44360 28256 44376 28320
rect 44440 28256 44456 28320
rect 44520 28256 44528 28320
rect 44208 27232 44528 28256
rect 44208 27168 44216 27232
rect 44280 27168 44296 27232
rect 44360 27168 44376 27232
rect 44440 27168 44456 27232
rect 44520 27168 44528 27232
rect 44208 26144 44528 27168
rect 44208 26080 44216 26144
rect 44280 26080 44296 26144
rect 44360 26080 44376 26144
rect 44440 26080 44456 26144
rect 44520 26080 44528 26144
rect 44208 25056 44528 26080
rect 44208 24992 44216 25056
rect 44280 24992 44296 25056
rect 44360 24992 44376 25056
rect 44440 24992 44456 25056
rect 44520 24992 44528 25056
rect 44208 23968 44528 24992
rect 44208 23904 44216 23968
rect 44280 23904 44296 23968
rect 44360 23904 44376 23968
rect 44440 23904 44456 23968
rect 44520 23904 44528 23968
rect 44208 22880 44528 23904
rect 44208 22816 44216 22880
rect 44280 22816 44296 22880
rect 44360 22816 44376 22880
rect 44440 22816 44456 22880
rect 44520 22816 44528 22880
rect 44208 21792 44528 22816
rect 44208 21728 44216 21792
rect 44280 21728 44296 21792
rect 44360 21728 44376 21792
rect 44440 21728 44456 21792
rect 44520 21728 44528 21792
rect 44208 20704 44528 21728
rect 44208 20640 44216 20704
rect 44280 20640 44296 20704
rect 44360 20640 44376 20704
rect 44440 20640 44456 20704
rect 44520 20640 44528 20704
rect 44208 19616 44528 20640
rect 44208 19552 44216 19616
rect 44280 19552 44296 19616
rect 44360 19552 44376 19616
rect 44440 19552 44456 19616
rect 44520 19552 44528 19616
rect 44208 18528 44528 19552
rect 44208 18464 44216 18528
rect 44280 18464 44296 18528
rect 44360 18464 44376 18528
rect 44440 18464 44456 18528
rect 44520 18464 44528 18528
rect 44208 17440 44528 18464
rect 44208 17376 44216 17440
rect 44280 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44528 17440
rect 44208 16352 44528 17376
rect 44208 16288 44216 16352
rect 44280 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44528 16352
rect 44208 15264 44528 16288
rect 44208 15200 44216 15264
rect 44280 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44528 15264
rect 44208 14176 44528 15200
rect 44208 14112 44216 14176
rect 44280 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44528 14176
rect 44208 13088 44528 14112
rect 44208 13024 44216 13088
rect 44280 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44528 13088
rect 44208 12000 44528 13024
rect 44208 11936 44216 12000
rect 44280 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44528 12000
rect 44208 10912 44528 11936
rect 44208 10848 44216 10912
rect 44280 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44528 10912
rect 44208 9824 44528 10848
rect 44208 9760 44216 9824
rect 44280 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44528 9824
rect 44208 8736 44528 9760
rect 44208 8672 44216 8736
rect 44280 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44528 8736
rect 44208 7648 44528 8672
rect 44208 7584 44216 7648
rect 44280 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44528 7648
rect 44208 6560 44528 7584
rect 44208 6496 44216 6560
rect 44280 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44528 6560
rect 44208 5472 44528 6496
rect 44208 5408 44216 5472
rect 44280 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44528 5472
rect 44208 4384 44528 5408
rect 44208 4320 44216 4384
rect 44280 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44528 4384
rect 44208 3296 44528 4320
rect 44208 3232 44216 3296
rect 44280 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44528 3296
rect 44208 2208 44528 3232
rect 44208 2144 44216 2208
rect 44280 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44528 2208
rect 44208 2128 44528 2144
use sky130_fd_sc_hd__decap_12  FILLER_6_496
timestamp 1626105910
transform 1 0 46736 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_508
timestamp 1626105910
transform 1 0 47840 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_484
timestamp 1626105910
transform 1 0 45632 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1626105910
transform 1 0 45540 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_475
timestamp 1626105910
transform 1 0 44804 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_463
timestamp 1626105910
transform 1 0 43700 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_478
timestamp 1626105910
transform 1 0 45080 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_478
timestamp 1626105910
transform 1 0 45080 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__D
timestamp 1626105910
transform -1 0 45632 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1626105910
transform 1 0 48300 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_482
timestamp 1626105910
transform 1 0 45448 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _109_
timestamp 1626105910
transform -1 0 45080 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1626105910
transform -1 0 48852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1626105910
transform 1 0 48116 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1626105910
transform 1 0 48208 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_491
timestamp 1626105910
transform 1 0 46276 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_503
timestamp 1626105910
transform 1 0 47380 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_479
timestamp 1626105910
transform 1 0 45172 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_467
timestamp 1626105910
transform 1 0 44068 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_455
timestamp 1626105910
transform 1 0 42964 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_509
timestamp 1626105910
transform 1 0 47932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__CLK
timestamp 1626105910
transform -1 0 43332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_467
timestamp 1626105910
transform 1 0 44068 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_461
timestamp 1626105910
transform 1 0 43516 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1626105910
transform 1 0 42964 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_455
timestamp 1626105910
transform 1 0 42964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A3
timestamp 1626105910
transform 1 0 43332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1626105910
transform -1 0 48852 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_496
timestamp 1626105910
transform 1 0 46736 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_508
timestamp 1626105910
transform 1 0 47840 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_484
timestamp 1626105910
transform 1 0 45632 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1626105910
transform 1 0 45540 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_475
timestamp 1626105910
transform 1 0 44804 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_463
timestamp 1626105910
transform 1 0 43700 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A2
timestamp 1626105910
transform 1 0 43884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_497
timestamp 1626105910
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_485
timestamp 1626105910
transform 1 0 45724 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_471
timestamp 1626105910
transform 1 0 44436 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1626105910
transform 1 0 45632 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1626105910
transform -1 0 48852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1626105910
transform 1 0 48116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1626105910
transform 1 0 48208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1626105910
transform -1 0 48852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1626105910
transform 1 0 48116 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1626105910
transform 1 0 48208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_491
timestamp 1626105910
transform 1 0 46276 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_503
timestamp 1626105910
transform 1 0 47380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_479
timestamp 1626105910
transform 1 0 45172 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_467
timestamp 1626105910
transform 1 0 44068 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_455
timestamp 1626105910
transform 1 0 42964 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_493
timestamp 1626105910
transform 1 0 46460 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_505
timestamp 1626105910
transform 1 0 47564 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_481
timestamp 1626105910
transform 1 0 45356 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_469
timestamp 1626105910
transform 1 0 44252 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp 1626105910
transform 1 0 45540 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_455
timestamp 1626105910
transform 1 0 42964 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_463
timestamp 1626105910
transform 1 0 43700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__B1
timestamp 1626105910
transform 1 0 43516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A1
timestamp 1626105910
transform 1 0 44068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1626105910
transform -1 0 48852 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_514
timestamp 1626105910
transform 1 0 48392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1626105910
transform -1 0 48852 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1626105910
transform -1 0 48852 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1626105910
transform 1 0 48116 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1626105910
transform 1 0 48208 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_496
timestamp 1626105910
transform 1 0 46736 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_491
timestamp 1626105910
transform 1 0 46276 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_508
timestamp 1626105910
transform 1 0 47840 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_503
timestamp 1626105910
transform 1 0 47380 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_484
timestamp 1626105910
transform 1 0 45632 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_479
timestamp 1626105910
transform 1 0 45172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1626105910
transform 1 0 45540 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_475
timestamp 1626105910
transform 1 0 44804 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_463
timestamp 1626105910
transform 1 0 43700 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_459
timestamp 1626105910
transform 1 0 43332 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_467
timestamp 1626105910
transform 1 0 44068 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_455
timestamp 1626105910
transform 1 0 42964 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1626105910
transform 1 0 42964 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_456
timestamp 1626105910
transform 1 0 43056 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1626105910
transform -1 0 48852 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1626105910
transform -1 0 48852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1626105910
transform 1 0 48116 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1626105910
transform 1 0 48208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_496
timestamp 1626105910
transform 1 0 46736 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_496
timestamp 1626105910
transform 1 0 46736 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_508
timestamp 1626105910
transform 1 0 47840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_508
timestamp 1626105910
transform 1 0 47840 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _099_
timestamp 1626105910
transform 1 0 44436 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_2_484
timestamp 1626105910
transform 1 0 45632 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_484
timestamp 1626105910
transform 1 0 45632 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1626105910
transform 1 0 45540 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1626105910
transform -1 0 48852 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_438
timestamp 1626105910
transform 1 0 41400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__B1
timestamp 1626105910
transform 1 0 41584 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_426
timestamp 1626105910
transform 1 0 40296 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_414
timestamp 1626105910
transform 1 0 39192 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1626105910
transform -1 0 38732 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_452
timestamp 1626105910
transform 1 0 42688 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_404
timestamp 1626105910
transform 1 0 38272 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1626105910
transform 1 0 37628 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_442
timestamp 1626105910
transform 1 0 41768 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A3
timestamp 1626105910
transform -1 0 41952 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A2
timestamp 1626105910
transform 1 0 41584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_444
timestamp 1626105910
transform 1 0 41952 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_434
timestamp 1626105910
transform 1 0 41032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _086_
timestamp 1626105910
transform 1 0 37904 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_436
timestamp 1626105910
transform 1 0 41216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_438
timestamp 1626105910
transform 1 0 41400 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__C1
timestamp 1626105910
transform -1 0 41400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A1
timestamp 1626105910
transform -1 0 41216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_433
timestamp 1626105910
transform 1 0 40940 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_412
timestamp 1626105910
transform 1 0 39008 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_414
timestamp 1626105910
transform 1 0 39192 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_424
timestamp 1626105910
transform 1 0 40112 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1626105910
transform 1 0 40296 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_427
timestamp 1626105910
transform 1 0 40388 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_426
timestamp 1626105910
transform 1 0 40296 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_402
timestamp 1626105910
transform 1 0 38088 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_402
timestamp 1626105910
transform 1 0 38088 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1626105910
transform 1 0 37628 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1626105910
transform 1 0 37628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1626105910
transform 1 0 37628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_439
timestamp 1626105910
transform 1 0 41492 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_427
timestamp 1626105910
transform 1 0 40388 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_424
timestamp 1626105910
transform 1 0 40112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1626105910
transform 1 0 40296 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_416
timestamp 1626105910
transform 1 0 39376 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1626105910
transform 1 0 37628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_407
timestamp 1626105910
transform 1 0 38548 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A2
timestamp 1626105910
transform -1 0 38088 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_450
timestamp 1626105910
transform 1 0 42504 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_430
timestamp 1626105910
transform 1 0 40664 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_442
timestamp 1626105910
transform 1 0 41768 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__CLK
timestamp 1626105910
transform 1 0 42320 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_1  _060_
timestamp 1626105910
transform 1 0 39468 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_424
timestamp 1626105910
transform 1 0 40112 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_413
timestamp 1626105910
transform 1 0 39100 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A1
timestamp 1626105910
transform 1 0 38916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A3
timestamp 1626105910
transform 1 0 40480 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_410
timestamp 1626105910
transform 1 0 38824 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1626105910
transform 1 0 37628 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_452
timestamp 1626105910
transform 1 0 42688 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1626105910
transform 1 0 37628 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1626105910
transform -1 0 38088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_439
timestamp 1626105910
transform 1 0 41492 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A3
timestamp 1626105910
transform 1 0 37904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_402
timestamp 1626105910
transform 1 0 38088 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_400
timestamp 1626105910
transform 1 0 37904 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1626105910
transform 1 0 37628 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_408
timestamp 1626105910
transform 1 0 38640 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1626105910
transform 1 0 37628 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_402
timestamp 1626105910
transform 1 0 38088 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_COMP_INP
timestamp 1626105910
transform 1 0 38456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B2
timestamp 1626105910
transform 1 0 37904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_432
timestamp 1626105910
transform 1 0 40848 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1626105910
transform -1 0 38180 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_409
timestamp 1626105910
transform 1 0 38732 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1626105910
transform 1 0 37628 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1626105910
transform 1 0 38180 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_444
timestamp 1626105910
transform 1 0 41952 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_427
timestamp 1626105910
transform 1 0 40388 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_420
timestamp 1626105910
transform 1 0 39744 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1626105910
transform 1 0 40296 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_421
timestamp 1626105910
transform 1 0 39836 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_415
timestamp 1626105910
transform 1 0 39284 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__B1
timestamp 1626105910
transform -1 0 39836 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A2
timestamp 1626105910
transform -1 0 39284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_425
timestamp 1626105910
transform 1 0 40204 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_412
timestamp 1626105910
transform 1 0 39008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B1
timestamp 1626105910
transform -1 0 38088 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_439
timestamp 1626105910
transform 1 0 41492 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_427
timestamp 1626105910
transform 1 0 40388 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1626105910
transform 1 0 40296 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_421
timestamp 1626105910
transform 1 0 39836 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_425
timestamp 1626105910
transform 1 0 40204 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1626105910
transform 1 0 37904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_453
timestamp 1626105910
transform 1 0 42780 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_437
timestamp 1626105910
transform 1 0 41308 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp 1626105910
transform 1 0 42412 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_425
timestamp 1626105910
transform 1 0 40204 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_413
timestamp 1626105910
transform 1 0 39100 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A1
timestamp 1626105910
transform 1 0 38916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_400
timestamp 1626105910
transform 1 0 37904 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_439
timestamp 1626105910
transform 1 0 41492 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_427
timestamp 1626105910
transform 1 0 40388 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_414
timestamp 1626105910
transform 1 0 39192 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1626105910
transform 1 0 40296 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_402
timestamp 1626105910
transform 1 0 38088 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_442
timestamp 1626105910
transform 1 0 41768 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_400
timestamp 1626105910
transform 1 0 37904 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_450
timestamp 1626105910
transform 1 0 42504 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_452
timestamp 1626105910
transform 1 0 42688 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_450
timestamp 1626105910
transform 1 0 42504 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_440
timestamp 1626105910
transform 1 0 41584 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_428
timestamp 1626105910
transform 1 0 40480 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_416
timestamp 1626105910
transform 1 0 39376 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_410
timestamp 1626105910
transform 1 0 38824 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1626105910
transform 1 0 39192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_438
timestamp 1626105910
transform 1 0 41400 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_426
timestamp 1626105910
transform 1 0 40296 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_414
timestamp 1626105910
transform 1 0 39192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1626105910
transform 1 0 37628 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1626105910
transform 1 0 37628 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_400
timestamp 1626105910
transform 1 0 37904 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _093_
timestamp 1626105910
transform -1 0 38364 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_17_400
timestamp 1626105910
transform 1 0 37904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_439
timestamp 1626105910
transform 1 0 41492 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_427
timestamp 1626105910
transform 1 0 40388 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_412
timestamp 1626105910
transform 1 0 39008 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_424
timestamp 1626105910
transform 1 0 40112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1626105910
transform 1 0 40296 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_402
timestamp 1626105910
transform 1 0 38088 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1626105910
transform 1 0 37628 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1626105910
transform 1 0 37628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_438
timestamp 1626105910
transform 1 0 41400 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1626105910
transform 1 0 37628 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_405
timestamp 1626105910
transform 1 0 38364 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__B
timestamp 1626105910
transform -1 0 38916 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_439
timestamp 1626105910
transform 1 0 41492 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_427
timestamp 1626105910
transform 1 0 40388 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_412
timestamp 1626105910
transform 1 0 39008 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_424
timestamp 1626105910
transform 1 0 40112 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_436
timestamp 1626105910
transform 1 0 41216 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_448
timestamp 1626105910
transform 1 0 42320 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_424
timestamp 1626105910
transform 1 0 40112 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_412
timestamp 1626105910
transform 1 0 39008 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1626105910
transform 1 0 40296 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1626105910
transform -1 0 38088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_400
timestamp 1626105910
transform 1 0 37904 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_402
timestamp 1626105910
transform 1 0 38088 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_400
timestamp 1626105910
transform 1 0 37904 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1626105910
transform 1 0 37628 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1626105910
transform 1 0 37628 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1626105910
transform 1 0 37628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_COMP_INN
timestamp 1626105910
transform 1 0 37904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_439
timestamp 1626105910
transform 1 0 41492 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_427
timestamp 1626105910
transform 1 0 40388 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1626105910
transform 1 0 37628 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_439
timestamp 1626105910
transform 1 0 41492 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_450
timestamp 1626105910
transform 1 0 42504 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A1
timestamp 1626105910
transform 1 0 37904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_411
timestamp 1626105910
transform 1 0 38916 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_426
timestamp 1626105910
transform 1 0 40296 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_414
timestamp 1626105910
transform 1 0 39192 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_427
timestamp 1626105910
transform 1 0 40388 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_412
timestamp 1626105910
transform 1 0 39008 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_424
timestamp 1626105910
transform 1 0 40112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1626105910
transform 1 0 40296 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_438
timestamp 1626105910
transform 1 0 41400 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_426
timestamp 1626105910
transform 1 0 40296 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_414
timestamp 1626105910
transform 1 0 39192 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_402
timestamp 1626105910
transform 1 0 38088 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_423
timestamp 1626105910
transform 1 0 40020 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1626105910
transform 1 0 40296 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _059_
timestamp 1626105910
transform 1 0 38272 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_467
timestamp 1626105910
transform 1 0 44068 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_455
timestamp 1626105910
transform 1 0 42964 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_491
timestamp 1626105910
transform 1 0 46276 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1626105910
transform -1 0 48852 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_496
timestamp 1626105910
transform 1 0 46736 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_508
timestamp 1626105910
transform 1 0 47840 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_484
timestamp 1626105910
transform 1 0 45632 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1626105910
transform 1 0 45540 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_475
timestamp 1626105910
transform 1 0 44804 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_463
timestamp 1626105910
transform 1 0 43700 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_496
timestamp 1626105910
transform 1 0 46736 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1626105910
transform -1 0 48852 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1626105910
transform 1 0 48116 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_512
timestamp 1626105910
transform 1 0 48208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_510
timestamp 1626105910
transform 1 0 48024 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_498
timestamp 1626105910
transform 1 0 46920 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_486
timestamp 1626105910
transform 1 0 45816 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _106_
timestamp 1626105910
transform 1 0 44068 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_15_503
timestamp 1626105910
transform 1 0 47380 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_455
timestamp 1626105910
transform 1 0 42964 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_463
timestamp 1626105910
transform 1 0 43700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__D
timestamp 1626105910
transform -1 0 43700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1626105910
transform -1 0 48852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_496
timestamp 1626105910
transform 1 0 46736 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_508
timestamp 1626105910
transform 1 0 47840 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_484
timestamp 1626105910
transform 1 0 45632 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1626105910
transform 1 0 45540 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1626105910
transform 1 0 44988 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_465
timestamp 1626105910
transform 1 0 43884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_508
timestamp 1626105910
transform 1 0 47840 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__CLK
timestamp 1626105910
transform 1 0 43700 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_479
timestamp 1626105910
transform 1 0 45172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_484
timestamp 1626105910
transform 1 0 45632 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1626105910
transform -1 0 48852 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1626105910
transform 1 0 48116 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1626105910
transform 1 0 48208 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_491
timestamp 1626105910
transform 1 0 46276 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_503
timestamp 1626105910
transform 1 0 47380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_479
timestamp 1626105910
transform 1 0 45172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_467
timestamp 1626105910
transform 1 0 44068 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_455
timestamp 1626105910
transform 1 0 42964 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1626105910
transform 1 0 45540 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1626105910
transform -1 0 48852 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1626105910
transform 1 0 48208 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1626105910
transform -1 0 48208 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_496
timestamp 1626105910
transform 1 0 46736 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_505
timestamp 1626105910
transform 1 0 47564 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1626105910
transform -1 0 47564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_502
timestamp 1626105910
transform 1 0 47288 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_484
timestamp 1626105910
transform 1 0 45632 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1626105910
transform 1 0 45540 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_475
timestamp 1626105910
transform 1 0 44804 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_463
timestamp 1626105910
transform 1 0 43700 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_475
timestamp 1626105910
transform 1 0 44804 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1626105910
transform -1 0 48852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1626105910
transform 1 0 48116 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1626105910
transform 1 0 48208 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_491
timestamp 1626105910
transform 1 0 46276 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_503
timestamp 1626105910
transform 1 0 47380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_479
timestamp 1626105910
transform 1 0 45172 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_467
timestamp 1626105910
transform 1 0 44068 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_455
timestamp 1626105910
transform 1 0 42964 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_467
timestamp 1626105910
transform 1 0 44068 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_455
timestamp 1626105910
transform 1 0 42964 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_463
timestamp 1626105910
transform 1 0 43700 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_503
timestamp 1626105910
transform 1 0 47380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_479
timestamp 1626105910
transform 1 0 45172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1626105910
transform -1 0 48852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1626105910
transform 1 0 48116 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_512
timestamp 1626105910
transform 1 0 48208 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1626105910
transform -1 0 48852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1626105910
transform -1 0 48852 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_491
timestamp 1626105910
transform 1 0 46276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1626105910
transform 1 0 48116 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_512
timestamp 1626105910
transform 1 0 48208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1626105910
transform 1 0 42872 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_451
timestamp 1626105910
transform 1 0 42596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1626105910
transform 1 0 42872 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_451
timestamp 1626105910
transform 1 0 42596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1626105910
transform 1 0 37628 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_407
timestamp 1626105910
transform 1 0 38548 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1626105910
transform 1 0 42872 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_451
timestamp 1626105910
transform 1 0 42596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1626105910
transform 1 0 42872 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1626105910
transform -1 0 48852 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_496
timestamp 1626105910
transform 1 0 46736 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_508
timestamp 1626105910
transform 1 0 47840 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_484
timestamp 1626105910
transform 1 0 45632 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_471
timestamp 1626105910
transform 1 0 44436 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1626105910
transform 1 0 45540 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _110_
timestamp 1626105910
transform 1 0 42688 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_10_439
timestamp 1626105910
transform 1 0 41492 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_448
timestamp 1626105910
transform 1 0 42320 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__D
timestamp 1626105910
transform 1 0 42136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_445
timestamp 1626105910
transform 1 0 42044 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_427
timestamp 1626105910
transform 1 0 40388 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1626105910
transform 1 0 40296 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_419
timestamp 1626105910
transform 1 0 39652 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_413
timestamp 1626105910
transform 1 0 39100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__B1
timestamp 1626105910
transform -1 0 39652 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A2
timestamp 1626105910
transform 1 0 38916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_425
timestamp 1626105910
transform 1 0 40204 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1626105910
transform 1 0 42872 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_451
timestamp 1626105910
transform 1 0 42596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1626105910
transform 1 0 42872 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_451
timestamp 1626105910
transform 1 0 42596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1626105910
transform 1 0 42872 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_451
timestamp 1626105910
transform 1 0 42596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1626105910
transform 1 0 42872 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1626105910
transform 1 0 42872 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_2  _064_
timestamp 1626105910
transform -1 0 42964 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_451
timestamp 1626105910
transform 1 0 42596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_2  _066_
timestamp 1626105910
transform 1 0 37904 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_14_451
timestamp 1626105910
transform 1 0 42596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1626105910
transform 1 0 42872 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_270
timestamp 1626105910
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1626105910
transform -1 0 25944 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_265
timestamp 1626105910
transform 1 0 25484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_266
timestamp 1626105910
transform 1 0 25576 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_298
timestamp 1626105910
transform 1 0 28520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1626105910
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_306
timestamp 1626105910
transform 1 0 29256 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_294
timestamp 1626105910
transform 1 0 28152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_282
timestamp 1626105910
transform 1 0 27048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_286
timestamp 1626105910
transform 1 0 27416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1626105910
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_306
timestamp 1626105910
transform 1 0 29256 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_294
timestamp 1626105910
transform 1 0 28152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1626105910
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_277
timestamp 1626105910
transform 1 0 26588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1626105910
transform 1 0 26496 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1626105910
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1626105910
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1626105910
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_262
timestamp 1626105910
transform 1 0 25208 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1626105910
transform 1 0 25116 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_301
timestamp 1626105910
transform 1 0 28796 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_289
timestamp 1626105910
transform 1 0 27692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1626105910
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__B
timestamp 1626105910
transform -1 0 27692 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_286
timestamp 1626105910
transform 1 0 27416 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_277
timestamp 1626105910
transform 1 0 26588 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1626105910
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1626105910
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1626105910
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1626105910
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1626105910
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1626105910
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1626105910
transform 1 0 26312 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_277
timestamp 1626105910
transform 1 0 26588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_310
timestamp 1626105910
transform 1 0 29624 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_265
timestamp 1626105910
transform 1 0 25484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_298
timestamp 1626105910
transform 1 0 28520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1626105910
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1626105910
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_298
timestamp 1626105910
transform 1 0 28520 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1626105910
transform 1 0 30452 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__CLK
timestamp 1626105910
transform 1 0 28888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_304
timestamp 1626105910
transform 1 0 29072 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1626105910
transform 1 0 30544 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _114_
timestamp 1626105910
transform 1 0 26956 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_32_318
timestamp 1626105910
transform 1 0 30360 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_312
timestamp 1626105910
transform 1 0 29808 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_305
timestamp 1626105910
transform 1 0 29164 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1626105910
transform 1 0 29532 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _100_
timestamp 1626105910
transform -1 0 27324 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_32_293
timestamp 1626105910
transform 1 0 28060 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1626105910
transform 1 0 27784 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_274
timestamp 1626105910
transform 1 0 26312 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_285
timestamp 1626105910
transform 1 0 27324 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1626105910
transform 1 0 27876 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_289
timestamp 1626105910
transform 1 0 27692 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_277
timestamp 1626105910
transform 1 0 26588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__D
timestamp 1626105910
transform 1 0 26404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_312
timestamp 1626105910
transform 1 0 29808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_300
timestamp 1626105910
transform 1 0 28704 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_310
timestamp 1626105910
transform 1 0 29624 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1626105910
transform 1 0 28520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_312
timestamp 1626105910
transform 1 0 29808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1626105910
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_288
timestamp 1626105910
transform 1 0 27600 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_310
timestamp 1626105910
transform 1 0 29624 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1626105910
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1626105910
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_363
timestamp 1626105910
transform 1 0 34500 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1626105910
transform 1 0 33396 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_339
timestamp 1626105910
transform 1 0 32292 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_327
timestamp 1626105910
transform 1 0 31188 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1626105910
transform 1 0 31188 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1626105910
transform 1 0 31188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1626105910
transform 1 0 34868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1626105910
transform 1 0 33764 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1626105910
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1626105910
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_341
timestamp 1626105910
transform 1 0 32476 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_325
timestamp 1626105910
transform 1 0 31004 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1626105910
transform 1 0 32108 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _050_
timestamp 1626105910
transform 1 0 35696 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1626105910
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_361
timestamp 1626105910
transform 1 0 34316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1626105910
transform 1 0 35788 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_373
timestamp 1626105910
transform 1 0 35420 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_349
timestamp 1626105910
transform 1 0 33212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1626105910
transform 1 0 33120 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_343
timestamp 1626105910
transform 1 0 32660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__B
timestamp 1626105910
transform 1 0 32476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_347
timestamp 1626105910
transform 1 0 33028 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1626105910
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_337
timestamp 1626105910
transform 1 0 32108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_331
timestamp 1626105910
transform 1 0 31556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1626105910
transform 1 0 31924 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_376
timestamp 1626105910
transform 1 0 35696 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_367
timestamp 1626105910
transform 1 0 34868 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__A
timestamp 1626105910
transform 1 0 35512 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_373
timestamp 1626105910
transform 1 0 35420 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1626105910
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1626105910
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1626105910
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_372
timestamp 1626105910
transform 1 0 35328 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_334
timestamp 1626105910
transform 1 0 31832 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_372
timestamp 1626105910
transform 1 0 35328 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_367
timestamp 1626105910
transform 1 0 34868 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_355
timestamp 1626105910
transform 1 0 33764 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_343
timestamp 1626105910
transform 1 0 32660 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1626105910
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_363
timestamp 1626105910
transform 1 0 34500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_372
timestamp 1626105910
transform 1 0 35328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_334
timestamp 1626105910
transform 1 0 31832 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1626105910
transform 1 0 34868 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1626105910
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_363
timestamp 1626105910
transform 1 0 34500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1626105910
transform 1 0 33396 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1626105910
transform 1 0 32292 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_355
timestamp 1626105910
transform 1 0 33764 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_343
timestamp 1626105910
transform 1 0 32660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1626105910
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_327
timestamp 1626105910
transform 1 0 31188 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1626105910
transform 1 0 33396 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_334
timestamp 1626105910
transform 1 0 31832 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1626105910
transform 1 0 32292 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_372
timestamp 1626105910
transform 1 0 35328 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1626105910
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_363
timestamp 1626105910
transform 1 0 34500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1626105910
transform 1 0 33396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1626105910
transform 1 0 32292 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_315
timestamp 1626105910
transform 1 0 30084 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1626105910
transform 1 0 30084 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_313
timestamp 1626105910
transform 1 0 29900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _056_
timestamp 1626105910
transform 1 0 30912 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_39_322
timestamp 1626105910
transform 1 0 30728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_322
timestamp 1626105910
transform 1 0 30728 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1626105910
transform 1 0 30728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_315
timestamp 1626105910
transform 1 0 30084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1626105910
transform 1 0 30084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_467
timestamp 1626105910
transform 1 0 44068 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_455
timestamp 1626105910
transform 1 0 42964 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1626105910
transform 1 0 48208 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_496
timestamp 1626105910
transform 1 0 46736 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_491
timestamp 1626105910
transform 1 0 46276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_508
timestamp 1626105910
transform 1 0 47840 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1626105910
transform -1 0 48852 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1626105910
transform 1 0 48116 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_512
timestamp 1626105910
transform 1 0 48208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_491
timestamp 1626105910
transform 1 0 46276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1626105910
transform -1 0 48852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_496
timestamp 1626105910
transform 1 0 46736 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_508
timestamp 1626105910
transform 1 0 47840 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_484
timestamp 1626105910
transform 1 0 45632 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1626105910
transform 1 0 45540 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_475
timestamp 1626105910
transform 1 0 44804 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_463
timestamp 1626105910
transform 1 0 43700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_503
timestamp 1626105910
transform 1 0 47380 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_479
timestamp 1626105910
transform 1 0 45172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_467
timestamp 1626105910
transform 1 0 44068 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_455
timestamp 1626105910
transform 1 0 42964 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_503
timestamp 1626105910
transform 1 0 47380 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_484
timestamp 1626105910
transform 1 0 45632 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1626105910
transform -1 0 48852 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1626105910
transform 1 0 48116 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_512
timestamp 1626105910
transform 1 0 48208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_491
timestamp 1626105910
transform 1 0 46276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_503
timestamp 1626105910
transform 1 0 47380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_479
timestamp 1626105910
transform 1 0 45172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_467
timestamp 1626105910
transform 1 0 44068 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_455
timestamp 1626105910
transform 1 0 42964 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_479
timestamp 1626105910
transform 1 0 45172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1626105910
transform 1 0 45540 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_475
timestamp 1626105910
transform 1 0 44804 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_463
timestamp 1626105910
transform 1 0 43700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_455
timestamp 1626105910
transform 1 0 42964 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_467
timestamp 1626105910
transform 1 0 44068 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1626105910
transform -1 0 48852 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1626105910
transform 1 0 48116 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_512
timestamp 1626105910
transform 1 0 48208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_503
timestamp 1626105910
transform 1 0 47380 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_491
timestamp 1626105910
transform 1 0 46276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_479
timestamp 1626105910
transform 1 0 45172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_467
timestamp 1626105910
transform 1 0 44068 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_455
timestamp 1626105910
transform 1 0 42964 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1626105910
transform -1 0 48852 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1626105910
transform -1 0 48852 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_496
timestamp 1626105910
transform 1 0 46736 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_508
timestamp 1626105910
transform 1 0 47840 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_484
timestamp 1626105910
transform 1 0 45632 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1626105910
transform -1 0 48852 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_508
timestamp 1626105910
transform 1 0 47840 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_496
timestamp 1626105910
transform 1 0 46736 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_484
timestamp 1626105910
transform 1 0 45632 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1626105910
transform 1 0 45540 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_475
timestamp 1626105910
transform 1 0 44804 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_463
timestamp 1626105910
transform 1 0 43700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1626105910
transform 1 0 45540 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_482
timestamp 1626105910
transform 1 0 45448 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_474
timestamp 1626105910
transform 1 0 44712 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_462
timestamp 1626105910
transform 1 0 43608 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1626105910
transform -1 0 48852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1626105910
transform 1 0 48116 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1626105910
transform -1 0 48852 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1626105910
transform 1 0 48116 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_512
timestamp 1626105910
transform 1 0 48208 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_503
timestamp 1626105910
transform 1 0 47380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_491
timestamp 1626105910
transform 1 0 46276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_479
timestamp 1626105910
transform 1 0 45172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_424
timestamp 1626105910
transform 1 0 40112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1626105910
transform 1 0 40296 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_427
timestamp 1626105910
transform 1 0 40388 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_451
timestamp 1626105910
transform 1 0 42596 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_412
timestamp 1626105910
transform 1 0 39008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_431
timestamp 1626105910
transform 1 0 40756 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_443
timestamp 1626105910
transform 1 0 41860 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_412
timestamp 1626105910
transform 1 0 39008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_424
timestamp 1626105910
transform 1 0 40112 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__D
timestamp 1626105910
transform -1 0 40756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_428
timestamp 1626105910
transform 1 0 40480 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_424
timestamp 1626105910
transform 1 0 40112 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1626105910
transform 1 0 40296 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_400
timestamp 1626105910
transform 1 0 37904 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1626105910
transform 1 0 37628 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_400
timestamp 1626105910
transform 1 0 37904 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1626105910
transform 1 0 37628 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_400
timestamp 1626105910
transform 1 0 37904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1626105910
transform 1 0 37628 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_400
timestamp 1626105910
transform 1 0 37904 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1626105910
transform 1 0 37628 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_400
timestamp 1626105910
transform 1 0 37904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_400
timestamp 1626105910
transform 1 0 37904 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_400
timestamp 1626105910
transform 1 0 37904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1626105910
transform 1 0 37628 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1626105910
transform 1 0 37628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1626105910
transform 1 0 37628 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_400
timestamp 1626105910
transform 1 0 37904 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_400
timestamp 1626105910
transform 1 0 37904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1626105910
transform 1 0 37628 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1626105910
transform 1 0 37628 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_439
timestamp 1626105910
transform 1 0 41492 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_448
timestamp 1626105910
transform 1 0 42320 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_436
timestamp 1626105910
transform 1 0 41216 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_424
timestamp 1626105910
transform 1 0 40112 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_412
timestamp 1626105910
transform 1 0 39008 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_436
timestamp 1626105910
transform 1 0 41216 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_439
timestamp 1626105910
transform 1 0 41492 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_427
timestamp 1626105910
transform 1 0 40388 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_412
timestamp 1626105910
transform 1 0 39008 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_424
timestamp 1626105910
transform 1 0 40112 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1626105910
transform 1 0 40296 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_452
timestamp 1626105910
transform 1 0 42688 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_448
timestamp 1626105910
transform 1 0 42320 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_444
timestamp 1626105910
transform 1 0 41952 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _112_
timestamp 1626105910
transform -1 0 41952 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_27_423
timestamp 1626105910
transform 1 0 40020 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__CLK
timestamp 1626105910
transform 1 0 39836 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_420
timestamp 1626105910
transform 1 0 39744 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_412
timestamp 1626105910
transform 1 0 39008 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_427
timestamp 1626105910
transform 1 0 40388 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_439
timestamp 1626105910
transform 1 0 41492 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_427
timestamp 1626105910
transform 1 0 40388 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_412
timestamp 1626105910
transform 1 0 39008 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_424
timestamp 1626105910
transform 1 0 40112 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1626105910
transform 1 0 40296 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_412
timestamp 1626105910
transform 1 0 39008 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_453
timestamp 1626105910
transform 1 0 42780 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_441
timestamp 1626105910
transform 1 0 41676 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1626105910
transform 1 0 40572 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_412
timestamp 1626105910
transform 1 0 39008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_424
timestamp 1626105910
transform 1 0 40112 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__CLK
timestamp 1626105910
transform 1 0 40388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_424
timestamp 1626105910
transform 1 0 40112 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _107_
timestamp 1626105910
transform -1 0 42504 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_24_412
timestamp 1626105910
transform 1 0 39008 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_400
timestamp 1626105910
transform 1 0 37904 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1626105910
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_391
timestamp 1626105910
transform 1 0 37076 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_405
timestamp 1626105910
transform 1 0 38364 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_407
timestamp 1626105910
transform 1 0 38548 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1626105910
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_390
timestamp 1626105910
transform 1 0 36984 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1626105910
transform 1 0 38088 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_393
timestamp 1626105910
transform 1 0 37260 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_396
timestamp 1626105910
transform 1 0 37536 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_408
timestamp 1626105910
transform 1 0 38640 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_441
timestamp 1626105910
transform 1 0 41676 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_429
timestamp 1626105910
transform 1 0 40572 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_400
timestamp 1626105910
transform 1 0 37904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_400
timestamp 1626105910
transform 1 0 37904 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_436
timestamp 1626105910
transform 1 0 41216 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1626105910
transform 1 0 40480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_424
timestamp 1626105910
transform 1 0 40112 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_412
timestamp 1626105910
transform 1 0 39008 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_420
timestamp 1626105910
transform 1 0 39744 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_396
timestamp 1626105910
transform 1 0 37536 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_408
timestamp 1626105910
transform 1 0 38640 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_441
timestamp 1626105910
transform 1 0 41676 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_441
timestamp 1626105910
transform 1 0 41676 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_429
timestamp 1626105910
transform 1 0 40572 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1626105910
transform 1 0 40480 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_425
timestamp 1626105910
transform 1 0 40204 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_417
timestamp 1626105910
transform 1 0 39468 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_429
timestamp 1626105910
transform 1 0 40572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1626105910
transform 1 0 40480 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_420
timestamp 1626105910
transform 1 0 39744 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_396
timestamp 1626105910
transform 1 0 37536 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1626105910
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_441
timestamp 1626105910
transform 1 0 41676 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_429
timestamp 1626105910
transform 1 0 40572 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1626105910
transform 1 0 40480 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_420
timestamp 1626105910
transform 1 0 39744 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1626105910
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_436
timestamp 1626105910
transform 1 0 41216 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_424
timestamp 1626105910
transform 1 0 40112 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_412
timestamp 1626105910
transform 1 0 39008 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_408
timestamp 1626105910
transform 1 0 38640 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_436
timestamp 1626105910
transform 1 0 41216 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1626105910
transform 1 0 41124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_431
timestamp 1626105910
transform 1 0 40756 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_419
timestamp 1626105910
transform 1 0 39652 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_396
timestamp 1626105910
transform 1 0 37536 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_391
timestamp 1626105910
transform 1 0 37076 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_436
timestamp 1626105910
transform 1 0 41216 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_424
timestamp 1626105910
transform 1 0 40112 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_436
timestamp 1626105910
transform 1 0 41216 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_424
timestamp 1626105910
transform 1 0 40112 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_412
timestamp 1626105910
transform 1 0 39008 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_412
timestamp 1626105910
transform 1 0 39008 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_400
timestamp 1626105910
transform 1 0 37904 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1626105910
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_391
timestamp 1626105910
transform 1 0 37076 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1626105910
transform 1 0 43056 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_460
timestamp 1626105910
transform 1 0 43424 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1626105910
transform -1 0 48852 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_514
timestamp 1626105910
transform 1 0 48392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1626105910
transform -1 0 48852 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_510
timestamp 1626105910
transform 1 0 48024 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_498
timestamp 1626105910
transform 1 0 46920 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_486
timestamp 1626105910
transform 1 0 45816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1626105910
transform 1 0 45724 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_465
timestamp 1626105910
transform 1 0 43884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_477
timestamp 1626105910
transform 1 0 44988 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_506
timestamp 1626105910
transform 1 0 47656 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1626105910
transform -1 0 48852 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_514
timestamp 1626105910
transform 1 0 48392 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1626105910
transform 1 0 48300 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1626105910
transform 1 0 47564 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_493
timestamp 1626105910
transform 1 0 46460 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_481
timestamp 1626105910
transform 1 0 45356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_469
timestamp 1626105910
transform 1 0 44252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_457
timestamp 1626105910
transform 1 0 43148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1626105910
transform 1 0 43056 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_494
timestamp 1626105910
transform 1 0 46552 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1626105910
transform -1 0 48852 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1626105910
transform -1 0 48852 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_514
timestamp 1626105910
transform 1 0 48392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1626105910
transform 1 0 48300 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_510
timestamp 1626105910
transform 1 0 48024 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1626105910
transform 1 0 47564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_498
timestamp 1626105910
transform 1 0 46920 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_486
timestamp 1626105910
transform 1 0 45816 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_493
timestamp 1626105910
transform 1 0 46460 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1626105910
transform 1 0 45724 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_465
timestamp 1626105910
transform 1 0 43884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_481
timestamp 1626105910
transform 1 0 45356 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_469
timestamp 1626105910
transform 1 0 44252 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1626105910
transform 1 0 44988 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1626105910
transform 1 0 46460 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_457
timestamp 1626105910
transform 1 0 43148 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1626105910
transform 1 0 43056 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_489
timestamp 1626105910
transform 1 0 46092 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1626105910
transform -1 0 48852 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_510
timestamp 1626105910
transform 1 0 48024 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_498
timestamp 1626105910
transform 1 0 46920 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_486
timestamp 1626105910
transform 1 0 45816 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1626105910
transform 1 0 45724 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_465
timestamp 1626105910
transform 1 0 43884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_477
timestamp 1626105910
transform 1 0 44988 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1626105910
transform 1 0 44988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1626105910
transform -1 0 48852 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_514
timestamp 1626105910
transform 1 0 48392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1626105910
transform 1 0 48300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1626105910
transform 1 0 47564 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_493
timestamp 1626105910
transform 1 0 46460 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_481
timestamp 1626105910
transform 1 0 45356 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_469
timestamp 1626105910
transform 1 0 44252 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_457
timestamp 1626105910
transform 1 0 43148 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1626105910
transform 1 0 43056 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_465
timestamp 1626105910
transform 1 0 43884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1626105910
transform -1 0 48852 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_510
timestamp 1626105910
transform 1 0 48024 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_498
timestamp 1626105910
transform 1 0 46920 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_486
timestamp 1626105910
transform 1 0 45816 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1626105910
transform 1 0 45724 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_465
timestamp 1626105910
transform 1 0 43884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_477
timestamp 1626105910
transform 1 0 44988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1626105910
transform 1 0 43792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1626105910
transform -1 0 48852 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_514
timestamp 1626105910
transform 1 0 48392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1626105910
transform 1 0 48300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1626105910
transform 1 0 47564 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_493
timestamp 1626105910
transform 1 0 46460 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_481
timestamp 1626105910
transform 1 0 45356 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_469
timestamp 1626105910
transform 1 0 44252 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_457
timestamp 1626105910
transform 1 0 43148 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_400
timestamp 1626105910
transform 1 0 37904 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_400
timestamp 1626105910
transform 1 0 37904 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1626105910
transform 1 0 37628 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1626105910
transform 1 0 37628 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_453
timestamp 1626105910
transform 1 0 42780 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_448
timestamp 1626105910
transform 1 0 42320 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_453
timestamp 1626105910
transform 1 0 42780 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_448
timestamp 1626105910
transform 1 0 42320 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_453
timestamp 1626105910
transform 1 0 42780 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_448
timestamp 1626105910
transform 1 0 42320 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_453
timestamp 1626105910
transform 1 0 42780 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_448
timestamp 1626105910
transform 1 0 42320 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_448
timestamp 1626105910
transform 1 0 42320 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1626105910
transform -1 0 48852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1626105910
transform -1 0 48852 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1626105910
transform 1 0 48116 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1626105910
transform 1 0 48208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_503
timestamp 1626105910
transform 1 0 47380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_508
timestamp 1626105910
transform 1 0 47840 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_491
timestamp 1626105910
transform 1 0 46276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_496
timestamp 1626105910
transform 1 0 46736 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_484
timestamp 1626105910
transform 1 0 45632 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1626105910
transform 1 0 45540 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_479
timestamp 1626105910
transform 1 0 45172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_467
timestamp 1626105910
transform 1 0 44068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_475
timestamp 1626105910
transform 1 0 44804 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_455
timestamp 1626105910
transform 1 0 42964 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_463
timestamp 1626105910
transform 1 0 43700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_451
timestamp 1626105910
transform 1 0 42596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1626105910
transform 1 0 42872 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_448
timestamp 1626105910
transform 1 0 42320 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_436
timestamp 1626105910
transform 1 0 41216 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_439
timestamp 1626105910
transform 1 0 41492 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_424
timestamp 1626105910
transform 1 0 40112 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_412
timestamp 1626105910
transform 1 0 39008 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_427
timestamp 1626105910
transform 1 0 40388 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_412
timestamp 1626105910
transform 1 0 39008 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_424
timestamp 1626105910
transform 1 0 40112 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1626105910
transform 1 0 40296 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1626105910
transform 1 0 42872 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_451
timestamp 1626105910
transform 1 0 42596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1626105910
transform 1 0 42872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_451
timestamp 1626105910
transform 1 0 42596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1626105910
transform 1 0 42872 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_450
timestamp 1626105910
transform 1 0 42504 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1626105910
transform 1 0 42872 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_451
timestamp 1626105910
transform 1 0 42596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1626105910
transform 1 0 42872 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1626105910
transform 1 0 35972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_378
timestamp 1626105910
transform 1 0 35880 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_400
timestamp 1626105910
transform 1 0 37904 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1626105910
transform 1 0 37628 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1626105910
transform -1 0 48852 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_496
timestamp 1626105910
transform 1 0 46736 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_508
timestamp 1626105910
transform 1 0 47840 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_484
timestamp 1626105910
transform 1 0 45632 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1626105910
transform 1 0 45540 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_475
timestamp 1626105910
transform 1 0 44804 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_463
timestamp 1626105910
transform 1 0 43700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_451
timestamp 1626105910
transform 1 0 42596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_439
timestamp 1626105910
transform 1 0 41492 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_427
timestamp 1626105910
transform 1 0 40388 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_412
timestamp 1626105910
transform 1 0 39008 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_424
timestamp 1626105910
transform 1 0 40112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1626105910
transform 1 0 40296 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_381
timestamp 1626105910
transform 1 0 36156 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_388
timestamp 1626105910
transform 1 0 36800 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_384
timestamp 1626105910
transform 1 0 36432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_379
timestamp 1626105910
transform 1 0 35972 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_384
timestamp 1626105910
transform 1 0 36432 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_379
timestamp 1626105910
transform 1 0 35972 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_384
timestamp 1626105910
transform 1 0 36432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1626105910
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_188
timestamp 1626105910
transform 1 0 18400 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1626105910
transform -1 0 18952 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1626105910
transform -1 0 18952 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_190
timestamp 1626105910
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_184
timestamp 1626105910
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_180
timestamp 1626105910
transform 1 0 17664 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1626105910
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1626105910
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1626105910
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1626105910
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1626105910
transform 1 0 15456 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1626105910
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1626105910
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1626105910
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1626105910
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1626105910
transform -1 0 18952 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1626105910
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1626105910
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1626105910
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1626105910
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_158
timestamp 1626105910
transform 1 0 15640 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1626105910
transform 1 0 14536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1626105910
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1626105910
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1626105910
transform -1 0 18952 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_187
timestamp 1626105910
transform 1 0 18308 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1626105910
transform 1 0 17756 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1626105910
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_COMP_clk
timestamp 1626105910
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A2
timestamp 1626105910
transform 1 0 18124 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_178
timestamp 1626105910
transform 1 0 17480 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1626105910
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_172
timestamp 1626105910
transform 1 0 16928 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1626105910
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1626105910
transform 1 0 14996 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_172
timestamp 1626105910
transform 1 0 16928 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1626105910
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1626105910
transform -1 0 18952 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1626105910
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1626105910
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A1
timestamp 1626105910
transform -1 0 18308 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_184
timestamp 1626105910
transform 1 0 18032 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1626105910
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1626105910
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1626105910
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1626105910
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1626105910
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1626105910
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1626105910
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1626105910
transform -1 0 18952 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1626105910
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_190
timestamp 1626105910
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1626105910
transform -1 0 18952 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_184
timestamp 1626105910
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _082_
timestamp 1626105910
transform -1 0 18308 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1626105910
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1626105910
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_187
timestamp 1626105910
transform 1 0 18308 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_163
timestamp 1626105910
transform 1 0 16100 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_177
timestamp 1626105910
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_172
timestamp 1626105910
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1626105910
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1626105910
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1626105910
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1626105910
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1626105910
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1626105910
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1626105910
transform 1 0 14996 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1626105910
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1626105910
transform -1 0 18952 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1626105910
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_187
timestamp 1626105910
transform 1 0 18308 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_180
timestamp 1626105910
transform 1 0 17664 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__C1
timestamp 1626105910
transform -1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_184
timestamp 1626105910
transform 1 0 18032 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1626105910
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1626105910
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1626105910
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1626105910
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1626105910
transform -1 0 18952 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1626105910
transform -1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _070_
timestamp 1626105910
transform -1 0 18308 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1626105910
transform 1 0 18308 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1626105910
transform 1 0 18308 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__B1
timestamp 1626105910
transform 1 0 18124 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1626105910
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1626105910
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1626105910
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1626105910
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1626105910
transform 1 0 17204 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_168
timestamp 1626105910
transform 1 0 16560 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1626105910
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A3
timestamp 1626105910
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_134
timestamp 1626105910
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1626105910
transform -1 0 18952 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1626105910
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_190
timestamp 1626105910
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1626105910
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1626105910
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1626105910
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1626105910
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1626105910
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1626105910
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1626105910
transform -1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_188
timestamp 1626105910
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_180
timestamp 1626105910
transform 1 0 17664 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1626105910
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1626105910
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1626105910
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1626105910
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1626105910
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1626105910
transform -1 0 18952 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1626105910
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_190
timestamp 1626105910
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1626105910
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1626105910
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1626105910
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1626105910
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1626105910
transform -1 0 18952 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_188
timestamp 1626105910
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_180
timestamp 1626105910
transform 1 0 17664 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1626105910
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1626105910
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1626105910
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1626105910
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1626105910
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1626105910
transform -1 0 18952 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1626105910
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_190
timestamp 1626105910
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1626105910
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1626105910
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1626105910
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1626105910
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1626105910
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1626105910
transform -1 0 18952 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_188
timestamp 1626105910
transform 1 0 18400 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_180
timestamp 1626105910
transform 1 0 17664 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1626105910
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1626105910
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1626105910
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1626105910
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1626105910
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_188
timestamp 1626105910
transform 1 0 18400 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1626105910
transform -1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1626105910
transform -1 0 18952 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_190
timestamp 1626105910
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1626105910
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_180
timestamp 1626105910
transform 1 0 17664 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1626105910
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1626105910
transform 1 0 16560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1626105910
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1626105910
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1626105910
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1626105910
transform 1 0 15456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1626105910
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1626105910
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1626105910
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1626105910
transform -1 0 18952 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_187
timestamp 1626105910
transform 1 0 18308 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 1626105910
transform 1 0 18124 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1626105910
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1626105910
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1626105910
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1626105910
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1626105910
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1626105910
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_136
timestamp 1626105910
transform 1 0 13616 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1626105910
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1626105910
transform -1 0 18952 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _092_
timestamp 1626105910
transform -1 0 18308 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1626105910
transform 1 0 18308 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1626105910
transform 1 0 17480 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1626105910
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_168
timestamp 1626105910
transform 1 0 16560 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1626105910
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1626105910
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1626105910
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1626105910
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1626105910
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1626105910
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_95
timestamp 1626105910
transform 1 0 9844 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1626105910
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_107
timestamp 1626105910
transform 1 0 10948 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1626105910
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1626105910
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1626105910
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_106
timestamp 1626105910
transform 1 0 10856 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1626105910
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1626105910
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1626105910
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1626105910
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1626105910
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1626105910
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1626105910
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1626105910
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1626105910
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_83
timestamp 1626105910
transform 1 0 8740 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1626105910
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1626105910
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1626105910
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1626105910
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1626105910
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_71
timestamp 1626105910
transform 1 0 7636 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1626105910
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1626105910
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1626105910
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1626105910
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1626105910
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1626105910
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1626105910
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1626105910
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1626105910
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1626105910
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1626105910
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__049__A
timestamp 1626105910
transform -1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104
timestamp 1626105910
transform 1 0 10672 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107
timestamp 1626105910
transform 1 0 10948 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1626105910
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1626105910
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1626105910
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1626105910
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1626105910
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1626105910
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1626105910
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1626105910
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1626105910
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1626105910
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_65
timestamp 1626105910
transform 1 0 7084 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1626105910
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1626105910
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1626105910
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1626105910
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1626105910
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1626105910
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1626105910
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1626105910
transform 1 0 11500 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1626105910
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1626105910
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1626105910
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1626105910
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1626105910
transform 1 0 11500 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _049_
timestamp 1626105910
transform -1 0 10764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1626105910
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_105
timestamp 1626105910
transform 1 0 10764 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_94
timestamp 1626105910
transform 1 0 9752 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1626105910
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1626105910
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1626105910
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1626105910
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1626105910
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1626105910
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1626105910
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1626105910
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1626105910
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1626105910
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1626105910
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1626105910
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1626105910
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1626105910
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_58
timestamp 1626105910
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1626105910
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1626105910
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1626105910
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1626105910
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1626105910
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1626105910
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1626105910
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_12
timestamp 1626105910
transform 1 0 2208 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1626105910
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1626105910
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1626105910
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1626105910
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1626105910
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1626105910
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1626105910
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1626105910
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1626105910
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1626105910
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1626105910
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1626105910
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1626105910
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1626105910
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1626105910
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1626105910
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1626105910
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1626105910
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1626105910
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6
timestamp 1626105910
transform 1 0 1656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1626105910
transform -1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1626105910
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1626105910
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1626105910
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1626105910
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1626105910
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51
timestamp 1626105910
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1626105910
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1626105910
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1626105910
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1626105910
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1626105910
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1626105910
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1626105910
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1626105910
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1626105910
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1626105910
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1626105910
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1626105910
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1626105910
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1626105910
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1626105910
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1626105910
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1626105910
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1626105910
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1626105910
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1626105910
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1626105910
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1626105910
transform 1 0 5428 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_35
timestamp 1626105910
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_23
timestamp 1626105910
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output14
timestamp 1626105910
transform -1 0 2116 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_11
timestamp 1626105910
transform 1 0 2116 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1626105910
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1626105910
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1626105910
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1626105910
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1626105910
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1626105910
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1626105910
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1626105910
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1626105910
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1626105910
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1626105910
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1626105910
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1626105910
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1626105910
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1626105910
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1626105910
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1626105910
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1626105910
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1626105910
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1626105910
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1626105910
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1626105910
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1626105910
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1626105910
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1626105910
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1626105910
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1626105910
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1626105910
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1626105910
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1626105910
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1626105910
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1626105910
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1626105910
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1626105910
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1626105910
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1626105910
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1626105910
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1626105910
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1626105910
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1626105910
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1626105910
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1626105910
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1626105910
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1626105910
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1626105910
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1626105910
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1626105910
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1626105910
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1626105910
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1626105910
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1626105910
transform -1 0 2116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_17
timestamp 1626105910
transform 1 0 2668 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1626105910
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1626105910
transform 1 0 2116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1626105910
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output6_A
timestamp 1626105910
transform -1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1626105910
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1626105910
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1626105910
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1626105910
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1626105910
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1626105910
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1626105910
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1626105910
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1626105910
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1626105910
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1626105910
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1626105910
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1626105910
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1626105910
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1626105910
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1626105910
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1626105910
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1626105910
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1626105910
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1626105910
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1626105910
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1626105910
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1626105910
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1626105910
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1626105910
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1626105910
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1626105910
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1626105910
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1626105910
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1626105910
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1626105910
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1626105910
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_106
timestamp 1626105910
transform 1 0 10856 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_112
timestamp 1626105910
transform 1 0 11408 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A2
timestamp 1626105910
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_107
timestamp 1626105910
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_99
timestamp 1626105910
transform 1 0 10212 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1626105910
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1626105910
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1626105910
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1626105910
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1626105910
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1626105910
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1626105910
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1626105910
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B1
timestamp 1626105910
transform 1 0 12236 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A3
timestamp 1626105910
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_2  _072_
timestamp 1626105910
transform -1 0 10856 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1626105910
transform 1 0 9752 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_98
timestamp 1626105910
transform 1 0 10120 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1626105910
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1626105910
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1626105910
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1626105910
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1626105910
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_110
timestamp 1626105910
transform 1 0 11224 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A1
timestamp 1626105910
transform -1 0 11224 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_107
timestamp 1626105910
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_99
timestamp 1626105910
transform 1 0 10212 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1626105910
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1626105910
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1626105910
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1626105910
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1626105910
transform 1 0 11316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1626105910
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1626105910
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1626105910
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1626105910
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1626105910
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1626105910
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1626105910
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1626105910
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1626105910
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1626105910
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1626105910
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1626105910
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1626105910
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1626105910
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1626105910
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1626105910
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1626105910
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1626105910
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1626105910
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1626105910
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1626105910
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1626105910
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1626105910
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1626105910
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1626105910
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1626105910
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1626105910
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1626105910
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1626105910
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1626105910
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1626105910
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1626105910
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1626105910
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1626105910
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1626105910
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1626105910
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1626105910
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1626105910
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1626105910
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1626105910
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1626105910
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1626105910
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1626105910
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1626105910
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1626105910
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1626105910
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1626105910
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1626105910
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1626105910
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1626105910
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1626105910
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1626105910
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1626105910
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1626105910
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1626105910
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1626105910
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1626105910
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1626105910
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1626105910
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1626105910
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1626105910
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1626105910
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1626105910
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1626105910
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1626105910
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1626105910
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1626105910
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1626105910
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1626105910
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1626105910
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1626105910
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1626105910
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1626105910
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1626105910
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1626105910
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1626105910
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1626105910
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1626105910
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1626105910
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1626105910
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1626105910
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1626105910
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1626105910
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1626105910
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1626105910
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_119
timestamp 1626105910
transform 1 0 12052 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1626105910
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_111
timestamp 1626105910
transform 1 0 11316 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1626105910
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1626105910
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1626105910
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1626105910
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1626105910
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1626105910
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1626105910
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1626105910
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1626105910
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1626105910
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1626105910
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1626105910
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1626105910
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1626105910
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1626105910
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1626105910
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1626105910
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1626105910
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1626105910
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1626105910
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1626105910
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1626105910
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1626105910
transform -1 0 2116 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_17
timestamp 1626105910
transform 1 0 2668 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1626105910
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1626105910
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1626105910
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1626105910
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1626105910
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1626105910
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1626105910
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1626105910
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1626105910
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1626105910
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1626105910
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1626105910
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1626105910
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1626105910
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1626105910
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1626105910
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1626105910
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_51
timestamp 1626105910
transform 1 0 5796 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1626105910
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1626105910
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1626105910
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1626105910
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1626105910
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1626105910
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1626105910
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1626105910
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1626105910
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output7_A
timestamp 1626105910
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1626105910
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1626105910
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1626105910
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1626105910
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1626105910
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1626105910
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1626105910
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1626105910
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1626105910
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1626105910
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1626105910
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1626105910
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1626105910
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1626105910
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1626105910
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1626105910
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1626105910
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1626105910
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1626105910
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_11
timestamp 1626105910
transform 1 0 2116 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1626105910
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1626105910
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1626105910
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1626105910
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1626105910
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1626105910
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1626105910
transform 1 0 6440 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1626105910
transform 1 0 6072 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1626105910
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1626105910
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1626105910
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1626105910
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1626105910
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1626105910
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1626105910
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1626105910
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1626105910
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1626105910
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1626105910
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1626105910
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1626105910
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1626105910
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1626105910
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1626105910
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1626105910
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1626105910
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1626105910
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1626105910
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1626105910
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1626105910
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_51
timestamp 1626105910
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1626105910
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_51
timestamp 1626105910
transform 1 0 5796 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1626105910
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1626105910
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1626105910
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1626105910
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1626105910
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1626105910
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1626105910
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1626105910
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1626105910
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1626105910
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1626105910
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1626105910
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1626105910
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1626105910
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1626105910
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1626105910
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1626105910
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1626105910
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1626105910
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1626105910
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_41
timestamp 1626105910
transform 1 0 4876 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1626105910
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_53
timestamp 1626105910
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1626105910
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_29
timestamp 1626105910
transform 1 0 3772 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1626105910
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1626105910
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1626105910
transform -1 0 2116 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1626105910
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1626105910
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_17
timestamp 1626105910
transform 1 0 2668 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1626105910
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1626105910
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_11
timestamp 1626105910
transform 1 0 2116 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1626105910
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_A
timestamp 1626105910
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1626105910
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1626105910
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1626105910
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1626105910
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1626105910
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1626105910
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1626105910
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1626105910
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1626105910
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1626105910
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1626105910
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1626105910
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1626105910
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1626105910
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1626105910
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1626105910
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1626105910
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1626105910
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1626105910
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1626105910
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1626105910
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1626105910
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_100
timestamp 1626105910
transform 1 0 10304 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_111
timestamp 1626105910
transform 1 0 11316 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1626105910
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1626105910
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_106
timestamp 1626105910
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_99
timestamp 1626105910
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_87
timestamp 1626105910
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1626105910
transform 1 0 9752 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1626105910
transform 1 0 8648 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1626105910
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1626105910
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1626105910
transform 1 0 7544 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_78
timestamp 1626105910
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1626105910
transform 1 0 11776 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_112
timestamp 1626105910
transform 1 0 11408 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_111
timestamp 1626105910
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_99
timestamp 1626105910
transform 1 0 10212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1626105910
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1626105910
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1626105910
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1626105910
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_88
timestamp 1626105910
transform 1 0 9200 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1626105910
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1626105910
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1626105910
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1626105910
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1626105910
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1626105910
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1626105910
transform 1 0 9108 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1626105910
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1626105910
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1626105910
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1626105910
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1626105910
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_78
timestamp 1626105910
transform 1 0 8280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_83
timestamp 1626105910
transform 1 0 8740 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_71
timestamp 1626105910
transform 1 0 7636 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1626105910
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1626105910
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1626105910
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1626105910
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1626105910
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1626105910
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1626105910
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1626105910
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1626105910
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1626105910
transform 1 0 6072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_58
timestamp 1626105910
transform 1 0 6440 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1626105910
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1626105910
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1626105910
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1626105910
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1626105910
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_59
timestamp 1626105910
transform 1 0 6532 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1626105910
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1626105910
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1626105910
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1626105910
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1626105910
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1626105910
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1626105910
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1626105910
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1626105910
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1626105910
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_74
timestamp 1626105910
transform 1 0 7912 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_62
timestamp 1626105910
transform 1 0 6808 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1626105910
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_44
timestamp 1626105910
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_50
timestamp 1626105910
transform 1 0 5704 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1626105910
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A2
timestamp 1626105910
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_56
timestamp 1626105910
transform 1 0 6256 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_38
timestamp 1626105910
transform 1 0 4600 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_30
timestamp 1626105910
transform 1 0 3864 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_38
timestamp 1626105910
transform 1 0 4600 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_32
timestamp 1626105910
transform 1 0 4048 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__B2
timestamp 1626105910
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A1
timestamp 1626105910
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _097_
timestamp 1626105910
transform 1 0 3404 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1626105910
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1626105910
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1626105910
transform 1 0 3036 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1626105910
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1626105910
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1626105910
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1626105910
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1626105910
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1626105910
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__B1
timestamp 1626105910
transform -1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1626105910
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1626105910
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1626105910
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B2
timestamp 1626105910
transform 1 0 18124 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_184
timestamp 1626105910
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1626105910
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_180
timestamp 1626105910
transform 1 0 17664 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1626105910
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1626105910
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1626105910
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1626105910
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1626105910
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1626105910
transform 1 0 16928 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1626105910
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1626105910
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1626105910
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1626105910
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1626105910
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1626105910
transform -1 0 18952 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _091_
timestamp 1626105910
transform -1 0 18308 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1626105910
transform 1 0 18308 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1626105910
transform 1 0 17296 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B1
timestamp 1626105910
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1626105910
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_168
timestamp 1626105910
transform 1 0 16560 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1626105910
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1626105910
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1626105910
transform -1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1626105910
transform 1 0 18308 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1626105910
transform 1 0 17756 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_175
timestamp 1626105910
transform 1 0 17204 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__CLK
timestamp 1626105910
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__D
timestamp 1626105910
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A1
timestamp 1626105910
transform 1 0 18124 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1626105910
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_172
timestamp 1626105910
transform 1 0 16928 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1626105910
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1626105910
transform 1 0 15548 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__B
timestamp 1626105910
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1626105910
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A2
timestamp 1626105910
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _095_
timestamp 1626105910
transform -1 0 15548 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_142
timestamp 1626105910
transform 1 0 14168 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__CLK
timestamp 1626105910
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1626105910
transform -1 0 18952 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1626105910
transform -1 0 18952 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1626105910
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_190
timestamp 1626105910
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1626105910
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1626105910
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_167
timestamp 1626105910
transform 1 0 16468 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_155
timestamp 1626105910
transform 1 0 15364 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_143
timestamp 1626105910
transform 1 0 14260 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1626105910
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__CLK
timestamp 1626105910
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1626105910
transform -1 0 18952 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_190
timestamp 1626105910
transform 1 0 18584 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_182
timestamp 1626105910
transform 1 0 17848 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_176
timestamp 1626105910
transform 1 0 17296 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1626105910
transform 1 0 16744 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__CLK
timestamp 1626105910
transform 1 0 17664 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__RESET_B
timestamp 1626105910
transform 1 0 17112 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _101_
timestamp 1626105910
transform 1 0 14812 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1626105910
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1626105910
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1626105910
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1626105910
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_148
timestamp 1626105910
transform 1 0 14720 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1626105910
transform -1 0 18952 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_184
timestamp 1626105910
transform 1 0 18032 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_190
timestamp 1626105910
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1626105910
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1626105910
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_165
timestamp 1626105910
transform 1 0 16284 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_153
timestamp 1626105910
transform 1 0 15180 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_141
timestamp 1626105910
transform 1 0 14076 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__D
timestamp 1626105910
transform -1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1626105910
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1626105910
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1626105910
transform -1 0 18952 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1626105910
transform 1 0 18308 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _111_
timestamp 1626105910
transform -1 0 18308 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_22_163
timestamp 1626105910
transform 1 0 16100 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1626105910
transform 1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__C
timestamp 1626105910
transform -1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1626105910
transform 1 0 16652 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_160
timestamp 1626105910
transform 1 0 15824 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1626105910
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1626105910
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1626105910
transform -1 0 18952 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1626105910
transform -1 0 18952 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _083_
timestamp 1626105910
transform 1 0 17664 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_187
timestamp 1626105910
transform 1 0 18308 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_188
timestamp 1626105910
transform 1 0 18400 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_176
timestamp 1626105910
transform 1 0 17296 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_178
timestamp 1626105910
transform 1 0 17480 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A1
timestamp 1626105910
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1626105910
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1626105910
transform 1 0 18308 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_146
timestamp 1626105910
transform 1 0 14536 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1626105910
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1626105910
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1626105910
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_156
timestamp 1626105910
transform 1 0 15456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1626105910
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1626105910
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1626105910
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1626105910
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _118_
timestamp 1626105910
transform -1 0 18952 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_40_168
timestamp 1626105910
transform 1 0 16560 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_174
timestamp 1626105910
transform 1 0 17112 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1626105910
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1626105910
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1626105910
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1626105910
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1626105910
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1626105910
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1626105910
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_135
timestamp 1626105910
transform 1 0 13524 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1626105910
transform 1 0 13524 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1626105910
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1626105910
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1626105910
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_163
timestamp 1626105910
transform 1 0 16100 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_151
timestamp 1626105910
transform 1 0 14996 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_139
timestamp 1626105910
transform 1 0 13892 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1626105910
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_175
timestamp 1626105910
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1626105910
transform 1 0 17112 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1626105910
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1626105910
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1626105910
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1626105910
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_151
timestamp 1626105910
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1626105910
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1626105910
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1626105910
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1626105910
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1626105910
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1626105910
transform 1 0 16744 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_158
timestamp 1626105910
transform 1 0 15640 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1626105910
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1626105910
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1626105910
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1626105910
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_163
timestamp 1626105910
transform 1 0 16100 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1626105910
transform 1 0 15456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_144
timestamp 1626105910
transform 1 0 14352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1626105910
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1626105910
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1626105910
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1626105910
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_251
timestamp 1626105910
transform 1 0 24196 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1626105910
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1626105910
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1626105910
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_203
timestamp 1626105910
transform 1 0 19780 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1626105910
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_245
timestamp 1626105910
transform 1 0 23644 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__CLK
timestamp 1626105910
transform -1 0 19780 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1626105910
transform 1 0 23276 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_229
timestamp 1626105910
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1626105910
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1626105910
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1626105910
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1626105910
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1626105910
transform 1 0 22540 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1626105910
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_249
timestamp 1626105910
transform 1 0 24012 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1626105910
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_225
timestamp 1626105910
transform 1 0 21804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1626105910
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1626105910
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1626105910
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1626105910
transform 1 0 20700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1626105910
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_220
timestamp 1626105910
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1626105910
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1626105910
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1626105910
transform 1 0 22448 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1626105910
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1626105910
transform 1 0 22080 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1626105910
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1626105910
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1626105910
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1626105910
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1626105910
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1626105910
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1626105910
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_216
timestamp 1626105910
transform 1 0 20976 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1626105910
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1626105910
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1626105910
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1626105910
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_220
timestamp 1626105910
transform 1 0 21344 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1626105910
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_204
timestamp 1626105910
transform 1 0 19872 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1626105910
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_249
timestamp 1626105910
transform 1 0 24012 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1626105910
transform 1 0 22908 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_225
timestamp 1626105910
transform 1 0 21804 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_213
timestamp 1626105910
transform 1 0 20700 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1626105910
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1626105910
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1626105910
transform 1 0 19780 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1626105910
transform 1 0 23276 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_229
timestamp 1626105910
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1626105910
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1626105910
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1626105910
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1626105910
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_199
timestamp 1626105910
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_194
timestamp 1626105910
transform 1 0 18952 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1626105910
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1626105910
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_192
timestamp 1626105910
transform 1 0 18768 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_192
timestamp 1626105910
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1626105910
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_192
timestamp 1626105910
transform 1 0 18768 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1626105910
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1626105910
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_188
timestamp 1626105910
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1626105910
transform -1 0 18952 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1626105910
transform -1 0 18952 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_184
timestamp 1626105910
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_190
timestamp 1626105910
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1626105910
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1626105910
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1626105910
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1626105910
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_180
timestamp 1626105910
transform 1 0 17664 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1626105910
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1626105910
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1626105910
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1626105910
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1626105910
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_135
timestamp 1626105910
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1626105910
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1626105910
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1626105910
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1626105910
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _103_
timestamp 1626105910
transform 1 0 12052 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1626105910
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1626105910
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1626105910
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1626105910
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1626105910
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1626105910
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1626105910
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1626105910
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1626105910
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1626105910
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1626105910
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1626105910
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1626105910
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1626105910
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1626105910
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1626105910
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1626105910
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1626105910
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_124
timestamp 1626105910
transform 1 0 12512 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1626105910
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_122
timestamp 1626105910
transform 1 0 12328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1626105910
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1626105910
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1626105910
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1626105910
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1626105910
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1626105910
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1626105910
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1626105910
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1626105910
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1626105910
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1626105910
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1626105910
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1626105910
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1626105910
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1626105910
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_129
timestamp 1626105910
transform 1 0 12972 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1626105910
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1626105910
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_123
timestamp 1626105910
transform 1 0 12420 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1626105910
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1626105910
transform 1 0 12420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_127
timestamp 1626105910
transform 1 0 12788 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1626105910
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1626105910
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1626105910
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1626105910
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1626105910
transform 1 0 12420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1626105910
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _117_
timestamp 1626105910
transform -1 0 13892 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_27_127
timestamp 1626105910
transform 1 0 12788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1626105910
transform -1 0 18952 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1626105910
transform 1 0 18308 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1626105910
transform 1 0 17756 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A2
timestamp 1626105910
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B1
timestamp 1626105910
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_167
timestamp 1626105910
transform 1 0 16468 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_156
timestamp 1626105910
transform 1 0 15456 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 1626105910
transform 1 0 15916 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__D
timestamp 1626105910
transform -1 0 16468 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1626105910
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1626105910
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1626105910
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_243
timestamp 1626105910
transform 1 0 23460 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_249
timestamp 1626105910
transform 1 0 24012 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_231
timestamp 1626105910
transform 1 0 22356 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1626105910
transform 1 0 23276 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_229
timestamp 1626105910
transform 1 0 22172 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1626105910
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1626105910
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1626105910
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1626105910
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_225
timestamp 1626105910
transform 1 0 21804 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_237
timestamp 1626105910
transform 1 0 22908 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_225
timestamp 1626105910
transform 1 0 21804 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B2
timestamp 1626105910
transform 1 0 22172 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_213
timestamp 1626105910
transform 1 0 20700 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_213
timestamp 1626105910
transform 1 0 20700 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_201
timestamp 1626105910
transform 1 0 19596 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1626105910
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1626105910
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_201
timestamp 1626105910
transform 1 0 19596 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1626105910
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1626105910
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_249
timestamp 1626105910
transform 1 0 24012 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_237
timestamp 1626105910
transform 1 0 22908 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_225
timestamp 1626105910
transform 1 0 21804 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1626105910
transform 1 0 23276 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_229
timestamp 1626105910
transform 1 0 22172 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1626105910
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_213
timestamp 1626105910
transform 1 0 20700 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1626105910
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_220
timestamp 1626105910
transform 1 0 21344 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1626105910
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1626105910
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1626105910
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1626105910
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_225
timestamp 1626105910
transform 1 0 21804 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_245
timestamp 1626105910
transform 1 0 23644 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1626105910
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A2
timestamp 1626105910
transform 1 0 22356 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1626105910
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1626105910
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1626105910
transform 1 0 23828 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A1
timestamp 1626105910
transform 1 0 24196 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _088_
timestamp 1626105910
transform 1 0 22540 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1626105910
transform 1 0 22540 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1626105910
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1626105910
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_201
timestamp 1626105910
transform 1 0 19596 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1626105910
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_249
timestamp 1626105910
transform 1 0 24012 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_241
timestamp 1626105910
transform 1 0 23276 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1626105910
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1626105910
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1626105910
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_220
timestamp 1626105910
transform 1 0 21344 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1626105910
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_241
timestamp 1626105910
transform 1 0 23276 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_229
timestamp 1626105910
transform 1 0 22172 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B1
timestamp 1626105910
transform 1 0 23644 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1626105910
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_220
timestamp 1626105910
transform 1 0 21344 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1626105910
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1626105910
transform 1 0 22908 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1626105910
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_255
timestamp 1626105910
transform 1 0 24564 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1626105910
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1626105910
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1626105910
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_135
timestamp 1626105910
transform 1 0 13524 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1626105910
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_163
timestamp 1626105910
transform 1 0 16100 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1626105910
transform 1 0 16928 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1626105910
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_163
timestamp 1626105910
transform 1 0 16100 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1626105910
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1626105910
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1626105910
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1626105910
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_151
timestamp 1626105910
transform 1 0 14996 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1626105910
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_135
timestamp 1626105910
transform 1 0 13524 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_139
timestamp 1626105910
transform 1 0 13892 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1626105910
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_180
timestamp 1626105910
transform 1 0 17664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_168
timestamp 1626105910
transform 1 0 16560 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_135
timestamp 1626105910
transform 1 0 13524 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_172
timestamp 1626105910
transform 1 0 16928 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_163
timestamp 1626105910
transform 1 0 16100 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_156
timestamp 1626105910
transform 1 0 15456 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_144
timestamp 1626105910
transform 1 0 14352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_151
timestamp 1626105910
transform 1 0 14996 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_139
timestamp 1626105910
transform 1 0 13892 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1626105910
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_168
timestamp 1626105910
transform 1 0 16560 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_180
timestamp 1626105910
transform 1 0 17664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_168
timestamp 1626105910
transform 1 0 16560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_156
timestamp 1626105910
transform 1 0 15456 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_144
timestamp 1626105910
transform 1 0 14352 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1626105910
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_135
timestamp 1626105910
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_156
timestamp 1626105910
transform 1 0 15456 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_151
timestamp 1626105910
transform 1 0 14996 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1626105910
transform 1 0 17664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_168
timestamp 1626105910
transform 1 0 16560 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_139
timestamp 1626105910
transform 1 0 13892 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_172
timestamp 1626105910
transform 1 0 16928 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1626105910
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_163
timestamp 1626105910
transform 1 0 16100 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_156
timestamp 1626105910
transform 1 0 15456 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_144
timestamp 1626105910
transform 1 0 14352 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_144
timestamp 1626105910
transform 1 0 14352 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1626105910
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1626105910
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_135
timestamp 1626105910
transform 1 0 13524 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_180
timestamp 1626105910
transform 1 0 17664 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1626105910
transform 1 0 16928 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1626105910
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_140
timestamp 1626105910
transform 1 0 13984 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 1626105910
transform 1 0 13248 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_163
timestamp 1626105910
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1626105910
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1626105910
transform 1 0 17664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_168
timestamp 1626105910
transform 1 0 16560 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_162
timestamp 1626105910
transform 1 0 16008 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__A
timestamp 1626105910
transform 1 0 16376 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_135
timestamp 1626105910
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _054_
timestamp 1626105910
transform -1 0 16008 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_144
timestamp 1626105910
transform 1 0 14352 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_172
timestamp 1626105910
transform 1 0 16928 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_157
timestamp 1626105910
transform 1 0 15548 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1626105910
transform 1 0 16652 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1626105910
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_145
timestamp 1626105910
transform 1 0 14444 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1626105910
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1626105910
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_139
timestamp 1626105910
transform 1 0 13892 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1626105910
transform 1 0 16928 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1626105910
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_163
timestamp 1626105910
transform 1 0 16100 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_151
timestamp 1626105910
transform 1 0 14996 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_139
timestamp 1626105910
transform 1 0 13892 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1626105910
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_168
timestamp 1626105910
transform 1 0 16560 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1626105910
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1626105910
transform 1 0 16928 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1626105910
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_156
timestamp 1626105910
transform 1 0 15456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_135
timestamp 1626105910
transform 1 0 13524 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_135
timestamp 1626105910
transform 1 0 13524 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_180
timestamp 1626105910
transform 1 0 17664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_144
timestamp 1626105910
transform 1 0 14352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1626105910
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_133
timestamp 1626105910
transform 1 0 13340 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_168
timestamp 1626105910
transform 1 0 16560 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1626105910
transform 1 0 16928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1626105910
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_163
timestamp 1626105910
transform 1 0 16100 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_156
timestamp 1626105910
transform 1 0 15456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_144
timestamp 1626105910
transform 1 0 14352 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1626105910
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_139
timestamp 1626105910
transform 1 0 13892 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1626105910
transform 1 0 14260 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A1
timestamp 1626105910
transform 1 0 13156 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1626105910
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_163
timestamp 1626105910
transform 1 0 16100 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_156
timestamp 1626105910
transform 1 0 15456 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1626105910
transform 1 0 14352 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_180
timestamp 1626105910
transform 1 0 17664 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1626105910
transform 1 0 14996 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_139
timestamp 1626105910
transform 1 0 13892 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1626105910
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_180
timestamp 1626105910
transform 1 0 17664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1626105910
transform 1 0 16928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1626105910
transform 1 0 16560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1626105910
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1626105910
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1626105910
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_201
timestamp 1626105910
transform 1 0 19596 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1626105910
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1626105910
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_241
timestamp 1626105910
transform 1 0 23276 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_229
timestamp 1626105910
transform 1 0 22172 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1626105910
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_220
timestamp 1626105910
transform 1 0 21344 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1626105910
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1626105910
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_213
timestamp 1626105910
transform 1 0 20700 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1626105910
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_249
timestamp 1626105910
transform 1 0 24012 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_237
timestamp 1626105910
transform 1 0 22908 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1626105910
transform 1 0 24748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_237
timestamp 1626105910
transform 1 0 22908 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_225
timestamp 1626105910
transform 1 0 21804 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_241
timestamp 1626105910
transform 1 0 23276 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_249
timestamp 1626105910
transform 1 0 24012 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_225
timestamp 1626105910
transform 1 0 21804 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_229
timestamp 1626105910
transform 1 0 22172 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1626105910
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_220
timestamp 1626105910
transform 1 0 21344 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_213
timestamp 1626105910
transform 1 0 20700 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_201
timestamp 1626105910
transform 1 0 19596 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1626105910
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1626105910
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1626105910
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_241
timestamp 1626105910
transform 1 0 23276 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_229
timestamp 1626105910
transform 1 0 22172 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_213
timestamp 1626105910
transform 1 0 20700 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_201
timestamp 1626105910
transform 1 0 19596 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1626105910
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_237
timestamp 1626105910
transform 1 0 22908 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_249
timestamp 1626105910
transform 1 0 24012 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_225
timestamp 1626105910
transform 1 0 21804 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_213
timestamp 1626105910
transform 1 0 20700 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1626105910
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1626105910
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1626105910
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1626105910
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_220
timestamp 1626105910
transform 1 0 21344 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1626105910
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1626105910
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1626105910
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1626105910
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_241
timestamp 1626105910
transform 1 0 23276 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_255
timestamp 1626105910
transform 1 0 24564 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_247
timestamp 1626105910
transform 1 0 23828 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_235
timestamp 1626105910
transform 1 0 22724 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_223
timestamp 1626105910
transform 1 0 21620 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_229
timestamp 1626105910
transform 1 0 22172 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1626105910
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_217
timestamp 1626105910
transform 1 0 21068 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1626105910
transform 1 0 21436 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_220
timestamp 1626105910
transform 1 0 21344 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1626105910
transform 1 0 20792 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_201
timestamp 1626105910
transform 1 0 19596 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_241
timestamp 1626105910
transform 1 0 23276 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_229
timestamp 1626105910
transform 1 0 22172 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1626105910
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_220
timestamp 1626105910
transform 1 0 21344 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1626105910
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1626105910
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1626105910
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1626105910
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_237
timestamp 1626105910
transform 1 0 22908 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_249
timestamp 1626105910
transform 1 0 24012 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_225
timestamp 1626105910
transform 1 0 21804 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_213
timestamp 1626105910
transform 1 0 20700 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1626105910
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1626105910
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_192
timestamp 1626105910
transform 1 0 18768 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1626105910
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1626105910
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_192
timestamp 1626105910
transform 1 0 18768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_192
timestamp 1626105910
transform 1 0 18768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_192
timestamp 1626105910
transform 1 0 18768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_241
timestamp 1626105910
transform 1 0 23276 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_229
timestamp 1626105910
transform 1 0 22172 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1626105910
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1626105910
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_220
timestamp 1626105910
transform 1 0 21344 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1626105910
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1626105910
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_192
timestamp 1626105910
transform 1 0 18768 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_172
timestamp 1626105910
transform 1 0 16928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1626105910
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_163
timestamp 1626105910
transform 1 0 16100 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_151
timestamp 1626105910
transform 1 0 14996 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_139
timestamp 1626105910
transform 1 0 13892 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1626105910
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_192
timestamp 1626105910
transform 1 0 18768 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1626105910
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1626105910
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_192
timestamp 1626105910
transform 1 0 18768 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_192
timestamp 1626105910
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1626105910
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1626105910
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_192
timestamp 1626105910
transform 1 0 18768 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_192
timestamp 1626105910
transform 1 0 18768 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_115
timestamp 1626105910
transform 1 0 11684 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1626105910
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1626105910
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_99
timestamp 1626105910
transform 1 0 10212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_111
timestamp 1626105910
transform 1 0 11316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_99
timestamp 1626105910
transform 1 0 10212 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1626105910
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1626105910
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1626105910
transform 1 0 7176 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_78
timestamp 1626105910
transform 1 0 8280 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_87
timestamp 1626105910
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1626105910
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1626105910
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1626105910
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_74
timestamp 1626105910
transform 1 0 7912 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_66
timestamp 1626105910
transform 1 0 7176 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1626105910
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1626105910
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1626105910
transform 1 0 11316 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_99
timestamp 1626105910
transform 1 0 10212 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_87
timestamp 1626105910
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1626105910
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_78
timestamp 1626105910
transform 1 0 8280 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_87
timestamp 1626105910
transform 1 0 9108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_66
timestamp 1626105910
transform 1 0 7176 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_78
timestamp 1626105910
transform 1 0 8280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_111
timestamp 1626105910
transform 1 0 11316 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1626105910
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_115
timestamp 1626105910
transform 1 0 11684 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1626105910
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1626105910
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_94
timestamp 1626105910
transform 1 0 9752 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_82
timestamp 1626105910
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_70
timestamp 1626105910
transform 1 0 7544 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_106
timestamp 1626105910
transform 1 0 10856 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1626105910
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1626105910
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1626105910
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_111
timestamp 1626105910
transform 1 0 11316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_99
timestamp 1626105910
transform 1 0 10212 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_87
timestamp 1626105910
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1626105910
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1626105910
transform 1 0 7176 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1626105910
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_115
timestamp 1626105910
transform 1 0 11684 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_94
timestamp 1626105910
transform 1 0 9752 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_82
timestamp 1626105910
transform 1 0 8648 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_70
timestamp 1626105910
transform 1 0 7544 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1626105910
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_82
timestamp 1626105910
transform 1 0 8648 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_70
timestamp 1626105910
transform 1 0 7544 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_99
timestamp 1626105910
transform 1 0 10212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_111
timestamp 1626105910
transform 1 0 11316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_31
timestamp 1626105910
transform 1 0 3956 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_27
timestamp 1626105910
transform 1 0 3588 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1626105910
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_32
timestamp 1626105910
transform 1 0 4048 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_25
timestamp 1626105910
transform 1 0 3404 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B2
timestamp 1626105910
transform 1 0 3772 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A1
timestamp 1626105910
transform 1 0 4416 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1626105910
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B1
timestamp 1626105910
transform 1 0 3864 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _090_
timestamp 1626105910
transform -1 0 3404 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1626105910
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1626105910
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1626105910
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1626105910
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1626105910
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1626105910
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1626105910
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_27
timestamp 1626105910
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1626105910
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1626105910
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_42
timestamp 1626105910
transform 1 0 4968 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_30
timestamp 1626105910
transform 1 0 3864 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1626105910
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1626105910
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1626105910
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1626105910
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1626105910
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_15
timestamp 1626105910
transform 1 0 2484 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1626105910
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1626105910
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1626105910
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1626105910
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1626105910
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1626105910
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1626105910
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1626105910
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_51
timestamp 1626105910
transform 1 0 5796 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1626105910
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1626105910
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1626105910
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1626105910
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1626105910
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1626105910
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1626105910
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1626105910
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1626105910
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1626105910
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1626105910
transform -1 0 2116 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_17
timestamp 1626105910
transform 1 0 2668 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1626105910
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_11
timestamp 1626105910
transform 1 0 2116 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1626105910
transform 1 0 1380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output9_A
timestamp 1626105910
transform 1 0 2484 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1626105910
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1626105910
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_45
timestamp 1626105910
transform 1 0 5244 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1626105910
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_33
timestamp 1626105910
transform 1 0 4140 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_27
timestamp 1626105910
transform 1 0 3588 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A2
timestamp 1626105910
transform 1 0 3956 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1626105910
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1626105910
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1626105910
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1626105910
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1626105910
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_51
timestamp 1626105910
transform 1 0 5796 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_50
timestamp 1626105910
transform 1 0 5704 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1626105910
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_43
timestamp 1626105910
transform 1 0 5060 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_55
timestamp 1626105910
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1626105910
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_38
timestamp 1626105910
transform 1 0 4600 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_23
timestamp 1626105910
transform 1 0 3220 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_15
timestamp 1626105910
transform 1 0 2484 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_21
timestamp 1626105910
transform 1 0 3036 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1626105910
transform 1 0 2484 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A1
timestamp 1626105910
transform -1 0 3220 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A3
timestamp 1626105910
transform 1 0 3404 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1626105910
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A2
timestamp 1626105910
transform 1 0 2852 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_2  _067_
timestamp 1626105910
transform 1 0 1656 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1626105910
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1626105910
transform 1 0 1380 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1626105910
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1626105910
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1626105910
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1626105910
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1626105910
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1626105910
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1626105910
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1626105910
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1626105910
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1626105910
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1626105910
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1626105910
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1626105910
transform 1 0 2484 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B1
timestamp 1626105910
transform 1 0 2852 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1626105910
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1626105910
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1626105910
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1626105910
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1626105910
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_33
timestamp 1626105910
transform 1 0 4140 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1626105910
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1626105910
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1626105910
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1626105910
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1626105910
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_42
timestamp 1626105910
transform 1 0 4968 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_30
timestamp 1626105910
transform 1 0 3864 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1626105910
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1626105910
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1626105910
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1626105910
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1626105910
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_27
timestamp 1626105910
transform 1 0 3588 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__C1
timestamp 1626105910
transform -1 0 4140 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1626105910
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1626105910
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1626105910
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_53
timestamp 1626105910
transform 1 0 5980 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_41
timestamp 1626105910
transform 1 0 4876 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_29
timestamp 1626105910
transform 1 0 3772 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1626105910
transform 1 0 6348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1626105910
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_51
timestamp 1626105910
transform 1 0 5796 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1626105910
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1626105910
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1626105910
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1626105910
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1626105910
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1626105910
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_51
timestamp 1626105910
transform 1 0 5796 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1626105910
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1626105910
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1626105910
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1626105910
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_17
timestamp 1626105910
transform 1 0 2668 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output10_A
timestamp 1626105910
transform -1 0 2668 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1626105910
transform -1 0 2116 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1626105910
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_11
timestamp 1626105910
transform 1 0 2116 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1626105910
transform 1 0 1380 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_21
timestamp 1626105910
transform 1 0 3036 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_45
timestamp 1626105910
transform 1 0 5244 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1626105910
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1626105910
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1626105910
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_51
timestamp 1626105910
transform 1 0 5796 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1626105910
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1626105910
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1626105910
transform 1 0 3588 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1626105910
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_82
timestamp 1626105910
transform 1 0 8648 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_70
timestamp 1626105910
transform 1 0 7544 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1626105910
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_78
timestamp 1626105910
transform 1 0 8280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_111
timestamp 1626105910
transform 1 0 11316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1626105910
transform 1 0 10212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1626105910
transform 1 0 9108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1626105910
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_78
timestamp 1626105910
transform 1 0 8280 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_66
timestamp 1626105910
transform 1 0 7176 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_66
timestamp 1626105910
transform 1 0 7176 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_115
timestamp 1626105910
transform 1 0 11684 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1626105910
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_106
timestamp 1626105910
transform 1 0 10856 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1626105910
transform 1 0 9752 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_111
timestamp 1626105910
transform 1 0 11316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_99
timestamp 1626105910
transform 1 0 10212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1626105910
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1626105910
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1626105910
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1626105910
transform 1 0 8648 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1626105910
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_70
timestamp 1626105910
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_111
timestamp 1626105910
transform 1 0 11316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_115
timestamp 1626105910
transform 1 0 11684 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_115
timestamp 1626105910
transform 1 0 11684 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1626105910
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_106
timestamp 1626105910
transform 1 0 10856 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1626105910
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_82
timestamp 1626105910
transform 1 0 8648 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_70
timestamp 1626105910
transform 1 0 7544 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1626105910
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_106
timestamp 1626105910
transform 1 0 10856 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_111
timestamp 1626105910
transform 1 0 11316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_115
timestamp 1626105910
transform 1 0 11684 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1626105910
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_106
timestamp 1626105910
transform 1 0 10856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_99
timestamp 1626105910
transform 1 0 10212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_94
timestamp 1626105910
transform 1 0 9752 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_87
timestamp 1626105910
transform 1 0 9108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_82
timestamp 1626105910
transform 1 0 8648 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1626105910
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_78
timestamp 1626105910
transform 1 0 8280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1626105910
transform 1 0 7176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_70
timestamp 1626105910
transform 1 0 7544 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_99
timestamp 1626105910
transform 1 0 10212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_94
timestamp 1626105910
transform 1 0 9752 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_78
timestamp 1626105910
transform 1 0 8280 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_108
timestamp 1626105910
transform 1 0 11040 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A
timestamp 1626105910
transform 1 0 10856 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  _058_
timestamp 1626105910
transform -1 0 10488 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_102
timestamp 1626105910
transform 1 0 10488 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_95
timestamp 1626105910
transform 1 0 9844 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1626105910
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_87
timestamp 1626105910
transform 1 0 9108 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1626105910
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1626105910
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_87
timestamp 1626105910
transform 1 0 9108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_82
timestamp 1626105910
transform 1 0 8648 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_115
timestamp 1626105910
transform 1 0 11684 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1626105910
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_106
timestamp 1626105910
transform 1 0 10856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1626105910
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_54
timestamp 1626105910
transform 1 0 6072 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_58
timestamp 1626105910
transform 1 0 6440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1626105910
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1626105910
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1626105910
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1626105910
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_115
timestamp 1626105910
transform 1 0 11684 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1626105910
transform 1 0 6072 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_54
timestamp 1626105910
transform 1 0 6072 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_58
timestamp 1626105910
transform 1 0 6440 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_62
timestamp 1626105910
transform 1 0 6808 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1626105910
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1626105910
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_58
timestamp 1626105910
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1626105910
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_51
timestamp 1626105910
transform 1 0 5796 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_70
timestamp 1626105910
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_106
timestamp 1626105910
transform 1 0 10856 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_94
timestamp 1626105910
transform 1 0 9752 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1626105910
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_58
timestamp 1626105910
transform 1 0 6440 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_82
timestamp 1626105910
transform 1 0 8648 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1626105910
transform 1 0 6072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_58
timestamp 1626105910
transform 1 0 6440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1626105910
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_54
timestamp 1626105910
transform 1 0 6072 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_58
timestamp 1626105910
transform 1 0 6440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1626105910
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_54
timestamp 1626105910
transform 1 0 6072 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_58
timestamp 1626105910
transform 1 0 6440 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_54
timestamp 1626105910
transform 1 0 6072 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_58
timestamp 1626105910
transform 1 0 6440 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_106
timestamp 1626105910
transform 1 0 10856 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_94
timestamp 1626105910
transform 1 0 9752 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_82
timestamp 1626105910
transform 1 0 8648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_70
timestamp 1626105910
transform 1 0 7544 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_111
timestamp 1626105910
transform 1 0 11316 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_99
timestamp 1626105910
transform 1 0 10212 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_87
timestamp 1626105910
transform 1 0 9108 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1626105910
transform 1 0 9016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_78
timestamp 1626105910
transform 1 0 8280 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_66
timestamp 1626105910
transform 1 0 7176 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_82
timestamp 1626105910
transform 1 0 8648 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_70
timestamp 1626105910
transform 1 0 7544 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_70
timestamp 1626105910
transform 1 0 7544 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1626105910
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_115
timestamp 1626105910
transform 1 0 11684 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1626105910
transform 1 0 11592 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_106
timestamp 1626105910
transform 1 0 10856 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_94
timestamp 1626105910
transform 1 0 9752 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_82
timestamp 1626105910
transform 1 0 8648 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1626105910
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_116
timestamp 1626105910
transform 1 0 11776 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_115
timestamp 1626105910
transform 1 0 11684 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_104
timestamp 1626105910
transform 1 0 10672 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1626105910
transform 1 0 11592 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_106
timestamp 1626105910
transform 1 0 10856 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_4  _080_
timestamp 1626105910
transform -1 0 10120 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_67_94
timestamp 1626105910
transform 1 0 9752 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_98
timestamp 1626105910
transform 1 0 10120 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1626105910
transform 1 0 10488 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_82
timestamp 1626105910
transform 1 0 8648 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1626105910
transform 1 0 9016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_80
timestamp 1626105910
transform 1 0 8464 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_87
timestamp 1626105910
transform 1 0 9108 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_70
timestamp 1626105910
transform 1 0 7544 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1626105910
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_106
timestamp 1626105910
transform 1 0 10856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_111
timestamp 1626105910
transform 1 0 11316 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_111
timestamp 1626105910
transform 1 0 11316 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_99
timestamp 1626105910
transform 1 0 10212 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_87
timestamp 1626105910
transform 1 0 9108 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1626105910
transform 1 0 9016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_78
timestamp 1626105910
transform 1 0 8280 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_66
timestamp 1626105910
transform 1 0 7176 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_99
timestamp 1626105910
transform 1 0 10212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_87
timestamp 1626105910
transform 1 0 9108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1626105910
transform 1 0 9016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_78
timestamp 1626105910
transform 1 0 8280 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_115
timestamp 1626105910
transform 1 0 11684 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_115
timestamp 1626105910
transform 1 0 11684 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1626105910
transform 1 0 11592 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_106
timestamp 1626105910
transform 1 0 10856 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_94
timestamp 1626105910
transform 1 0 9752 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_82
timestamp 1626105910
transform 1 0 8648 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_70
timestamp 1626105910
transform 1 0 7544 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_66
timestamp 1626105910
transform 1 0 7176 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_115
timestamp 1626105910
transform 1 0 11684 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1626105910
transform 1 0 11592 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1626105910
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1626105910
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1626105910
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_42
timestamp 1626105910
transform 1 0 4968 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_30
timestamp 1626105910
transform 1 0 3864 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_27
timestamp 1626105910
transform 1 0 3588 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1626105910
transform 1 0 3772 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1626105910
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1626105910
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1626105910
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_11
timestamp 1626105910
transform 1 0 2116 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1626105910
transform 1 0 6348 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1626105910
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1626105910
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1626105910
transform 1 0 6348 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1626105910
transform 1 0 6072 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  _084_
timestamp 1626105910
transform 1 0 5152 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1626105910
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_42
timestamp 1626105910
transform 1 0 4968 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_51
timestamp 1626105910
transform 1 0 5796 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_50
timestamp 1626105910
transform 1 0 5704 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1626105910
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_30
timestamp 1626105910
transform 1 0 3864 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_27
timestamp 1626105910
transform 1 0 3588 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1626105910
transform 1 0 3772 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1626105910
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1626105910
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1626105910
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1626105910
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1626105910
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1626105910
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1626105910
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1626105910
transform 1 0 6348 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1626105910
transform 1 0 6348 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1626105910
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_51
timestamp 1626105910
transform 1 0 5796 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1626105910
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1626105910
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1626105910
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1626105910
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_51
timestamp 1626105910
transform 1 0 5796 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1626105910
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1626105910
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_42
timestamp 1626105910
transform 1 0 4968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_51
timestamp 1626105910
transform 1 0 5796 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1626105910
transform 1 0 6348 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1626105910
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1626105910
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_17
timestamp 1626105910
transform 1 0 2668 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_51
timestamp 1626105910
transform 1 0 5796 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1626105910
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1626105910
transform -1 0 2116 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1626105910
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1626105910
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1626105910
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1626105910
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1626105910
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1626105910
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1626105910
transform 1 0 1380 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1626105910
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1626105910
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_42
timestamp 1626105910
transform 1 0 4968 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_30
timestamp 1626105910
transform 1 0 3864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_30
timestamp 1626105910
transform 1 0 3864 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output11_A
timestamp 1626105910
transform 1 0 2484 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_27
timestamp 1626105910
transform 1 0 3588 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1626105910
transform 1 0 3772 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1626105910
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_30
timestamp 1626105910
transform 1 0 3864 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_27
timestamp 1626105910
transform 1 0 3588 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1626105910
transform 1 0 3772 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1626105910
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1626105910
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1626105910
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_51
timestamp 1626105910
transform 1 0 5796 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1626105910
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1626105910
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1626105910
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1626105910
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1626105910
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_51
timestamp 1626105910
transform 1 0 5796 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1626105910
transform 1 0 6348 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1626105910
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_51
timestamp 1626105910
transform 1 0 5796 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1626105910
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1626105910
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1626105910
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1626105910
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1626105910
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1626105910
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1626105910
transform 1 0 6348 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1626105910
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1626105910
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_42
timestamp 1626105910
transform 1 0 4968 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_30
timestamp 1626105910
transform 1 0 3864 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_42
timestamp 1626105910
transform 1 0 4968 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_42
timestamp 1626105910
transform 1 0 4968 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_30
timestamp 1626105910
transform 1 0 3864 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_42
timestamp 1626105910
transform 1 0 4968 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1626105910
transform 1 0 6440 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1626105910
transform 1 0 6348 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_51
timestamp 1626105910
transform 1 0 5796 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_54
timestamp 1626105910
transform 1 0 6072 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_30
timestamp 1626105910
transform 1 0 3864 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1626105910
transform 1 0 4692 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1626105910
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_30
timestamp 1626105910
transform 1 0 3864 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_27
timestamp 1626105910
transform 1 0 3588 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1626105910
transform 1 0 3772 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1626105910
transform 1 0 3772 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output13
timestamp 1626105910
transform -1 0 2116 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_17
timestamp 1626105910
transform 1 0 2668 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1626105910
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_11
timestamp 1626105910
transform 1 0 2116 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1626105910
transform 1 0 1380 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output13_A
timestamp 1626105910
transform 1 0 2484 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1626105910
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1626105910
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1626105910
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1626105910
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1626105910
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1626105910
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_27
timestamp 1626105910
transform 1 0 3588 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1626105910
transform 1 0 3772 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1626105910
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1626105910
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1626105910
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1626105910
transform 1 0 3772 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_17
timestamp 1626105910
transform 1 0 2668 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1626105910
transform 1 0 6348 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1626105910
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_51
timestamp 1626105910
transform 1 0 5796 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1626105910
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1626105910
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1626105910
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1626105910
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1626105910
transform 1 0 2484 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1626105910
transform -1 0 2116 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1626105910
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_11
timestamp 1626105910
transform 1 0 2116 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1626105910
transform 1 0 1380 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1626105910
transform 1 0 6348 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1626105910
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_42
timestamp 1626105910
transform 1 0 4968 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_70
timestamp 1626105910
transform 1 0 7544 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1626105910
transform 1 0 11592 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_111
timestamp 1626105910
transform 1 0 11316 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_99
timestamp 1626105910
transform 1 0 10212 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_87
timestamp 1626105910
transform 1 0 9108 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1626105910
transform 1 0 9016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_117
timestamp 1626105910
transform 1 0 11868 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_115
timestamp 1626105910
transform 1 0 11684 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_111
timestamp 1626105910
transform 1 0 11316 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1626105910
transform 1 0 11776 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1626105910
transform 1 0 11592 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_112
timestamp 1626105910
transform 1 0 11408 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_106
timestamp 1626105910
transform 1 0 10856 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_100
timestamp 1626105910
transform 1 0 10304 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_88
timestamp 1626105910
transform 1 0 9200 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_94
timestamp 1626105910
transform 1 0 9752 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_82
timestamp 1626105910
transform 1 0 8648 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_99
timestamp 1626105910
transform 1 0 10212 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_87
timestamp 1626105910
transform 1 0 9108 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1626105910
transform 1 0 9108 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1626105910
transform 1 0 9016 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_83
timestamp 1626105910
transform 1 0 8740 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1626105910
transform 1 0 7636 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_70
timestamp 1626105910
transform 1 0 7544 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_66
timestamp 1626105910
transform 1 0 7176 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_78
timestamp 1626105910
transform 1 0 8280 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_78
timestamp 1626105910
transform 1 0 8280 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_66
timestamp 1626105910
transform 1 0 7176 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_106
timestamp 1626105910
transform 1 0 10856 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_115
timestamp 1626105910
transform 1 0 11684 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1626105910
transform 1 0 11592 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_106
timestamp 1626105910
transform 1 0 10856 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_94
timestamp 1626105910
transform 1 0 9752 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_82
timestamp 1626105910
transform 1 0 8648 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_70
timestamp 1626105910
transform 1 0 7544 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_94
timestamp 1626105910
transform 1 0 9752 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_111
timestamp 1626105910
transform 1 0 11316 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_99
timestamp 1626105910
transform 1 0 10212 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_87
timestamp 1626105910
transform 1 0 9108 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1626105910
transform 1 0 9016 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_78
timestamp 1626105910
transform 1 0 8280 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_66
timestamp 1626105910
transform 1 0 7176 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_70
timestamp 1626105910
transform 1 0 7544 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_115
timestamp 1626105910
transform 1 0 11684 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1626105910
transform 1 0 11592 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_106
timestamp 1626105910
transform 1 0 10856 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_94
timestamp 1626105910
transform 1 0 9752 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_82
timestamp 1626105910
transform 1 0 8648 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_70
timestamp 1626105910
transform 1 0 7544 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_115
timestamp 1626105910
transform 1 0 11684 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_111
timestamp 1626105910
transform 1 0 11316 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_99
timestamp 1626105910
transform 1 0 10212 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_87
timestamp 1626105910
transform 1 0 9108 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1626105910
transform 1 0 9016 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_78
timestamp 1626105910
transform 1 0 8280 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_66
timestamp 1626105910
transform 1 0 7176 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_82
timestamp 1626105910
transform 1 0 8648 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_115
timestamp 1626105910
transform 1 0 11684 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1626105910
transform 1 0 11592 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_106
timestamp 1626105910
transform 1 0 10856 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_94
timestamp 1626105910
transform 1 0 9752 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_82
timestamp 1626105910
transform 1 0 8648 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_54
timestamp 1626105910
transform 1 0 6072 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_58
timestamp 1626105910
transform 1 0 6440 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_58
timestamp 1626105910
transform 1 0 6440 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1626105910
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_58
timestamp 1626105910
transform 1 0 6440 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_54
timestamp 1626105910
transform 1 0 6072 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_59
timestamp 1626105910
transform 1 0 6532 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_58
timestamp 1626105910
transform 1 0 6440 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_54
timestamp 1626105910
transform 1 0 6072 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_58
timestamp 1626105910
transform 1 0 6440 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_54
timestamp 1626105910
transform 1 0 6072 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_58
timestamp 1626105910
transform 1 0 6440 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_54
timestamp 1626105910
transform 1 0 6072 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_58
timestamp 1626105910
transform 1 0 6440 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_54
timestamp 1626105910
transform 1 0 6072 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_123
timestamp 1626105910
transform 1 0 12420 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_127
timestamp 1626105910
transform 1 0 12788 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_111
timestamp 1626105910
transform 1 0 11316 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_99
timestamp 1626105910
transform 1 0 10212 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_87
timestamp 1626105910
transform 1 0 9108 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_83
timestamp 1626105910
transform 1 0 8740 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1626105910
transform 1 0 9016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_71
timestamp 1626105910
transform 1 0 7636 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_65
timestamp 1626105910
transform 1 0 7084 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1626105910
transform 1 0 7452 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_4  _081_
timestamp 1626105910
transform -1 0 7084 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_73_58
timestamp 1626105910
transform 1 0 6440 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_54
timestamp 1626105910
transform 1 0 6072 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_42
timestamp 1626105910
transform 1 0 4968 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_30
timestamp 1626105910
transform 1 0 3864 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_27
timestamp 1626105910
transform 1 0 3588 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1626105910
transform 1 0 3772 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1626105910
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1626105910
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1626105910
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_58
timestamp 1626105910
transform 1 0 6440 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_54
timestamp 1626105910
transform 1 0 6072 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_58
timestamp 1626105910
transform 1 0 6440 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_196
timestamp 1626105910
transform 1 0 19136 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1626105910
transform 1 0 19504 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_241
timestamp 1626105910
transform 1 0 23276 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_229
timestamp 1626105910
transform 1 0 22172 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1626105910
transform 1 0 22080 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_220
timestamp 1626105910
transform 1 0 21344 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1626105910
transform 1 0 23276 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1626105910
transform 1 0 22172 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_216
timestamp 1626105910
transform 1 0 20976 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1626105910
transform 1 0 22080 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_204
timestamp 1626105910
transform 1 0 19872 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_201
timestamp 1626105910
transform 1 0 19596 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_241
timestamp 1626105910
transform 1 0 23276 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_201
timestamp 1626105910
transform 1 0 19596 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1626105910
transform 1 0 19504 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_229
timestamp 1626105910
transform 1 0 22172 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1626105910
transform 1 0 22080 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_220
timestamp 1626105910
transform 1 0 21344 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_208
timestamp 1626105910
transform 1 0 20240 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_196
timestamp 1626105910
transform 1 0 19136 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1626105910
transform 1 0 19504 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_208
timestamp 1626105910
transform 1 0 20240 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1626105910
transform 1 0 24748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_256
timestamp 1626105910
transform 1 0 24656 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_252
timestamp 1626105910
transform 1 0 24288 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_246
timestamp 1626105910
transform 1 0 23736 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_240
timestamp 1626105910
transform 1 0 23184 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A1
timestamp 1626105910
transform 1 0 24104 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B1
timestamp 1626105910
transform 1 0 23552 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_1  _079_
timestamp 1626105910
transform 1 0 22448 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_228
timestamp 1626105910
transform 1 0 22080 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A3
timestamp 1626105910
transform 1 0 21896 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_225
timestamp 1626105910
transform 1 0 21804 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_213
timestamp 1626105910
transform 1 0 20700 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_196
timestamp 1626105910
transform 1 0 19136 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1626105910
transform 1 0 24748 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_237
timestamp 1626105910
transform 1 0 22908 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_249
timestamp 1626105910
transform 1 0 24012 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1626105910
transform 1 0 24748 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_237
timestamp 1626105910
transform 1 0 22908 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1626105910
transform 1 0 24748 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_249
timestamp 1626105910
transform 1 0 24012 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1626105910
transform -1 0 24748 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_237
timestamp 1626105910
transform 1 0 22908 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1626105910
transform 1 0 21804 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_241
timestamp 1626105910
transform 1 0 23276 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A2
timestamp 1626105910
transform 1 0 23552 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_246
timestamp 1626105910
transform 1 0 23736 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_249
timestamp 1626105910
transform 1 0 24012 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_213
timestamp 1626105910
transform 1 0 20700 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_229
timestamp 1626105910
transform 1 0 22172 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_225
timestamp 1626105910
transform 1 0 21804 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_213
timestamp 1626105910
transform 1 0 20700 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_225
timestamp 1626105910
transform 1 0 21804 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1626105910
transform 1 0 22080 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_220
timestamp 1626105910
transform 1 0 21344 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_208
timestamp 1626105910
transform 1 0 20240 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_213
timestamp 1626105910
transform 1 0 20700 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_201
timestamp 1626105910
transform 1 0 19596 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1626105910
transform 1 0 19504 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_196
timestamp 1626105910
transform 1 0 19136 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_201
timestamp 1626105910
transform 1 0 19596 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_241
timestamp 1626105910
transform 1 0 23276 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_229
timestamp 1626105910
transform 1 0 22172 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1626105910
transform 1 0 22080 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_220
timestamp 1626105910
transform 1 0 21344 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_208
timestamp 1626105910
transform 1 0 20240 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_180
timestamp 1626105910
transform 1 0 17664 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_182
timestamp 1626105910
transform 1 0 17848 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_168
timestamp 1626105910
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_156
timestamp 1626105910
transform 1 0 15456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_144
timestamp 1626105910
transform 1 0 14352 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1626105910
transform 1 0 14260 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_172
timestamp 1626105910
transform 1 0 16928 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_180
timestamp 1626105910
transform 1 0 17664 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__CLK
timestamp 1626105910
transform 1 0 17480 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1626105910
transform 1 0 16836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_174
timestamp 1626105910
transform 1 0 17112 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_167
timestamp 1626105910
transform 1 0 16468 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__D
timestamp 1626105910
transform -1 0 17112 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _113_
timestamp 1626105910
transform -1 0 16468 0 1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_63_147
timestamp 1626105910
transform 1 0 14628 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_151
timestamp 1626105910
transform 1 0 14996 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_139
timestamp 1626105910
transform 1 0 13892 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_172
timestamp 1626105910
transform 1 0 16928 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1626105910
transform 1 0 16836 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_170
timestamp 1626105910
transform 1 0 16744 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_164
timestamp 1626105910
transform 1 0 16192 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_165
timestamp 1626105910
transform 1 0 16284 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__A
timestamp 1626105910
transform 1 0 16560 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  _053_
timestamp 1626105910
transform -1 0 16192 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_153
timestamp 1626105910
transform 1 0 15180 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_152
timestamp 1626105910
transform 1 0 15088 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1626105910
transform 1 0 14260 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_144
timestamp 1626105910
transform 1 0 14352 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_135
timestamp 1626105910
transform 1 0 13524 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_135
timestamp 1626105910
transform 1 0 13524 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_135
timestamp 1626105910
transform 1 0 13524 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_135
timestamp 1626105910
transform 1 0 13524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A2
timestamp 1626105910
transform -1 0 13524 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_141
timestamp 1626105910
transform 1 0 14076 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_180
timestamp 1626105910
transform 1 0 17664 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B
timestamp 1626105910
transform 1 0 13892 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_172
timestamp 1626105910
transform 1 0 16928 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_168
timestamp 1626105910
transform 1 0 16560 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1626105910
transform 1 0 16836 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_163
timestamp 1626105910
transform 1 0 16100 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_151
timestamp 1626105910
transform 1 0 14996 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_139
timestamp 1626105910
transform 1 0 13892 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_156
timestamp 1626105910
transform 1 0 15456 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_144
timestamp 1626105910
transform 1 0 14352 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_140
timestamp 1626105910
transform 1 0 13984 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1626105910
transform 1 0 14260 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_180
timestamp 1626105910
transform 1 0 17664 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_172
timestamp 1626105910
transform 1 0 16928 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1626105910
transform 1 0 16836 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_163
timestamp 1626105910
transform 1 0 16100 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_151
timestamp 1626105910
transform 1 0 14996 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_139
timestamp 1626105910
transform 1 0 13892 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1626105910
transform 1 0 16836 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_168
timestamp 1626105910
transform 1 0 16560 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_156
timestamp 1626105910
transform 1 0 15456 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_144
timestamp 1626105910
transform 1 0 14352 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1626105910
transform 1 0 14260 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_163
timestamp 1626105910
transform 1 0 16100 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1626105910
transform 1 0 16836 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_163
timestamp 1626105910
transform 1 0 16100 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_151
timestamp 1626105910
transform 1 0 14996 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_139
timestamp 1626105910
transform 1 0 13892 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_172
timestamp 1626105910
transform 1 0 16928 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1626105910
transform 1 0 16836 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_163
timestamp 1626105910
transform 1 0 16100 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_151
timestamp 1626105910
transform 1 0 14996 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_139
timestamp 1626105910
transform 1 0 13892 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_156
timestamp 1626105910
transform 1 0 15456 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_144
timestamp 1626105910
transform 1 0 14352 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_180
timestamp 1626105910
transform 1 0 17664 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1626105910
transform 1 0 14260 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_168
timestamp 1626105910
transform 1 0 16560 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_156
timestamp 1626105910
transform 1 0 15456 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_144
timestamp 1626105910
transform 1 0 14352 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_180
timestamp 1626105910
transform 1 0 17664 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1626105910
transform 1 0 14260 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_168
timestamp 1626105910
transform 1 0 16560 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_156
timestamp 1626105910
transform 1 0 15456 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_144
timestamp 1626105910
transform 1 0 14352 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1626105910
transform 1 0 14260 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_163
timestamp 1626105910
transform 1 0 16100 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1626105910
transform 1 0 17664 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_172
timestamp 1626105910
transform 1 0 16928 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_151
timestamp 1626105910
transform 1 0 14996 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_139
timestamp 1626105910
transform 1 0 13892 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_175
timestamp 1626105910
transform 1 0 17204 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_158
timestamp 1626105910
transform 1 0 15640 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_172
timestamp 1626105910
transform 1 0 16928 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1626105910
transform 1 0 16560 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1626105910
transform 1 0 17112 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1626105910
transform 1 0 16836 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_170
timestamp 1626105910
transform 1 0 16744 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_163
timestamp 1626105910
transform 1 0 16100 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_146
timestamp 1626105910
transform 1 0 14536 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_151
timestamp 1626105910
transform 1 0 14996 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_139
timestamp 1626105910
transform 1 0 13892 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1626105910
transform 1 0 15456 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1626105910
transform 1 0 14352 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1626105910
transform 1 0 14444 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1626105910
transform 1 0 14260 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1626105910
transform 1 0 14076 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_135
timestamp 1626105910
transform 1 0 13524 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_180
timestamp 1626105910
transform 1 0 17664 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_135
timestamp 1626105910
transform 1 0 13524 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_135
timestamp 1626105910
transform 1 0 13524 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_135
timestamp 1626105910
transform 1 0 13524 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1626105910
transform 1 0 16836 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_168
timestamp 1626105910
transform 1 0 16560 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_172
timestamp 1626105910
transform 1 0 16928 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1626105910
transform 1 0 16836 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_163
timestamp 1626105910
transform 1 0 16100 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_151
timestamp 1626105910
transform 1 0 14996 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_139
timestamp 1626105910
transform 1 0 13892 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_172
timestamp 1626105910
transform 1 0 16928 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_229
timestamp 1626105910
transform 1 0 22172 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1626105910
transform 1 0 24748 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_245
timestamp 1626105910
transform 1 0 23644 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1626105910
transform 1 0 24748 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_249
timestamp 1626105910
transform 1 0 24012 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_233
timestamp 1626105910
transform 1 0 22540 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_241
timestamp 1626105910
transform 1 0 23276 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_229
timestamp 1626105910
transform 1 0 22172 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_237
timestamp 1626105910
transform 1 0 22908 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_225
timestamp 1626105910
transform 1 0 21804 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1626105910
transform 1 0 22448 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1626105910
transform 1 0 22080 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_228
timestamp 1626105910
transform 1 0 22080 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_216
timestamp 1626105910
transform 1 0 20976 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_204
timestamp 1626105910
transform 1 0 19872 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_208
timestamp 1626105910
transform 1 0 20240 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_213
timestamp 1626105910
transform 1 0 20700 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_201
timestamp 1626105910
transform 1 0 19596 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1626105910
transform 1 0 19780 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_220
timestamp 1626105910
transform 1 0 21344 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_237
timestamp 1626105910
transform 1 0 22908 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_196
timestamp 1626105910
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_249
timestamp 1626105910
transform 1 0 24012 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1626105910
transform 1 0 19504 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_199
timestamp 1626105910
transform 1 0 19412 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_225
timestamp 1626105910
transform 1 0 21804 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_213
timestamp 1626105910
transform 1 0 20700 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_201
timestamp 1626105910
transform 1 0 19596 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1626105910
transform 1 0 19504 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_196
timestamp 1626105910
transform 1 0 19136 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_254
timestamp 1626105910
transform 1 0 24472 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _104_
timestamp 1626105910
transform 1 0 22724 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1626105910
transform 1 0 22080 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_231
timestamp 1626105910
transform 1 0 22356 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__D
timestamp 1626105910
transform 1 0 22172 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_220
timestamp 1626105910
transform 1 0 21344 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_208
timestamp 1626105910
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_196
timestamp 1626105910
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1626105910
transform 1 0 22080 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1626105910
transform 1 0 24748 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_237
timestamp 1626105910
transform 1 0 22908 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_249
timestamp 1626105910
transform 1 0 24012 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_225
timestamp 1626105910
transform 1 0 21804 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_213
timestamp 1626105910
transform 1 0 20700 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_201
timestamp 1626105910
transform 1 0 19596 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1626105910
transform 1 0 19504 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_241
timestamp 1626105910
transform 1 0 23276 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_241
timestamp 1626105910
transform 1 0 23276 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_229
timestamp 1626105910
transform 1 0 22172 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1626105910
transform 1 0 22080 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_220
timestamp 1626105910
transform 1 0 21344 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_208
timestamp 1626105910
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_196
timestamp 1626105910
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_220
timestamp 1626105910
transform 1 0 21344 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1626105910
transform 1 0 24748 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_237
timestamp 1626105910
transform 1 0 22908 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_249
timestamp 1626105910
transform 1 0 24012 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_225
timestamp 1626105910
transform 1 0 21804 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_213
timestamp 1626105910
transform 1 0 20700 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_201
timestamp 1626105910
transform 1 0 19596 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1626105910
transform 1 0 19504 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_208
timestamp 1626105910
transform 1 0 20240 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_241
timestamp 1626105910
transform 1 0 23276 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_229
timestamp 1626105910
transform 1 0 22172 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1626105910
transform 1 0 22080 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_220
timestamp 1626105910
transform 1 0 21344 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_208
timestamp 1626105910
transform 1 0 20240 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_196
timestamp 1626105910
transform 1 0 19136 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_192
timestamp 1626105910
transform 1 0 18768 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_192
timestamp 1626105910
transform 1 0 18768 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_187
timestamp 1626105910
transform 1 0 18308 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_184
timestamp 1626105910
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_192
timestamp 1626105910
transform 1 0 18768 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_68_194
timestamp 1626105910
transform 1 0 18952 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1626105910
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_192
timestamp 1626105910
transform 1 0 18768 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1626105910
transform 1 0 18032 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_184
timestamp 1626105910
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_192
timestamp 1626105910
transform 1 0 18768 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_184
timestamp 1626105910
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_192
timestamp 1626105910
transform 1 0 18768 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_184
timestamp 1626105910
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_192
timestamp 1626105910
transform 1 0 18768 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1626105910
transform 1 0 24748 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_237
timestamp 1626105910
transform 1 0 22908 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_249
timestamp 1626105910
transform 1 0 24012 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_225
timestamp 1626105910
transform 1 0 21804 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_213
timestamp 1626105910
transform 1 0 20700 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_201
timestamp 1626105910
transform 1 0 19596 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1626105910
transform 1 0 19504 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_184
timestamp 1626105910
transform 1 0 18032 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_182
timestamp 1626105910
transform 1 0 17848 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_194
timestamp 1626105910
transform 1 0 18952 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_170
timestamp 1626105910
transform 1 0 16744 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_158
timestamp 1626105910
transform 1 0 15640 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_146
timestamp 1626105910
transform 1 0 14536 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1626105910
transform 1 0 14260 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_137
timestamp 1626105910
transform 1 0 13708 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1626105910
transform 1 0 14352 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1626105910
transform 1 0 18032 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_192
timestamp 1626105910
transform 1 0 18768 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_184
timestamp 1626105910
transform 1 0 18032 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1626105910
transform 1 0 24748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1626105910
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1626105910
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1626105910
transform 1 0 21804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_213
timestamp 1626105910
transform 1 0 20700 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1626105910
transform 1 0 19596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1626105910
transform 1 0 19504 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_180
timestamp 1626105910
transform 1 0 17664 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_192
timestamp 1626105910
transform 1 0 18768 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1626105910
transform 1 0 16560 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_156
timestamp 1626105910
transform 1 0 15456 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1626105910
transform 1 0 14352 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1626105910
transform 1 0 14260 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_127
timestamp 1626105910
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_129
timestamp 1626105910
transform 1 0 12972 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_127
timestamp 1626105910
transform 1 0 12788 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_123
timestamp 1626105910
transform 1 0 12420 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_127
timestamp 1626105910
transform 1 0 12788 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_123
timestamp 1626105910
transform 1 0 12420 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_127
timestamp 1626105910
transform 1 0 12788 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_123
timestamp 1626105910
transform 1 0 12420 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_127
timestamp 1626105910
transform 1 0 12788 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_123
timestamp 1626105910
transform 1 0 12420 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _098_
timestamp 1626105910
transform 1 0 12880 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_73_127
timestamp 1626105910
transform 1 0 12788 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_127
timestamp 1626105910
transform 1 0 12788 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_123
timestamp 1626105910
transform 1 0 12420 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_127
timestamp 1626105910
transform 1 0 12788 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_123
timestamp 1626105910
transform 1 0 12420 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_127
timestamp 1626105910
transform 1 0 12788 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_128
timestamp 1626105910
transform 1 0 12880 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_127
timestamp 1626105910
transform 1 0 12788 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_123
timestamp 1626105910
transform 1 0 12420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_127
timestamp 1626105910
transform 1 0 12788 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_129
timestamp 1626105910
transform 1 0 12972 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B1
timestamp 1626105910
transform 1 0 13340 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_135
timestamp 1626105910
transform 1 0 13524 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _087_
timestamp 1626105910
transform 1 0 12236 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_117
timestamp 1626105910
transform 1 0 11868 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_111
timestamp 1626105910
transform 1 0 11316 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B2
timestamp 1626105910
transform 1 0 11684 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1626105910
transform 1 0 10212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_87
timestamp 1626105910
transform 1 0 9108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1626105910
transform 1 0 9016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_78
timestamp 1626105910
transform 1 0 8280 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_66
timestamp 1626105910
transform 1 0 7176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_54
timestamp 1626105910
transform 1 0 6072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_42
timestamp 1626105910
transform 1 0 4968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1626105910
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_27
timestamp 1626105910
transform 1 0 3588 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1626105910
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1626105910
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1626105910
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1626105910
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_127
timestamp 1626105910
transform 1 0 12788 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1626105910
transform 1 0 12420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_127
timestamp 1626105910
transform 1 0 12788 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_120
timestamp 1626105910
transform 1 0 12144 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_127
timestamp 1626105910
transform 1 0 12788 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_123
timestamp 1626105910
transform 1 0 12420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_127
timestamp 1626105910
transform 1 0 12788 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_123
timestamp 1626105910
transform 1 0 12420 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_127
timestamp 1626105910
transform 1 0 12788 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_123
timestamp 1626105910
transform 1 0 12420 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_127
timestamp 1626105910
transform 1 0 12788 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_123
timestamp 1626105910
transform 1 0 12420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1626105910
transform 1 0 12788 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1626105910
transform 1 0 12420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1626105910
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_123
timestamp 1626105910
transform 1 0 12420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_123
timestamp 1626105910
transform 1 0 12420 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_127
timestamp 1626105910
transform 1 0 12788 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_123
timestamp 1626105910
transform 1 0 12420 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_477
timestamp 1626105910
transform 1 0 44988 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1626105910
transform -1 0 48208 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_457
timestamp 1626105910
transform 1 0 43148 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1626105910
transform 1 0 43056 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1626105910
transform -1 0 48852 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_514
timestamp 1626105910
transform 1 0 48392 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1626105910
transform 1 0 48300 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_512
timestamp 1626105910
transform 1 0 48208 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_504
timestamp 1626105910
transform 1 0 47472 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_492
timestamp 1626105910
transform 1 0 46368 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__o311a_1  _076_
timestamp 1626105910
transform 1 0 44528 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_480
timestamp 1626105910
transform 1 0 45264 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_468
timestamp 1626105910
transform 1 0 44160 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A2
timestamp 1626105910
transform 1 0 43976 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_465
timestamp 1626105910
transform 1 0 43884 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1626105910
transform 1 0 43056 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_457
timestamp 1626105910
transform 1 0 43148 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1626105910
transform -1 0 48852 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_514
timestamp 1626105910
transform 1 0 48392 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1626105910
transform 1 0 48300 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1626105910
transform 1 0 47564 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_493
timestamp 1626105910
transform 1 0 46460 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _085_
timestamp 1626105910
transform -1 0 46828 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1626105910
transform 1 0 45724 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_497
timestamp 1626105910
transform 1 0 46828 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1626105910
transform -1 0 48852 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_510
timestamp 1626105910
transform 1 0 48024 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_498
timestamp 1626105910
transform 1 0 46920 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_486
timestamp 1626105910
transform 1 0 45816 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_482
timestamp 1626105910
transform 1 0 45448 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1626105910
transform 1 0 45724 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_470
timestamp 1626105910
transform 1 0 44344 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_465
timestamp 1626105910
transform 1 0 43884 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_486
timestamp 1626105910
transform 1 0 45816 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_465
timestamp 1626105910
transform 1 0 43884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_477
timestamp 1626105910
transform 1 0 44988 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_481
timestamp 1626105910
transform 1 0 45356 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A2
timestamp 1626105910
transform 1 0 45172 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_481
timestamp 1626105910
transform 1 0 45356 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B1
timestamp 1626105910
transform 1 0 44160 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_469
timestamp 1626105910
transform 1 0 44252 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_457
timestamp 1626105910
transform 1 0 43148 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1626105910
transform 1 0 43056 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1626105910
transform -1 0 48852 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1626105910
transform 1 0 48208 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_505
timestamp 1626105910
transform 1 0 47564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1626105910
transform -1 0 47564 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1626105910
transform -1 0 48852 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_514
timestamp 1626105910
transform 1 0 48392 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1626105910
transform 1 0 48300 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1626105910
transform 1 0 47564 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_500
timestamp 1626105910
transform 1 0 47104 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1626105910
transform -1 0 48852 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1626105910
transform -1 0 48852 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_514
timestamp 1626105910
transform 1 0 48392 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_493
timestamp 1626105910
transform 1 0 46460 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1626105910
transform -1 0 48852 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_481
timestamp 1626105910
transform 1 0 45356 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_469
timestamp 1626105910
transform 1 0 44252 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_510
timestamp 1626105910
transform 1 0 48024 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_457
timestamp 1626105910
transform 1 0 43148 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1626105910
transform 1 0 43056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_498
timestamp 1626105910
transform 1 0 46920 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_486
timestamp 1626105910
transform 1 0 45816 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1626105910
transform 1 0 48300 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_510
timestamp 1626105910
transform 1 0 48024 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_512
timestamp 1626105910
transform 1 0 48208 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_483
timestamp 1626105910
transform 1 0 45540 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1626105910
transform 1 0 45724 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_498
timestamp 1626105910
transform 1 0 46920 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1626105910
transform -1 0 48852 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__A
timestamp 1626105910
transform 1 0 44620 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_475
timestamp 1626105910
transform 1 0 44804 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_510
timestamp 1626105910
transform 1 0 48024 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_468
timestamp 1626105910
transform 1 0 44160 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A3
timestamp 1626105910
transform 1 0 43976 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_498
timestamp 1626105910
transform 1 0 46920 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_472
timestamp 1626105910
transform 1 0 44528 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_465
timestamp 1626105910
transform 1 0 43884 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_486
timestamp 1626105910
transform 1 0 45816 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1626105910
transform 1 0 45724 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_486
timestamp 1626105910
transform 1 0 45816 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_488
timestamp 1626105910
transform 1 0 46000 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1626105910
transform 1 0 45724 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A1
timestamp 1626105910
transform 1 0 45816 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_485
timestamp 1626105910
transform 1 0 45724 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_465
timestamp 1626105910
transform 1 0 43884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_469
timestamp 1626105910
transform 1 0 44252 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_465
timestamp 1626105910
transform 1 0 43884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_477
timestamp 1626105910
transform 1 0 44988 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_481
timestamp 1626105910
transform 1 0 45356 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_408
timestamp 1626105910
transform 1 0 38640 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_396
timestamp 1626105910
transform 1 0 37536 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_398
timestamp 1626105910
transform 1 0 37720 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_396
timestamp 1626105910
transform 1 0 37536 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_400
timestamp 1626105910
transform 1 0 37904 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_391
timestamp 1626105910
transform 1 0 37076 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_408
timestamp 1626105910
transform 1 0 38640 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1626105910
transform 1 0 37812 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_396
timestamp 1626105910
transform 1 0 37536 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_400
timestamp 1626105910
transform 1 0 37904 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1626105910
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_408
timestamp 1626105910
transform 1 0 38640 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_408
timestamp 1626105910
transform 1 0 38640 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_412
timestamp 1626105910
transform 1 0 39008 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_400
timestamp 1626105910
transform 1 0 37904 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_396
timestamp 1626105910
transform 1 0 37536 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1626105910
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_424
timestamp 1626105910
transform 1 0 40112 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__D
timestamp 1626105910
transform -1 0 39008 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_406
timestamp 1626105910
transform 1 0 38456 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_420
timestamp 1626105910
transform 1 0 39744 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_429
timestamp 1626105910
transform 1 0 40572 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_400
timestamp 1626105910
transform 1 0 37904 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_441
timestamp 1626105910
transform 1 0 41676 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_441
timestamp 1626105910
transform 1 0 41676 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_429
timestamp 1626105910
transform 1 0 40572 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_441
timestamp 1626105910
transform 1 0 41676 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_429
timestamp 1626105910
transform 1 0 40572 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1626105910
transform 1 0 40480 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_436
timestamp 1626105910
transform 1 0 41216 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_424
timestamp 1626105910
transform 1 0 40112 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_420
timestamp 1626105910
transform 1 0 39744 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_412
timestamp 1626105910
transform 1 0 39008 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_436
timestamp 1626105910
transform 1 0 41216 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1626105910
transform 1 0 40480 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_424
timestamp 1626105910
transform 1 0 40112 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_412
timestamp 1626105910
transform 1 0 39008 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_436
timestamp 1626105910
transform 1 0 41216 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_424
timestamp 1626105910
transform 1 0 40112 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_412
timestamp 1626105910
transform 1 0 39008 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_420
timestamp 1626105910
transform 1 0 39744 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_436
timestamp 1626105910
transform 1 0 41216 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_424
timestamp 1626105910
transform 1 0 40112 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_412
timestamp 1626105910
transform 1 0 39008 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_441
timestamp 1626105910
transform 1 0 41676 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_429
timestamp 1626105910
transform 1 0 40572 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1626105910
transform 1 0 40480 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_441
timestamp 1626105910
transform 1 0 41676 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_429
timestamp 1626105910
transform 1 0 40572 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1626105910
transform 1 0 40480 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1626105910
transform 1 0 40480 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_420
timestamp 1626105910
transform 1 0 39744 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1626105910
transform 1 0 37812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_391
timestamp 1626105910
transform 1 0 37076 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_394
timestamp 1626105910
transform 1 0 37352 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_436
timestamp 1626105910
transform 1 0 41216 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1626105910
transform 1 0 40480 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_424
timestamp 1626105910
transform 1 0 40112 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_412
timestamp 1626105910
transform 1 0 39008 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_420
timestamp 1626105910
transform 1 0 39744 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_441
timestamp 1626105910
transform 1 0 41676 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_429
timestamp 1626105910
transform 1 0 40572 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_433
timestamp 1626105910
transform 1 0 40940 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1626105910
transform 1 0 40480 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_445
timestamp 1626105910
transform 1 0 42044 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_421
timestamp 1626105910
transform 1 0 39836 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_423
timestamp 1626105910
transform 1 0 40020 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__B1
timestamp 1626105910
transform -1 0 39836 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_441
timestamp 1626105910
transform 1 0 41676 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_429
timestamp 1626105910
transform 1 0 40572 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1626105910
transform 1 0 40480 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_425
timestamp 1626105910
transform 1 0 40204 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_417
timestamp 1626105910
transform 1 0 39468 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A3
timestamp 1626105910
transform 1 0 39836 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_427
timestamp 1626105910
transform 1 0 40388 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _063_
timestamp 1626105910
transform -1 0 39468 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_54_417
timestamp 1626105910
transform 1 0 39468 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_414
timestamp 1626105910
transform 1 0 39192 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__CLK
timestamp 1626105910
transform 1 0 39008 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_418
timestamp 1626105910
transform 1 0 39560 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1626105910
transform 1 0 38180 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1626105910
transform 1 0 37812 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A1
timestamp 1626105910
transform 1 0 37996 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_408
timestamp 1626105910
transform 1 0 38640 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_438
timestamp 1626105910
transform 1 0 41400 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_426
timestamp 1626105910
transform 1 0 40296 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_420
timestamp 1626105910
transform 1 0 39744 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_414
timestamp 1626105910
transform 1 0 39192 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A2
timestamp 1626105910
transform -1 0 40296 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A3
timestamp 1626105910
transform 1 0 39560 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_396
timestamp 1626105910
transform 1 0 37536 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_400
timestamp 1626105910
transform 1 0 37904 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_391
timestamp 1626105910
transform 1 0 37076 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_429
timestamp 1626105910
transform 1 0 40572 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _075_
timestamp 1626105910
transform -1 0 39008 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_56_396
timestamp 1626105910
transform 1 0 37536 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_401
timestamp 1626105910
transform 1 0 37996 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A3
timestamp 1626105910
transform 1 0 37812 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_436
timestamp 1626105910
transform 1 0 41216 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_441
timestamp 1626105910
transform 1 0 41676 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_429
timestamp 1626105910
transform 1 0 40572 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1626105910
transform 1 0 40480 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_420
timestamp 1626105910
transform 1 0 39744 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_441
timestamp 1626105910
transform 1 0 41676 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_429
timestamp 1626105910
transform 1 0 40572 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1626105910
transform 1 0 40480 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_424
timestamp 1626105910
transform 1 0 40112 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_418
timestamp 1626105910
transform 1 0 39560 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_412
timestamp 1626105910
transform 1 0 39008 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B1
timestamp 1626105910
transform 1 0 39928 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A2
timestamp 1626105910
transform 1 0 39376 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1626105910
transform 1 0 38180 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__D
timestamp 1626105910
transform -1 0 38824 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_407
timestamp 1626105910
transform 1 0 38548 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1626105910
transform 1 0 37812 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A1
timestamp 1626105910
transform 1 0 37996 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_400
timestamp 1626105910
transform 1 0 37904 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_400
timestamp 1626105910
transform 1 0 37904 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1626105910
transform 1 0 37812 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_391
timestamp 1626105910
transform 1 0 37076 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_391
timestamp 1626105910
transform 1 0 37076 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_424
timestamp 1626105910
transform 1 0 40112 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_406
timestamp 1626105910
transform 1 0 38456 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_408
timestamp 1626105910
transform 1 0 38640 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_431
timestamp 1626105910
transform 1 0 40756 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _115_
timestamp 1626105910
transform -1 0 40756 0 1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_55_410
timestamp 1626105910
transform 1 0 38824 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_408
timestamp 1626105910
transform 1 0 38640 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_396
timestamp 1626105910
transform 1 0 37536 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_400
timestamp 1626105910
transform 1 0 37904 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1626105910
transform 1 0 37812 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_391
timestamp 1626105910
transform 1 0 37076 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A2
timestamp 1626105910
transform 1 0 38456 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A1
timestamp 1626105910
transform 1 0 38272 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1626105910
transform 1 0 37812 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_400
timestamp 1626105910
transform 1 0 37904 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_396
timestamp 1626105910
transform 1 0 37536 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_391
timestamp 1626105910
transform 1 0 37076 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_412
timestamp 1626105910
transform 1 0 39008 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_405
timestamp 1626105910
transform 1 0 38364 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__B1
timestamp 1626105910
transform -1 0 38364 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_402
timestamp 1626105910
transform 1 0 38088 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_396
timestamp 1626105910
transform 1 0 37536 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_441
timestamp 1626105910
transform 1 0 41676 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_2  _069_
timestamp 1626105910
transform -1 0 39192 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1626105910
transform -1 0 48852 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_510
timestamp 1626105910
transform 1 0 48024 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_498
timestamp 1626105910
transform 1 0 46920 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_486
timestamp 1626105910
transform 1 0 45816 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1626105910
transform 1 0 45724 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_465
timestamp 1626105910
transform 1 0 43884 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_477
timestamp 1626105910
transform 1 0 44988 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1626105910
transform 1 0 45724 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_501
timestamp 1626105910
transform 1 0 47196 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1626105910
transform -1 0 48852 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_514
timestamp 1626105910
transform 1 0 48392 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1626105910
transform 1 0 48300 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A2
timestamp 1626105910
transform 1 0 47012 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_493
timestamp 1626105910
transform 1 0 46460 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_481
timestamp 1626105910
transform 1 0 45356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_469
timestamp 1626105910
transform 1 0 44252 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_457
timestamp 1626105910
transform 1 0 43148 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1626105910
transform 1 0 43056 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_465
timestamp 1626105910
transform 1 0 43884 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _089_
timestamp 1626105910
transform -1 0 48208 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1626105910
transform -1 0 48852 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1626105910
transform 1 0 48208 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_501
timestamp 1626105910
transform 1 0 47196 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B1
timestamp 1626105910
transform 1 0 47012 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1626105910
transform 1 0 45724 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_486
timestamp 1626105910
transform 1 0 45816 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_495
timestamp 1626105910
transform 1 0 46644 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B2
timestamp 1626105910
transform 1 0 46460 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_492
timestamp 1626105910
transform 1 0 46368 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_465
timestamp 1626105910
transform 1 0 43884 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_477
timestamp 1626105910
transform 1 0 44988 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_481
timestamp 1626105910
transform 1 0 45356 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1626105910
transform -1 0 48852 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_514
timestamp 1626105910
transform 1 0 48392 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_511
timestamp 1626105910
transform 1 0 48116 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1626105910
transform 1 0 48300 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A1
timestamp 1626105910
transform 1 0 47196 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_503
timestamp 1626105910
transform 1 0 47380 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_493
timestamp 1626105910
transform 1 0 46460 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_481
timestamp 1626105910
transform 1 0 45356 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_469
timestamp 1626105910
transform 1 0 44252 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_457
timestamp 1626105910
transform 1 0 43148 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1626105910
transform 1 0 43056 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_455
timestamp 1626105910
transform 1 0 42964 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_469
timestamp 1626105910
transform 1 0 44252 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1626105910
transform -1 0 48852 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1626105910
transform -1 0 48852 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_514
timestamp 1626105910
transform 1 0 48392 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1626105910
transform 1 0 48300 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_510
timestamp 1626105910
transform 1 0 48024 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1626105910
transform 1 0 47564 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_498
timestamp 1626105910
transform 1 0 46920 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_486
timestamp 1626105910
transform 1 0 45816 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_493
timestamp 1626105910
transform 1 0 46460 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1626105910
transform 1 0 45724 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_465
timestamp 1626105910
transform 1 0 43884 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_481
timestamp 1626105910
transform 1 0 45356 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_469
timestamp 1626105910
transform 1 0 44252 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_477
timestamp 1626105910
transform 1 0 44988 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_477
timestamp 1626105910
transform 1 0 44988 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_457
timestamp 1626105910
transform 1 0 43148 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1626105910
transform 1 0 43056 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1626105910
transform 1 0 43056 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1626105910
transform 1 0 47656 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1626105910
transform -1 0 48852 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_514
timestamp 1626105910
transform 1 0 48392 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1626105910
transform -1 0 48852 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_510
timestamp 1626105910
transform 1 0 48024 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_498
timestamp 1626105910
transform 1 0 46920 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_486
timestamp 1626105910
transform 1 0 45816 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1626105910
transform 1 0 45724 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_465
timestamp 1626105910
transform 1 0 43884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_477
timestamp 1626105910
transform 1 0 44988 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1626105910
transform 1 0 48300 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_509
timestamp 1626105910
transform 1 0 47932 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_502
timestamp 1626105910
transform 1 0 47288 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1626105910
transform -1 0 47288 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_499
timestamp 1626105910
transform 1 0 47012 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_493
timestamp 1626105910
transform 1 0 46460 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_481
timestamp 1626105910
transform 1 0 45356 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_469
timestamp 1626105910
transform 1 0 44252 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_457
timestamp 1626105910
transform 1 0 43148 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1626105910
transform 1 0 43056 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_457
timestamp 1626105910
transform 1 0 43148 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1626105910
transform -1 0 48852 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1626105910
transform -1 0 48852 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_514
timestamp 1626105910
transform 1 0 48392 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1626105910
transform 1 0 48300 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_510
timestamp 1626105910
transform 1 0 48024 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1626105910
transform 1 0 47564 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_498
timestamp 1626105910
transform 1 0 46920 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_486
timestamp 1626105910
transform 1 0 45816 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_493
timestamp 1626105910
transform 1 0 46460 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_453
timestamp 1626105910
transform 1 0 42780 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_450
timestamp 1626105910
transform 1 0 42504 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_453
timestamp 1626105910
transform 1 0 42780 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_443
timestamp 1626105910
transform 1 0 41860 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_453
timestamp 1626105910
transform 1 0 42780 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_453
timestamp 1626105910
transform 1 0 42780 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_400
timestamp 1626105910
transform 1 0 37904 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1626105910
transform 1 0 37812 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_395
timestamp 1626105910
transform 1 0 37444 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_453
timestamp 1626105910
transform 1 0 42780 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_510
timestamp 1626105910
transform 1 0 48024 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1626105910
transform -1 0 48852 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_514
timestamp 1626105910
transform 1 0 48392 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1626105910
transform 1 0 48300 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_498
timestamp 1626105910
transform 1 0 46920 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_486
timestamp 1626105910
transform 1 0 45816 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _051_
timestamp 1626105910
transform -1 0 45816 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_473
timestamp 1626105910
transform 1 0 44620 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_469
timestamp 1626105910
transform 1 0 44252 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__B
timestamp 1626105910
transform -1 0 44620 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_457
timestamp 1626105910
transform 1 0 43148 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_453
timestamp 1626105910
transform 1 0 42780 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1626105910
transform 1 0 43056 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_448
timestamp 1626105910
transform 1 0 42320 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_436
timestamp 1626105910
transform 1 0 41216 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_424
timestamp 1626105910
transform 1 0 40112 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_412
timestamp 1626105910
transform 1 0 39008 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_448
timestamp 1626105910
transform 1 0 42320 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_453
timestamp 1626105910
transform 1 0 42780 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_448
timestamp 1626105910
transform 1 0 42320 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_453
timestamp 1626105910
transform 1 0 42780 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_448
timestamp 1626105910
transform 1 0 42320 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_453
timestamp 1626105910
transform 1 0 42780 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_448
timestamp 1626105910
transform 1 0 42320 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_453
timestamp 1626105910
transform 1 0 42780 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_448
timestamp 1626105910
transform 1 0 42320 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_453
timestamp 1626105910
transform 1 0 42780 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_448
timestamp 1626105910
transform 1 0 42320 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_383
timestamp 1626105910
transform 1 0 36340 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1626105910
transform 1 0 35236 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__CLK
timestamp 1626105910
transform 1 0 36156 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_380
timestamp 1626105910
transform 1 0 36064 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_370
timestamp 1626105910
transform 1 0 35144 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_372
timestamp 1626105910
transform 1 0 35328 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_362
timestamp 1626105910
transform 1 0 34408 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_350
timestamp 1626105910
transform 1 0 33304 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_338
timestamp 1626105910
transform 1 0 32200 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_326
timestamp 1626105910
transform 1 0 31096 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1626105910
transform 1 0 35236 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_335
timestamp 1626105910
transform 1 0 31924 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1626105910
transform 1 0 33396 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__CLK
timestamp 1626105910
transform 1 0 32108 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1626105910
transform 1 0 34316 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1626105910
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_327
timestamp 1626105910
transform 1 0 31188 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1626105910
transform 1 0 34868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_375
timestamp 1626105910
transform 1 0 35604 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_363
timestamp 1626105910
transform 1 0 34500 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_351
timestamp 1626105910
transform 1 0 33396 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1626105910
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_345
timestamp 1626105910
transform 1 0 32844 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__C1
timestamp 1626105910
transform -1 0 33396 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__B1
timestamp 1626105910
transform 1 0 32660 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_1  _061_
timestamp 1626105910
transform 1 0 31464 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_340
timestamp 1626105910
transform 1 0 32384 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_338
timestamp 1626105910
transform 1 0 32200 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_326
timestamp 1626105910
transform 1 0 31096 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_328
timestamp 1626105910
transform 1 0 31280 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_334
timestamp 1626105910
transform 1 0 31832 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_370
timestamp 1626105910
transform 1 0 35144 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1626105910
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_364
timestamp 1626105910
transform 1 0 34592 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_364
timestamp 1626105910
transform 1 0 34592 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1626105910
transform 1 0 32292 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1626105910
transform 1 0 34960 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_363
timestamp 1626105910
transform 1 0 34500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_345
timestamp 1626105910
transform 1 0 32844 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1626105910
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1626105910
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_357
timestamp 1626105910
transform 1 0 33948 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1626105910
transform 1 0 33396 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_363
timestamp 1626105910
transform 1 0 34500 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_351
timestamp 1626105910
transform 1 0 33396 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_372
timestamp 1626105910
transform 1 0 35328 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_372
timestamp 1626105910
transform 1 0 35328 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_372
timestamp 1626105910
transform 1 0 35328 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_339
timestamp 1626105910
transform 1 0 32292 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__RESET_B
timestamp 1626105910
transform -1 0 32844 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_370
timestamp 1626105910
transform 1 0 35144 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_341
timestamp 1626105910
transform 1 0 32476 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1626105910
transform 1 0 32292 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_335
timestamp 1626105910
transform 1 0 31924 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_327
timestamp 1626105910
transform 1 0 31188 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_327
timestamp 1626105910
transform 1 0 31188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_334
timestamp 1626105910
transform 1 0 31832 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1626105910
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_363
timestamp 1626105910
transform 1 0 34500 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1626105910
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A2
timestamp 1626105910
transform 1 0 31096 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_355
timestamp 1626105910
transform 1 0 33764 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_355
timestamp 1626105910
transform 1 0 33764 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_343
timestamp 1626105910
transform 1 0 32660 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_352
timestamp 1626105910
transform 1 0 33488 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_367
timestamp 1626105910
transform 1 0 34868 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1626105910
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B1
timestamp 1626105910
transform 1 0 34684 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_343
timestamp 1626105910
transform 1 0 32660 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_372
timestamp 1626105910
transform 1 0 35328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_306
timestamp 1626105910
transform 1 0 29256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_323
timestamp 1626105910
transform 1 0 30820 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1626105910
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_315
timestamp 1626105910
transform 1 0 30084 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_306
timestamp 1626105910
transform 1 0 29256 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_294
timestamp 1626105910
transform 1 0 28152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_282
timestamp 1626105910
transform 1 0 27048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_322
timestamp 1626105910
transform 1 0 30728 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_284
timestamp 1626105910
transform 1 0 27232 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_310
timestamp 1626105910
transform 1 0 29624 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_298
timestamp 1626105910
transform 1 0 28520 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1626105910
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1626105910
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1626105910
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_294
timestamp 1626105910
transform 1 0 28152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1626105910
transform 1 0 27048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_279
timestamp 1626105910
transform 1 0 26772 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_310
timestamp 1626105910
transform 1 0 29624 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_298
timestamp 1626105910
transform 1 0 28520 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1626105910
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_306
timestamp 1626105910
transform 1 0 29256 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1626105910
transform 1 0 28152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_282
timestamp 1626105910
transform 1 0 27048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1626105910
transform 1 0 27416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A2
timestamp 1626105910
transform 1 0 27140 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1626105910
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_306
timestamp 1626105910
transform 1 0 29256 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_277
timestamp 1626105910
transform 1 0 26588 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A1
timestamp 1626105910
transform 1 0 26588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_276
timestamp 1626105910
transform 1 0 26496 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1626105910
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_310
timestamp 1626105910
transform 1 0 29624 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1626105910
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_310
timestamp 1626105910
transform 1 0 29624 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_298
timestamp 1626105910
transform 1 0 28520 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_286
timestamp 1626105910
transform 1 0 27416 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_298
timestamp 1626105910
transform 1 0 28520 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_286
timestamp 1626105910
transform 1 0 27416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_297
timestamp 1626105910
transform 1 0 28428 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1626105910
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_306
timestamp 1626105910
transform 1 0 29256 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1626105910
transform 1 0 28152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1626105910
transform 1 0 27048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1626105910
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1626105910
transform 1 0 25944 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_273
timestamp 1626105910
transform 1 0 26220 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _078_
timestamp 1626105910
transform 1 0 25576 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_50_309
timestamp 1626105910
transform 1 0 29532 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1626105910
transform 1 0 25944 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1626105910
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_262
timestamp 1626105910
transform 1 0 25208 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A3
timestamp 1626105910
transform 1 0 25024 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_264
timestamp 1626105910
transform 1 0 25392 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B1
timestamp 1626105910
transform 1 0 25208 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_261
timestamp 1626105910
transform 1 0 25116 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1626105910
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_270
timestamp 1626105910
transform 1 0 25944 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_265
timestamp 1626105910
transform 1 0 25484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_265
timestamp 1626105910
transform 1 0 25484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__D
timestamp 1626105910
transform -1 0 29624 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_313
timestamp 1626105910
transform 1 0 29900 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1626105910
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_285
timestamp 1626105910
transform 1 0 27324 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1626105910
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_315
timestamp 1626105910
transform 1 0 30084 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_270
timestamp 1626105910
transform 1 0 25944 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1626105910
transform 1 0 25484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_306
timestamp 1626105910
transform 1 0 29256 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1626105910
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_310
timestamp 1626105910
transform 1 0 29624 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_306
timestamp 1626105910
transform 1 0 29256 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_294
timestamp 1626105910
transform 1 0 28152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1626105910
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_310
timestamp 1626105910
transform 1 0 29624 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_298
timestamp 1626105910
transform 1 0 28520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1626105910
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1626105910
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_277
timestamp 1626105910
transform 1 0 26588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_315
timestamp 1626105910
transform 1 0 30084 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1626105910
transform -1 0 30728 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_306
timestamp 1626105910
transform 1 0 29256 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1626105910
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1626105910
transform 1 0 27048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_298
timestamp 1626105910
transform 1 0 28520 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_286
timestamp 1626105910
transform 1 0 27416 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_282
timestamp 1626105910
transform 1 0 27048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1626105910
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1626105910
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_270
timestamp 1626105910
transform 1 0 25944 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_310
timestamp 1626105910
transform 1 0 29624 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_298
timestamp 1626105910
transform 1 0 28520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1626105910
transform 1 0 29992 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_310
timestamp 1626105910
transform 1 0 29624 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_306
timestamp 1626105910
transform 1 0 29256 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1626105910
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_298
timestamp 1626105910
transform 1 0 28520 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1626105910
transform 1 0 27416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_282
timestamp 1626105910
transform 1 0 27048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1626105910
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_277
timestamp 1626105910
transform 1 0 26588 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1626105910
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1626105910
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_277
timestamp 1626105910
transform 1 0 26588 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_294
timestamp 1626105910
transform 1 0 28152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_282
timestamp 1626105910
transform 1 0 27048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1626105910
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_265
timestamp 1626105910
transform 1 0 25484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1626105910
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_306
timestamp 1626105910
transform 1 0 29256 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1626105910
transform 1 0 28152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_282
timestamp 1626105910
transform 1 0 27048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_270
timestamp 1626105910
transform 1 0 25944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_265
timestamp 1626105910
transform 1 0 25484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1626105910
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_265
timestamp 1626105910
transform 1 0 25484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1626105910
transform 1 0 25944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_265
timestamp 1626105910
transform 1 0 25484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_310
timestamp 1626105910
transform 1 0 29624 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_298
timestamp 1626105910
transform 1 0 28520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_286
timestamp 1626105910
transform 1 0 27416 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1626105910
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_277
timestamp 1626105910
transform 1 0 26588 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_334
timestamp 1626105910
transform 1 0 31832 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1626105910
transform 1 0 35328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1626105910
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_355
timestamp 1626105910
transform 1 0 33764 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_343
timestamp 1626105910
transform 1 0 32660 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1626105910
transform 1 0 32568 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_334
timestamp 1626105910
transform 1 0 31832 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1626105910
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1626105910
transform 1 0 35328 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1626105910
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1626105910
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_351
timestamp 1626105910
transform 1 0 33396 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_355
timestamp 1626105910
transform 1 0 33764 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_363
timestamp 1626105910
transform 1 0 34500 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_339
timestamp 1626105910
transform 1 0 32292 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_343
timestamp 1626105910
transform 1 0 32660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1626105910
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_327
timestamp 1626105910
transform 1 0 31188 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_334
timestamp 1626105910
transform 1 0 31832 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_365
timestamp 1626105910
transform 1 0 34684 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _105_
timestamp 1626105910
transform -1 0 34684 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_58_372
timestamp 1626105910
transform 1 0 35328 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1626105910
transform 1 0 35236 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_351
timestamp 1626105910
transform 1 0 33396 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_363
timestamp 1626105910
transform 1 0 34500 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_339
timestamp 1626105910
transform 1 0 32292 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1626105910
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_342
timestamp 1626105910
transform 1 0 32568 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1626105910
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_355
timestamp 1626105910
transform 1 0 33764 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1626105910
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1626105910
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_334
timestamp 1626105910
transform 1 0 31832 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__CLK
timestamp 1626105910
transform 1 0 32384 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_372
timestamp 1626105910
transform 1 0 35328 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1626105910
transform 1 0 35236 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_370
timestamp 1626105910
transform 1 0 35144 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_358
timestamp 1626105910
transform 1 0 34040 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_346
timestamp 1626105910
transform 1 0 32936 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_334
timestamp 1626105910
transform 1 0 31832 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_339
timestamp 1626105910
transform 1 0 32292 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1626105910
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1626105910
transform 1 0 33764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1626105910
transform 1 0 32660 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1626105910
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_334
timestamp 1626105910
transform 1 0 31832 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_327
timestamp 1626105910
transform 1 0 31188 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_372
timestamp 1626105910
transform 1 0 35328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1626105910
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1626105910
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_351
timestamp 1626105910
transform 1 0 33396 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1626105910
transform 1 0 33764 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_363
timestamp 1626105910
transform 1 0 34500 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_339
timestamp 1626105910
transform 1 0 32292 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1626105910
transform 1 0 32660 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1626105910
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_327
timestamp 1626105910
transform 1 0 31188 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A3
timestamp 1626105910
transform 1 0 30912 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A1
timestamp 1626105910
transform -1 0 31096 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_322
timestamp 1626105910
transform 1 0 30728 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_315
timestamp 1626105910
transform 1 0 30084 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_322
timestamp 1626105910
transform 1 0 30728 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1626105910
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1626105910
transform 1 0 30728 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_322
timestamp 1626105910
transform 1 0 30728 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1626105910
transform 1 0 30728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1626105910
transform 1 0 30084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_322
timestamp 1626105910
transform 1 0 30728 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_323
timestamp 1626105910
transform 1 0 30820 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_322
timestamp 1626105910
transform 1 0 30728 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_315
timestamp 1626105910
transform 1 0 30084 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _102_
timestamp 1626105910
transform 1 0 29992 0 1 26656
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_42_315
timestamp 1626105910
transform 1 0 30084 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1626105910
transform 1 0 25484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1626105910
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_377
timestamp 1626105910
transform 1 0 35788 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A2
timestamp 1626105910
transform 1 0 36156 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o311a_1  _073_
timestamp 1626105910
transform 1 0 35052 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_365
timestamp 1626105910
transform 1 0 34684 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A3
timestamp 1626105910
transform 1 0 34500 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1626105910
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_359
timestamp 1626105910
transform 1 0 34132 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_353
timestamp 1626105910
transform 1 0 33580 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__C1
timestamp 1626105910
transform -1 0 33580 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A1
timestamp 1626105910
transform -1 0 34132 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_343
timestamp 1626105910
transform 1 0 32660 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1626105910
transform 1 0 30728 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_334
timestamp 1626105910
transform 1 0 31832 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1626105910
transform 1 0 29624 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_298
timestamp 1626105910
transform 1 0 28520 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_315
timestamp 1626105910
transform 1 0 30084 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_286
timestamp 1626105910
transform 1 0 27416 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1626105910
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_277
timestamp 1626105910
transform 1 0 26588 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_322
timestamp 1626105910
transform 1 0 30728 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_372
timestamp 1626105910
transform 1 0 35328 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1626105910
transform 1 0 35236 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_327
timestamp 1626105910
transform 1 0 31188 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_351
timestamp 1626105910
transform 1 0 33396 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_363
timestamp 1626105910
transform 1 0 34500 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_339
timestamp 1626105910
transform 1 0 32292 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_363
timestamp 1626105910
transform 1 0 34500 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_339
timestamp 1626105910
transform 1 0 32292 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_327
timestamp 1626105910
transform 1 0 31188 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_372
timestamp 1626105910
transform 1 0 35328 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1626105910
transform 1 0 35236 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_351
timestamp 1626105910
transform 1 0 33396 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_363
timestamp 1626105910
transform 1 0 34500 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_339
timestamp 1626105910
transform 1 0 32292 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_327
timestamp 1626105910
transform 1 0 31188 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1626105910
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_355
timestamp 1626105910
transform 1 0 33764 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1626105910
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_355
timestamp 1626105910
transform 1 0 33764 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_343
timestamp 1626105910
transform 1 0 32660 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1626105910
transform 1 0 32568 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_334
timestamp 1626105910
transform 1 0 31832 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_327
timestamp 1626105910
transform 1 0 31188 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_355
timestamp 1626105910
transform 1 0 33764 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_343
timestamp 1626105910
transform 1 0 32660 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1626105910
transform 1 0 34868 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_377
timestamp 1626105910
transform 1 0 35788 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_355
timestamp 1626105910
transform 1 0 33764 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_365
timestamp 1626105910
transform 1 0 34684 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_372
timestamp 1626105910
transform 1 0 35328 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1626105910
transform 1 0 35236 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_353
timestamp 1626105910
transform 1 0 33580 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_359
timestamp 1626105910
transform 1 0 34132 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _057_
timestamp 1626105910
transform -1 0 33580 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_347
timestamp 1626105910
transform 1 0 33028 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1626105910
transform 1 0 32568 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_339
timestamp 1626105910
transform 1 0 32292 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_343
timestamp 1626105910
transform 1 0 32660 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A
timestamp 1626105910
transform 1 0 32844 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_341
timestamp 1626105910
transform 1 0 32476 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_329
timestamp 1626105910
transform 1 0 31372 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_327
timestamp 1626105910
transform 1 0 31188 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_343
timestamp 1626105910
transform 1 0 32660 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_339
timestamp 1626105910
transform 1 0 32292 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1626105910
transform 1 0 32568 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_372
timestamp 1626105910
transform 1 0 35328 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1626105910
transform 1 0 35236 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_351
timestamp 1626105910
transform 1 0 33396 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1626105910
transform 1 0 32568 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_334
timestamp 1626105910
transform 1 0 31832 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_367
timestamp 1626105910
transform 1 0 34868 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_343
timestamp 1626105910
transform 1 0 32660 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1626105910
transform 1 0 32568 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_334
timestamp 1626105910
transform 1 0 31832 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_303
timestamp 1626105910
transform 1 0 28980 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_310
timestamp 1626105910
transform 1 0 29624 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_298
timestamp 1626105910
transform 1 0 28520 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_286
timestamp 1626105910
transform 1 0 27416 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1626105910
transform 1 0 27324 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_277
timestamp 1626105910
transform 1 0 26588 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1626105910
transform 1 0 27324 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_277
timestamp 1626105910
transform 1 0 26588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1626105910
transform -1 0 25300 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_270
timestamp 1626105910
transform 1 0 25944 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1626105910
transform 1 0 29992 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_306
timestamp 1626105910
transform 1 0 29256 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_294
timestamp 1626105910
transform 1 0 28152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_282
timestamp 1626105910
transform 1 0 27048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_265
timestamp 1626105910
transform 1 0 25484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_270
timestamp 1626105910
transform 1 0 25944 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_265
timestamp 1626105910
transform 1 0 25484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_265
timestamp 1626105910
transform 1 0 25484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1626105910
transform 1 0 27324 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_277
timestamp 1626105910
transform 1 0 26588 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_298
timestamp 1626105910
transform 1 0 28520 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1626105910
transform 1 0 29992 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_306
timestamp 1626105910
transform 1 0 29256 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1626105910
transform 1 0 29992 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_313
timestamp 1626105910
transform 1 0 29900 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1626105910
transform 1 0 29164 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_309
timestamp 1626105910
transform 1 0 29532 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_303
timestamp 1626105910
transform 1 0 28980 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1626105910
transform -1 0 29164 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__C
timestamp 1626105910
transform -1 0 29532 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__D
timestamp 1626105910
transform 1 0 28796 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_294
timestamp 1626105910
transform 1 0 28152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_282
timestamp 1626105910
transform 1 0 27048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_286
timestamp 1626105910
transform 1 0 27416 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_263
timestamp 1626105910
transform 1 0 25300 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_302
timestamp 1626105910
transform 1 0 28888 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _094_
timestamp 1626105910
transform -1 0 28428 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_67_286
timestamp 1626105910
transform 1 0 27416 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_298
timestamp 1626105910
transform 1 0 28520 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_297
timestamp 1626105910
transform 1 0 28428 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_283
timestamp 1626105910
transform 1 0 27140 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1626105910
transform 1 0 27324 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_282
timestamp 1626105910
transform 1 0 27048 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_275
timestamp 1626105910
transform 1 0 26404 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__B
timestamp 1626105910
transform 1 0 28796 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_286
timestamp 1626105910
transform 1 0 27416 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_298
timestamp 1626105910
transform 1 0 28520 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1626105910
transform 1 0 27324 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_270
timestamp 1626105910
transform 1 0 25944 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_310
timestamp 1626105910
transform 1 0 29624 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_270
timestamp 1626105910
transform 1 0 25944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_310
timestamp 1626105910
transform 1 0 29624 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_298
timestamp 1626105910
transform 1 0 28520 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_286
timestamp 1626105910
transform 1 0 27416 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1626105910
transform 1 0 29992 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_306
timestamp 1626105910
transform 1 0 29256 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_294
timestamp 1626105910
transform 1 0 28152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_282
timestamp 1626105910
transform 1 0 27048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_265
timestamp 1626105910
transform 1 0 25484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_277
timestamp 1626105910
transform 1 0 26588 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_298
timestamp 1626105910
transform 1 0 28520 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_286
timestamp 1626105910
transform 1 0 27416 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_272
timestamp 1626105910
transform 1 0 26128 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_260
timestamp 1626105910
transform 1 0 25024 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_270
timestamp 1626105910
transform 1 0 25944 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_265
timestamp 1626105910
transform 1 0 25484 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1626105910
transform 1 0 27324 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_284
timestamp 1626105910
transform 1 0 27232 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_277
timestamp 1626105910
transform 1 0 26588 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_294
timestamp 1626105910
transform 1 0 28152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_282
timestamp 1626105910
transform 1 0 27048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_310
timestamp 1626105910
transform 1 0 29624 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1626105910
transform 1 0 29992 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_306
timestamp 1626105910
transform 1 0 29256 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_294
timestamp 1626105910
transform 1 0 28152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_282
timestamp 1626105910
transform 1 0 27048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1626105910
transform 1 0 29992 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_306
timestamp 1626105910
transform 1 0 29256 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_294
timestamp 1626105910
transform 1 0 28152 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_282
timestamp 1626105910
transform 1 0 27048 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_277
timestamp 1626105910
transform 1 0 26588 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_298
timestamp 1626105910
transform 1 0 28520 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_286
timestamp 1626105910
transform 1 0 27416 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1626105910
transform 1 0 27324 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1626105910
transform 1 0 29992 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_306
timestamp 1626105910
transform 1 0 29256 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_310
timestamp 1626105910
transform 1 0 29624 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1626105910
transform 1 0 30452 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_298
timestamp 1626105910
transform 1 0 28520 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_303
timestamp 1626105910
transform 1 0 28980 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_310
timestamp 1626105910
transform 1 0 29624 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_298
timestamp 1626105910
transform 1 0 28520 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_286
timestamp 1626105910
transform 1 0 27416 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1626105910
transform 1 0 29992 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_315
timestamp 1626105910
transform 1 0 30084 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_306
timestamp 1626105910
transform 1 0 29256 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_291
timestamp 1626105910
transform 1 0 27876 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_274
timestamp 1626105910
transform 1 0 26312 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_286
timestamp 1626105910
transform 1 0 27416 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_294
timestamp 1626105910
transform 1 0 28152 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_282
timestamp 1626105910
transform 1 0 27048 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1626105910
transform 1 0 27784 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1626105910
transform 1 0 27324 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_286
timestamp 1626105910
transform 1 0 27416 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_277
timestamp 1626105910
transform 1 0 26588 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_265
timestamp 1626105910
transform 1 0 25484 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_270
timestamp 1626105910
transform 1 0 25944 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_262
timestamp 1626105910
transform 1 0 25208 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1626105910
transform 1 0 25116 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_270
timestamp 1626105910
transform 1 0 25944 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_265
timestamp 1626105910
transform 1 0 25484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_270
timestamp 1626105910
transform 1 0 25944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_265
timestamp 1626105910
transform 1 0 25484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1626105910
transform 1 0 27324 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_277
timestamp 1626105910
transform 1 0 26588 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_310
timestamp 1626105910
transform 1 0 29624 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_298
timestamp 1626105910
transform 1 0 28520 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_286
timestamp 1626105910
transform 1 0 27416 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1626105910
transform 1 0 27324 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_310
timestamp 1626105910
transform 1 0 29624 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1626105910
transform 1 0 32568 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_334
timestamp 1626105910
transform 1 0 31832 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_343
timestamp 1626105910
transform 1 0 32660 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_372
timestamp 1626105910
transform 1 0 35328 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_361
timestamp 1626105910
transform 1 0 34316 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_367
timestamp 1626105910
transform 1 0 34868 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_372
timestamp 1626105910
transform 1 0 35328 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1626105910
transform 1 0 35788 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1626105910
transform 1 0 35236 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_373
timestamp 1626105910
transform 1 0 35420 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_363
timestamp 1626105910
transform 1 0 34500 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1626105910
transform 1 0 33212 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_355
timestamp 1626105910
transform 1 0 33764 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_343
timestamp 1626105910
transform 1 0 32660 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_351
timestamp 1626105910
transform 1 0 33396 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_339
timestamp 1626105910
transform 1 0 32292 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1626105910
transform 1 0 33120 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1626105910
transform 1 0 32568 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_344
timestamp 1626105910
transform 1 0 32752 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_332
timestamp 1626105910
transform 1 0 31648 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1626105910
transform 1 0 35236 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_351
timestamp 1626105910
transform 1 0 33396 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_327
timestamp 1626105910
transform 1 0 31188 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_334
timestamp 1626105910
transform 1 0 31832 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_363
timestamp 1626105910
transform 1 0 34500 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_367
timestamp 1626105910
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_355
timestamp 1626105910
transform 1 0 33764 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_343
timestamp 1626105910
transform 1 0 32660 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1626105910
transform 1 0 32568 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_334
timestamp 1626105910
transform 1 0 31832 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_339
timestamp 1626105910
transform 1 0 32292 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_327
timestamp 1626105910
transform 1 0 31188 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_372
timestamp 1626105910
transform 1 0 35328 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1626105910
transform 1 0 35236 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_351
timestamp 1626105910
transform 1 0 33396 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_363
timestamp 1626105910
transform 1 0 34500 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_339
timestamp 1626105910
transform 1 0 32292 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_327
timestamp 1626105910
transform 1 0 31188 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_355
timestamp 1626105910
transform 1 0 33764 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_367
timestamp 1626105910
transform 1 0 34868 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_355
timestamp 1626105910
transform 1 0 33764 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_343
timestamp 1626105910
transform 1 0 32660 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1626105910
transform 1 0 32568 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_334
timestamp 1626105910
transform 1 0 31832 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_334
timestamp 1626105910
transform 1 0 31832 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1626105910
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_372
timestamp 1626105910
transform 1 0 35328 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1626105910
transform 1 0 35236 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_351
timestamp 1626105910
transform 1 0 33396 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_363
timestamp 1626105910
transform 1 0 34500 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_339
timestamp 1626105910
transform 1 0 32292 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_327
timestamp 1626105910
transform 1 0 31188 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1626105910
transform 1 0 32568 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1626105910
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_355
timestamp 1626105910
transform 1 0 33764 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_343
timestamp 1626105910
transform 1 0 32660 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_322
timestamp 1626105910
transform 1 0 30728 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_315
timestamp 1626105910
transform 1 0 30084 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1626105910
transform 1 0 30268 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_315
timestamp 1626105910
transform 1 0 30084 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_320
timestamp 1626105910
transform 1 0 30544 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_322
timestamp 1626105910
transform 1 0 30728 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_315
timestamp 1626105910
transform 1 0 30084 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_322
timestamp 1626105910
transform 1 0 30728 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_315
timestamp 1626105910
transform 1 0 30084 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_315
timestamp 1626105910
transform 1 0 30084 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_322
timestamp 1626105910
transform 1 0 30728 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_270
timestamp 1626105910
transform 1 0 25944 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_315
timestamp 1626105910
transform 1 0 30084 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_322
timestamp 1626105910
transform 1 0 30728 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_315
timestamp 1626105910
transform 1 0 30084 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_315
timestamp 1626105910
transform 1 0 30084 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_372
timestamp 1626105910
transform 1 0 35328 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1626105910
transform 1 0 35236 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_351
timestamp 1626105910
transform 1 0 33396 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_363
timestamp 1626105910
transform 1 0 34500 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_339
timestamp 1626105910
transform 1 0 32292 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_327
timestamp 1626105910
transform 1 0 31188 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_322
timestamp 1626105910
transform 1 0 30728 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_315
timestamp 1626105910
transform 1 0 30084 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1626105910
transform 1 0 29992 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_306
timestamp 1626105910
transform 1 0 29256 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_294
timestamp 1626105910
transform 1 0 28152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_282
timestamp 1626105910
transform 1 0 27048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_322
timestamp 1626105910
transform 1 0 30728 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_315
timestamp 1626105910
transform 1 0 30084 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_322
timestamp 1626105910
transform 1 0 30728 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_486
timestamp 1626105910
transform 1 0 45816 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1626105910
transform 1 0 45724 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_481
timestamp 1626105910
transform 1 0 45356 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_469
timestamp 1626105910
transform 1 0 44252 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_465
timestamp 1626105910
transform 1 0 43884 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_477
timestamp 1626105910
transform 1 0 44988 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_457
timestamp 1626105910
transform 1 0 43148 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_486
timestamp 1626105910
transform 1 0 45816 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1626105910
transform 1 0 43056 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1626105910
transform 1 0 45724 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_465
timestamp 1626105910
transform 1 0 43884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_477
timestamp 1626105910
transform 1 0 44988 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_493
timestamp 1626105910
transform 1 0 46460 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_481
timestamp 1626105910
transform 1 0 45356 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_469
timestamp 1626105910
transform 1 0 44252 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1626105910
transform -1 0 48852 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_514
timestamp 1626105910
transform 1 0 48392 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1626105910
transform 1 0 48300 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1626105910
transform 1 0 47564 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_493
timestamp 1626105910
transform 1 0 46460 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_481
timestamp 1626105910
transform 1 0 45356 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_469
timestamp 1626105910
transform 1 0 44252 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_457
timestamp 1626105910
transform 1 0 43148 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1626105910
transform 1 0 43056 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_457
timestamp 1626105910
transform 1 0 43148 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1626105910
transform 1 0 43056 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1626105910
transform -1 0 48852 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_514
timestamp 1626105910
transform 1 0 48392 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1626105910
transform -1 0 48852 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_510
timestamp 1626105910
transform 1 0 48024 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_498
timestamp 1626105910
transform 1 0 46920 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_486
timestamp 1626105910
transform 1 0 45816 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1626105910
transform 1 0 45724 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_465
timestamp 1626105910
transform 1 0 43884 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_477
timestamp 1626105910
transform 1 0 44988 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1626105910
transform 1 0 48300 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1626105910
transform 1 0 47564 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_493
timestamp 1626105910
transform 1 0 46460 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_481
timestamp 1626105910
transform 1 0 45356 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_469
timestamp 1626105910
transform 1 0 44252 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1626105910
transform -1 0 48852 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_514
timestamp 1626105910
transform 1 0 48392 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1626105910
transform 1 0 48300 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1626105910
transform 1 0 47564 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_493
timestamp 1626105910
transform 1 0 46460 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_481
timestamp 1626105910
transform 1 0 45356 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_469
timestamp 1626105910
transform 1 0 44252 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_457
timestamp 1626105910
transform 1 0 43148 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1626105910
transform 1 0 43056 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_457
timestamp 1626105910
transform 1 0 43148 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1626105910
transform 1 0 43056 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1626105910
transform -1 0 48852 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_514
timestamp 1626105910
transform 1 0 48392 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1626105910
transform -1 0 48852 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_510
timestamp 1626105910
transform 1 0 48024 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_498
timestamp 1626105910
transform 1 0 46920 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_486
timestamp 1626105910
transform 1 0 45816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1626105910
transform 1 0 45724 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_465
timestamp 1626105910
transform 1 0 43884 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_477
timestamp 1626105910
transform 1 0 44988 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1626105910
transform 1 0 48300 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1626105910
transform 1 0 47564 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1626105910
transform -1 0 48852 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_510
timestamp 1626105910
transform 1 0 48024 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_498
timestamp 1626105910
transform 1 0 46920 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1626105910
transform -1 0 48852 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1626105910
transform -1 0 48852 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_514
timestamp 1626105910
transform 1 0 48392 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1626105910
transform 1 0 48300 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_510
timestamp 1626105910
transform 1 0 48024 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1626105910
transform 1 0 47564 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_493
timestamp 1626105910
transform 1 0 46460 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_498
timestamp 1626105910
transform 1 0 46920 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_391
timestamp 1626105910
transform 1 0 37076 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_408
timestamp 1626105910
transform 1 0 38640 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_408
timestamp 1626105910
transform 1 0 38640 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_396
timestamp 1626105910
transform 1 0 37536 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_396
timestamp 1626105910
transform 1 0 37536 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_408
timestamp 1626105910
transform 1 0 38640 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_436
timestamp 1626105910
transform 1 0 41216 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_424
timestamp 1626105910
transform 1 0 40112 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_412
timestamp 1626105910
transform 1 0 39008 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1626105910
transform 1 0 37812 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_441
timestamp 1626105910
transform 1 0 41676 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_429
timestamp 1626105910
transform 1 0 40572 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1626105910
transform 1 0 40480 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_420
timestamp 1626105910
transform 1 0 39744 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_400
timestamp 1626105910
transform 1 0 37904 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_436
timestamp 1626105910
transform 1 0 41216 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_424
timestamp 1626105910
transform 1 0 40112 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_412
timestamp 1626105910
transform 1 0 39008 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_397
timestamp 1626105910
transform 1 0 37628 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_441
timestamp 1626105910
transform 1 0 41676 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_429
timestamp 1626105910
transform 1 0 40572 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1626105910
transform 1 0 40480 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_420
timestamp 1626105910
transform 1 0 39744 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_400
timestamp 1626105910
transform 1 0 37904 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_400
timestamp 1626105910
transform 1 0 37904 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_436
timestamp 1626105910
transform 1 0 41216 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_441
timestamp 1626105910
transform 1 0 41676 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_429
timestamp 1626105910
transform 1 0 40572 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1626105910
transform 1 0 40480 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_424
timestamp 1626105910
transform 1 0 40112 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_412
timestamp 1626105910
transform 1 0 39008 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_420
timestamp 1626105910
transform 1 0 39744 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_391
timestamp 1626105910
transform 1 0 37076 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_436
timestamp 1626105910
transform 1 0 41216 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_424
timestamp 1626105910
transform 1 0 40112 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_412
timestamp 1626105910
transform 1 0 39008 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_396
timestamp 1626105910
transform 1 0 37536 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_441
timestamp 1626105910
transform 1 0 41676 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_429
timestamp 1626105910
transform 1 0 40572 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1626105910
transform 1 0 40480 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_420
timestamp 1626105910
transform 1 0 39744 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1626105910
transform 1 0 37812 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_436
timestamp 1626105910
transform 1 0 41216 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_424
timestamp 1626105910
transform 1 0 40112 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_412
timestamp 1626105910
transform 1 0 39008 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_391
timestamp 1626105910
transform 1 0 37076 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_408
timestamp 1626105910
transform 1 0 38640 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_400
timestamp 1626105910
transform 1 0 37904 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1626105910
transform 1 0 37812 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_396
timestamp 1626105910
transform 1 0 37536 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_391
timestamp 1626105910
transform 1 0 37076 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1626105910
transform 1 0 37812 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_400
timestamp 1626105910
transform 1 0 37904 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1626105910
transform 1 0 37812 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_400
timestamp 1626105910
transform 1 0 37904 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1626105910
transform 1 0 37812 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_436
timestamp 1626105910
transform 1 0 41216 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_424
timestamp 1626105910
transform 1 0 40112 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_412
timestamp 1626105910
transform 1 0 39008 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_441
timestamp 1626105910
transform 1 0 41676 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_429
timestamp 1626105910
transform 1 0 40572 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1626105910
transform 1 0 40480 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_420
timestamp 1626105910
transform 1 0 39744 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_391
timestamp 1626105910
transform 1 0 37076 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_408
timestamp 1626105910
transform 1 0 38640 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_396
timestamp 1626105910
transform 1 0 37536 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1626105910
transform 1 0 37812 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_400
timestamp 1626105910
transform 1 0 37904 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_391
timestamp 1626105910
transform 1 0 37076 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_400
timestamp 1626105910
transform 1 0 37904 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1626105910
transform 1 0 37812 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_451
timestamp 1626105910
transform 1 0 42596 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_391
timestamp 1626105910
transform 1 0 37076 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_436
timestamp 1626105910
transform 1 0 41216 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_424
timestamp 1626105910
transform 1 0 40112 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_412
timestamp 1626105910
transform 1 0 39008 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_408
timestamp 1626105910
transform 1 0 38640 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_431
timestamp 1626105910
transform 1 0 40756 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1626105910
transform 1 0 40480 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__A
timestamp 1626105910
transform 1 0 40572 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_436
timestamp 1626105910
transform 1 0 41216 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_436
timestamp 1626105910
transform 1 0 41216 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_443
timestamp 1626105910
transform 1 0 41860 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_441
timestamp 1626105910
transform 1 0 41676 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1626105910
transform 1 0 41124 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _052_
timestamp 1626105910
transform -1 0 39744 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_74_420
timestamp 1626105910
transform 1 0 39744 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_419
timestamp 1626105910
transform 1 0 39652 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_424
timestamp 1626105910
transform 1 0 40112 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_412
timestamp 1626105910
transform 1 0 39008 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_429
timestamp 1626105910
transform 1 0 40572 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1626105910
transform 1 0 40480 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_431
timestamp 1626105910
transform 1 0 40756 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_420
timestamp 1626105910
transform 1 0 39744 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_407
timestamp 1626105910
transform 1 0 38548 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_400
timestamp 1626105910
transform 1 0 37904 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_408
timestamp 1626105910
transform 1 0 38640 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1626105910
transform 1 0 38456 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1626105910
transform 1 0 37812 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_402
timestamp 1626105910
transform 1 0 38088 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_390
timestamp 1626105910
transform 1 0 36984 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_396
timestamp 1626105910
transform 1 0 37536 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_391
timestamp 1626105910
transform 1 0 37076 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_396
timestamp 1626105910
transform 1 0 37536 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_441
timestamp 1626105910
transform 1 0 41676 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_429
timestamp 1626105910
transform 1 0 40572 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1626105910
transform 1 0 40480 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_420
timestamp 1626105910
transform 1 0 39744 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_436
timestamp 1626105910
transform 1 0 41216 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_400
timestamp 1626105910
transform 1 0 37904 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1626105910
transform 1 0 37812 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_391
timestamp 1626105910
transform 1 0 37076 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_424
timestamp 1626105910
transform 1 0 40112 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_436
timestamp 1626105910
transform 1 0 41216 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_424
timestamp 1626105910
transform 1 0 40112 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_412
timestamp 1626105910
transform 1 0 39008 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_412
timestamp 1626105910
transform 1 0 39008 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_408
timestamp 1626105910
transform 1 0 38640 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_396
timestamp 1626105910
transform 1 0 37536 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1626105910
transform -1 0 48852 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1626105910
transform -1 0 48852 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1626105910
transform -1 0 48852 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_514
timestamp 1626105910
transform 1 0 48392 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_514
timestamp 1626105910
transform 1 0 48392 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1626105910
transform 1 0 48300 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_510
timestamp 1626105910
transform 1 0 48024 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_506
timestamp 1626105910
transform 1 0 47656 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1626105910
transform 1 0 47564 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_494
timestamp 1626105910
transform 1 0 46552 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_493
timestamp 1626105910
transform 1 0 46460 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_481
timestamp 1626105910
transform 1 0 45356 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_498
timestamp 1626105910
transform 1 0 46920 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_486
timestamp 1626105910
transform 1 0 45816 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1626105910
transform 1 0 46460 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1626105910
transform 1 0 45724 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_489
timestamp 1626105910
transform 1 0 46092 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_477
timestamp 1626105910
transform 1 0 44988 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_465
timestamp 1626105910
transform 1 0 43884 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_469
timestamp 1626105910
transform 1 0 44252 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_457
timestamp 1626105910
transform 1 0 43148 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_465
timestamp 1626105910
transform 1 0 43884 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1626105910
transform 1 0 43792 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_460
timestamp 1626105910
transform 1 0 43424 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_477
timestamp 1626105910
transform 1 0 44988 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1626105910
transform -1 0 48852 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__CLK
timestamp 1626105910
transform 1 0 43148 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1626105910
transform 1 0 43056 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_514
timestamp 1626105910
transform 1 0 48392 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1626105910
transform -1 0 48852 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_514
timestamp 1626105910
transform 1 0 48392 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1626105910
transform 1 0 48300 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1626105910
transform 1 0 47564 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_493
timestamp 1626105910
transform 1 0 46460 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_481
timestamp 1626105910
transform 1 0 45356 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_469
timestamp 1626105910
transform 1 0 44252 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_457
timestamp 1626105910
transform 1 0 43148 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1626105910
transform 1 0 43056 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1626105910
transform 1 0 48300 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1626105910
transform -1 0 48852 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_78_510
timestamp 1626105910
transform 1 0 48024 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_498
timestamp 1626105910
transform 1 0 46920 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_486
timestamp 1626105910
transform 1 0 45816 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1626105910
transform 1 0 45724 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_465
timestamp 1626105910
transform 1 0 43884 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_477
timestamp 1626105910
transform 1 0 44988 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_507
timestamp 1626105910
transform 1 0 47748 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1626105910
transform -1 0 48852 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_514
timestamp 1626105910
transform 1 0 48392 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1626105910
transform 1 0 48300 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1626105910
transform 1 0 47564 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_493
timestamp 1626105910
transform 1 0 46460 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_481
timestamp 1626105910
transform 1 0 45356 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_469
timestamp 1626105910
transform 1 0 44252 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_457
timestamp 1626105910
transform 1 0 43148 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1626105910
transform 1 0 43056 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1626105910
transform 1 0 43056 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1626105910
transform -1 0 48852 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_510
timestamp 1626105910
transform 1 0 48024 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_498
timestamp 1626105910
transform 1 0 46920 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_486
timestamp 1626105910
transform 1 0 45816 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1626105910
transform 1 0 45724 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_465
timestamp 1626105910
transform 1 0 43884 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_477
timestamp 1626105910
transform 1 0 44988 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_459
timestamp 1626105910
transform 1 0 43332 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1626105910
transform -1 0 48852 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_514
timestamp 1626105910
transform 1 0 48392 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1626105910
transform 1 0 48300 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1626105910
transform 1 0 47564 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_493
timestamp 1626105910
transform 1 0 46460 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_481
timestamp 1626105910
transform 1 0 45356 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_469
timestamp 1626105910
transform 1 0 44252 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_457
timestamp 1626105910
transform 1 0 43148 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1626105910
transform 1 0 43056 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_471
timestamp 1626105910
transform 1 0 44436 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1626105910
transform -1 0 48852 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_510
timestamp 1626105910
transform 1 0 48024 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_498
timestamp 1626105910
transform 1 0 46920 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_486
timestamp 1626105910
transform 1 0 45816 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1626105910
transform 1 0 45724 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_484
timestamp 1626105910
transform 1 0 45632 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_476
timestamp 1626105910
transform 1 0 44896 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _116_
timestamp 1626105910
transform 1 0 43332 0 -1 42976
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_74_455
timestamp 1626105910
transform 1 0 42964 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_495
timestamp 1626105910
transform 1 0 46644 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_483
timestamp 1626105910
transform 1 0 45540 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_448
timestamp 1626105910
transform 1 0 42320 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_453
timestamp 1626105910
transform 1 0 42780 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_448
timestamp 1626105910
transform 1 0 42320 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_448
timestamp 1626105910
transform 1 0 42320 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_453
timestamp 1626105910
transform 1 0 42780 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_448
timestamp 1626105910
transform 1 0 42320 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_453
timestamp 1626105910
transform 1 0 42780 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_448
timestamp 1626105910
transform 1 0 42320 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__D
timestamp 1626105910
transform 1 0 42780 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1626105910
transform 1 0 47840 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1626105910
transform -1 0 48852 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1626105910
transform 1 0 48208 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_504
timestamp 1626105910
transform 1 0 47472 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1626105910
transform 1 0 47288 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_486
timestamp 1626105910
transform 1 0 45816 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1626105910
transform 1 0 45724 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_498
timestamp 1626105910
transform 1 0 46920 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_465
timestamp 1626105910
transform 1 0 43884 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_477
timestamp 1626105910
transform 1 0 44988 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_453
timestamp 1626105910
transform 1 0 42780 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_448
timestamp 1626105910
transform 1 0 42320 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_441
timestamp 1626105910
transform 1 0 41676 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_429
timestamp 1626105910
transform 1 0 40572 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1626105910
transform 1 0 40480 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_420
timestamp 1626105910
transform 1 0 39744 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_448
timestamp 1626105910
transform 1 0 42320 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_453
timestamp 1626105910
transform 1 0 42780 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_448
timestamp 1626105910
transform 1 0 42320 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_453
timestamp 1626105910
transform 1 0 42780 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_453
timestamp 1626105910
transform 1 0 42780 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_448
timestamp 1626105910
transform 1 0 42320 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_448
timestamp 1626105910
transform 1 0 42320 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_453
timestamp 1626105910
transform 1 0 42780 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_448
timestamp 1626105910
transform 1 0 42320 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_408
timestamp 1626105910
transform 1 0 38640 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_396
timestamp 1626105910
transform 1 0 37536 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_378
timestamp 1626105910
transform 1 0 35880 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_379
timestamp 1626105910
transform 1 0 35972 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_384
timestamp 1626105910
transform 1 0 36432 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1626105910
transform -1 0 48852 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_510
timestamp 1626105910
transform 1 0 48024 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_498
timestamp 1626105910
transform 1 0 46920 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_486
timestamp 1626105910
transform 1 0 45816 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1626105910
transform 1 0 45724 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_465
timestamp 1626105910
transform 1 0 43884 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_477
timestamp 1626105910
transform 1 0 44988 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_453
timestamp 1626105910
transform 1 0 42780 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_441
timestamp 1626105910
transform 1 0 41676 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_429
timestamp 1626105910
transform 1 0 40572 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1626105910
transform 1 0 40480 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_420
timestamp 1626105910
transform 1 0 39744 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_379
timestamp 1626105910
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_384
timestamp 1626105910
transform 1 0 36432 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_379
timestamp 1626105910
transform 1 0 35972 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_384
timestamp 1626105910
transform 1 0 36432 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_379
timestamp 1626105910
transform 1 0 35972 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_384
timestamp 1626105910
transform 1 0 36432 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_379
timestamp 1626105910
transform 1 0 35972 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_384
timestamp 1626105910
transform 1 0 36432 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1626105910
transform 1 0 35972 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_384
timestamp 1626105910
transform 1 0 36432 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1626105910
transform 1 0 35972 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_384
timestamp 1626105910
transform 1 0 36432 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_389
timestamp 1626105910
transform 1 0 36892 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_384
timestamp 1626105910
transform 1 0 36432 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_379
timestamp 1626105910
transform 1 0 35972 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_384
timestamp 1626105910
transform 1 0 36432 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1626105910
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_408
timestamp 1626105910
transform 1 0 38640 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_396
timestamp 1626105910
transform 1 0 37536 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_384
timestamp 1626105910
transform 1 0 36432 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_372
timestamp 1626105910
transform 1 0 35328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1626105910
transform 1 0 35236 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1626105910
transform 1 0 33396 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_363
timestamp 1626105910
transform 1 0 34500 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1626105910
transform 1 0 32292 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1626105910
transform 1 0 31188 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1626105910
transform 1 0 30084 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1626105910
transform 1 0 29992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_306
timestamp 1626105910
transform 1 0 29256 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_294
timestamp 1626105910
transform 1 0 28152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_282
timestamp 1626105910
transform 1 0 27048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1626105910
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_384
timestamp 1626105910
transform 1 0 36432 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1626105910
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_384
timestamp 1626105910
transform 1 0 36432 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1626105910
transform 1 0 35972 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1626105910
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1626105910
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_384
timestamp 1626105910
transform 1 0 36432 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1626105910
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_270
timestamp 1626105910
transform 1 0 25944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_384
timestamp 1626105910
transform 1 0 36432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1626105910
transform 1 0 36432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_383
timestamp 1626105910
transform 1 0 36340 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_384
timestamp 1626105910
transform 1 0 36432 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1626105910
transform 1 0 35972 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _108_
timestamp 1626105910
transform -1 0 38456 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_47_387
timestamp 1626105910
transform 1 0 36708 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_384
timestamp 1626105910
transform 1 0 36432 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_382
timestamp 1626105910
transform 1 0 36248 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_384
timestamp 1626105910
transform 1 0 36432 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1626105910
transform 1 0 35972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_253
timestamp 1626105910
transform 1 0 24380 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_258
timestamp 1626105910
transform 1 0 24840 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_257
timestamp 1626105910
transform 1 0 24748 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__CLK
timestamp 1626105910
transform -1 0 25024 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_258
timestamp 1626105910
transform 1 0 24840 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_253
timestamp 1626105910
transform 1 0 24380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_258
timestamp 1626105910
transform 1 0 24840 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_253
timestamp 1626105910
transform 1 0 24380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_258
timestamp 1626105910
transform 1 0 24840 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_258
timestamp 1626105910
transform 1 0 24840 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_253
timestamp 1626105910
transform 1 0 24380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_253
timestamp 1626105910
transform 1 0 24380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_258
timestamp 1626105910
transform 1 0 24840 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_253
timestamp 1626105910
transform 1 0 24380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_258
timestamp 1626105910
transform 1 0 24840 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_258
timestamp 1626105910
transform 1 0 24840 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_257
timestamp 1626105910
transform 1 0 24748 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_253
timestamp 1626105910
transform 1 0 24380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_258
timestamp 1626105910
transform 1 0 24840 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1626105910
transform 1 0 24380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1626105910
transform 1 0 24840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_253
timestamp 1626105910
transform 1 0 24380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1626105910
transform 1 0 24840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_253
timestamp 1626105910
transform 1 0 24380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1626105910
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_253
timestamp 1626105910
transform 1 0 24380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1626105910
transform 1 0 24840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_253
timestamp 1626105910
transform 1 0 24380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_258
timestamp 1626105910
transform 1 0 24840 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_253
timestamp 1626105910
transform 1 0 24380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_510
timestamp 1626105910
transform 1 0 48024 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1626105910
transform -1 0 48852 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_514
timestamp 1626105910
transform 1 0 48392 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1626105910
transform 1 0 48300 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_502
timestamp 1626105910
transform 1 0 47288 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_490
timestamp 1626105910
transform 1 0 46184 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_484
timestamp 1626105910
transform 1 0 45632 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B2
timestamp 1626105910
transform 1 0 45448 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B1
timestamp 1626105910
transform 1 0 46000 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_469
timestamp 1626105910
transform 1 0 44252 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_481
timestamp 1626105910
transform 1 0 45356 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_457
timestamp 1626105910
transform 1 0 43148 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1626105910
transform 1 0 43056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_455
timestamp 1626105910
transform 1 0 42964 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_443
timestamp 1626105910
transform 1 0 41860 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_431
timestamp 1626105910
transform 1 0 40756 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _055_
timestamp 1626105910
transform -1 0 40756 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_412
timestamp 1626105910
transform 1 0 39008 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_421
timestamp 1626105910
transform 1 0 39836 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__A
timestamp 1626105910
transform 1 0 39652 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_418
timestamp 1626105910
transform 1 0 39560 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_400
timestamp 1626105910
transform 1 0 37904 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1626105910
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_391
timestamp 1626105910
transform 1 0 37076 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1626105910
transform 1 0 35972 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1626105910
transform 1 0 34868 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_355
timestamp 1626105910
transform 1 0 33764 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1626105910
transform 1 0 32660 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1626105910
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_330
timestamp 1626105910
transform 1 0 31464 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_318
timestamp 1626105910
transform 1 0 30360 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1626105910
transform 1 0 28520 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1626105910
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_286
timestamp 1626105910
transform 1 0 27416 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_294
timestamp 1626105910
transform 1 0 28152 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1626105910
transform -1 0 28152 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_277
timestamp 1626105910
transform 1 0 26588 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_258
timestamp 1626105910
transform 1 0 24840 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_253
timestamp 1626105910
transform 1 0 24380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_258
timestamp 1626105910
transform 1 0 24840 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_253
timestamp 1626105910
transform 1 0 24380 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_258
timestamp 1626105910
transform 1 0 24840 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1626105910
transform 1 0 24380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1626105910
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1626105910
transform 1 0 24380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1626105910
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1626105910
transform 1 0 24380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1626105910
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_265
timestamp 1626105910
transform 1 0 25484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1626105910
transform 1 0 24380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1626105910
transform 1 0 23276 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1626105910
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1626105910
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1626105910
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1626105910
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1626105910
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1626105910
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1626105910
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1626105910
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_163
timestamp 1626105910
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1626105910
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1626105910
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1626105910
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1626105910
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1626105910
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_258
timestamp 1626105910
transform 1 0 24840 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1626105910
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1626105910
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1626105910
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1626105910
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_257
timestamp 1626105910
transform 1 0 24748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1626105910
transform 1 0 12788 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_115
timestamp 1626105910
transform 1 0 11684 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1626105910
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1626105910
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1626105910
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1626105910
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1626105910
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1626105910
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1626105910
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_51
timestamp 1626105910
transform 1 0 5796 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1626105910
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1626105910
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1626105910
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1626105910
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1626105910
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use ACMP  COMP
timestamp 1626105910
transform 1 0 22000 0 1 2000
box 0 0 12564 14476
<< labels >>
rlabel metal2 s 12438 0 12494 800 4 clk
port 1 nsew
rlabel metal2 s 37370 0 37426 800 4 rstn
port 2 nsew
rlabel metal3 s 49200 24896 50000 25016 4 INN
port 3 nsew
rlabel metal3 s 49200 8304 50000 8424 4 INP
port 4 nsew
rlabel metal3 s 49200 41624 50000 41744 4 Q
port 5 nsew
rlabel metal3 s 0 12384 800 12504 4 data[0]
port 6 nsew
rlabel metal3 s 0 17416 800 17536 4 data[1]
port 7 nsew
rlabel metal3 s 0 22448 800 22568 4 data[2]
port 8 nsew
rlabel metal3 s 0 27480 800 27600 4 data[3]
port 9 nsew
rlabel metal3 s 0 32376 800 32496 4 data[4]
port 10 nsew
rlabel metal3 s 0 37408 800 37528 4 data[5]
port 11 nsew
rlabel metal3 s 0 42440 800 42560 4 data[6]
port 12 nsew
rlabel metal3 s 0 47472 800 47592 4 data[7]
port 13 nsew
rlabel metal3 s 0 7352 800 7472 4 done
port 14 nsew
rlabel metal3 s 0 2456 800 2576 4 start
port 15 nsew
rlabel metal4 s 44208 2128 44528 47376 4 VPWR
port 16 nsew
rlabel metal4 s 34208 2176 34528 47376 4 VPWR
port 16 nsew
rlabel metal4 s 24208 2176 24528 47376 4 VPWR
port 16 nsew
rlabel metal4 s 14208 2128 14528 47376 4 VPWR
port 16 nsew
rlabel metal4 s 4208 2128 4528 47376 4 VPWR
port 16 nsew
rlabel metal4 s 39208 2128 39528 47376 4 VGND
port 17 nsew
rlabel metal4 s 29208 2176 29528 47376 4 VGND
port 17 nsew
rlabel metal4 s 19208 2176 19528 47376 4 VGND
port 17 nsew
rlabel metal4 s 9208 2128 9528 47376 4 VGND
port 17 nsew
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string GDS_FILE ../gds/adc.gds
string GDS_END 1346242
string GDS_START 368140
<< end >>
