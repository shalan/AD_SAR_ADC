magic
tech sky130A
magscale 1 2
timestamp 0
<< checkpaint >>
rect -3932 -3932 3933 3933
<< end >>
