* NGSPICE file created from adc_wrapper.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__diode_2 VGND VPWR VPB VNB DIODE
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO VGND VPWR VPB VNB
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND X VPWR A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q VGND CLK VPWR VPB VNB D
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_1 VGND X B1 VPWR B2 A1 A2 VPB VNB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND X VPWR A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND X VPWR A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 RESET_B Q VGND CLK VPWR VPB VNB D
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 RESET_B Q VGND CLK VPWR VPB VNB D
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 VGND Y VPWR A VPB B VNB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 VGND Y VPWR A VPB VNB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_1 VGND X B1 C1 VPWR A1 A2 A3 VPB VNB
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND X B1 VPWR A1 A2 A3 VPB VNB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VGND X VPWR A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND X VPWR A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q VGND CLK VPWR VPB VNB D
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_8 S VGND X A0 VPWR A1 VPB VNB
X0 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_79_21# A0 a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_1259_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_1302_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_792_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1259_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_79_21# A1 a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 VGND a_1259_199# a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_79_21# A0 a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 VPWR S a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_792_297# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1302_47# a_1259_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VPWR a_1259_199# a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_1302_297# a_1259_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_792_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1302_297# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND S a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_79_21# A1 a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 a_792_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 Q VGND CLK VPWR VPB VNB D
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 VGND X VPWR A VPB VNB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND Y B1 VPWR A1 A2 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_1 VGND X B1 VPWR A1 A2 VPB VNB
X0 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 VGND Y VPWR A VPB B VNB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VGND X VPWR A VPB VNB
X0 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND Y VPWR A VPB B VNB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_4 VGND X VPWR A VPB B VNB C D
X0 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND X VPWR A VPB B VNB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hvl__decap_8 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
.ends

.subckt sky130_fd_sc_hvl__decap_4 VGND VPWR VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt sky130_fd_sc_hvl__inv_1 VGND Y VPWR A VPB VNB
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
.ends

.subckt sky130_fd_sc_hvl__diode_2 VGND VPWR VPB VNB DIODE
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 pj=3.16e+06u area=6.072e+11p
.ends

.subckt sky130_fd_sc_hvl__nor3_1 VGND Y VPWR A VPB B VNB C
X0 a_205_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1 a_347_443# B a_205_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2 Y C a_347_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 Y C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 VGND B Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
.ends

.subckt sky130_fd_sc_hvl__nand3_1 VGND Y VPWR A VPB B VNB C
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1 a_243_107# C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2 a_385_107# B a_243_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 Y C VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4 VPWR B Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X5 Y A a_385_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
.ends

.subckt sky130_fd_sc_hvl__inv_4 VGND Y VPWR A VPB VNB
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X6 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
.ends

.subckt ACMP_HVL clk INN INP Q vccd2 vssd2
XFILLER_12_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_9_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx0 vssd2 x0/Y vccd2 clk vccd2 vssd2 sky130_fd_sc_hvl__inv_1
XFILLER_6_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_100 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_15_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XANTENNA_x0_A vssd2 vccd2 vccd2 vssd2 clk sky130_fd_sc_hvl__diode_2
XFILLER_15_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_12_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_135 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_15_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx5 vssd2 Q vccd2 x5/A vccd2 x5/B vssd2 x6/Y sky130_fd_sc_hvl__nor3_1
XFILLER_13_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx2.x1 vssd2 x5/B vccd2 x0/Y vccd2 INP vssd2 x6/B sky130_fd_sc_hvl__nor3_1
XFILLER_13_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx6 vssd2 x6/Y vccd2 x6/A vccd2 x6/B vssd2 Q sky130_fd_sc_hvl__nor3_1
XFILLER_4_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XANTENNA_x2.x1_B vssd2 vccd2 vccd2 vssd2 INP sky130_fd_sc_hvl__diode_2
Xx2.x2 vssd2 x6/B vccd2 x0/Y vccd2 INN vssd2 x5/B sky130_fd_sc_hvl__nor3_1
XFILLER_15_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_4_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_107 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_2_118 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_2_129 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_13_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_5_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_132 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_13_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_124 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XANTENNA_x1.x1_A vssd2 vccd2 vccd2 vssd2 clk sky130_fd_sc_hvl__diode_2
XFILLER_15_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_12_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XANTENNA_x1.x1_B vssd2 vccd2 vccd2 vssd2 INP sky130_fd_sc_hvl__diode_2
XFILLER_2_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_137 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_4_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_5_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_1_107 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_1_118 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_15_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_8_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_129 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_118 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_14_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XANTENNA_x2.x2_B vssd2 vccd2 vccd2 vssd2 INN sky130_fd_sc_hvl__diode_2
XFILLER_5_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_4_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_11_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_8_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_11_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_2_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_2_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_135 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_10_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_5_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_8_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_7_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx1.x1 vssd2 x1.x4/A vccd2 clk vccd2 INP vssd2 x1.x3/A sky130_fd_sc_hvl__nand3_1
XFILLER_14_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_80 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_11_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_15_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx1.x2 vssd2 x1.x3/A vccd2 clk vccd2 INN vssd2 x1.x4/A sky130_fd_sc_hvl__nand3_1
XFILLER_14_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_14_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx1.x3 vssd2 x5/A vccd2 x1.x3/A vccd2 vssd2 sky130_fd_sc_hvl__inv_4
XFILLER_6_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_5_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_9_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
Xx1.x4 vssd2 x6/A vccd2 x1.x4/A vccd2 vssd2 sky130_fd_sc_hvl__inv_4
XFILLER_0_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_72 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_104 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XANTENNA_x1.x2_A vssd2 vccd2 vccd2 vssd2 clk sky130_fd_sc_hvl__diode_2
XFILLER_3_118 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_3_129 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_9_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_13_120 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_10_112 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XANTENNA_x1.x2_B vssd2 vccd2 vccd2 vssd2 INN sky130_fd_sc_hvl__diode_2
XFILLER_3_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_96 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_136 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_4
XFILLER_3_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_12_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_128 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_3_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_9_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_0_56 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_15_64 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
XFILLER_6_88 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hvl__decap_8
.ends

.subckt sky130_fd_sc_hd__buf_2 VGND X VPWR A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_4 VGND X VPWR A VPB B VNB
X0 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_4 VGND X VPWR A VPB B VNB C
X0 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_1 VGND Y VPWR A VPB VNB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND Y C1 B1 VPWR B2 A1 A2 VPB VNB
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221oi_1 VGND Y C1 B1 VPWR B2 A1 A2 VPB VNB
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_1 VGND Y VPWR A VPB B VNB C
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt ACMP INN INP Q VDD VSS clk vccd2 vssd2
XFILLER_23_53 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_12_12 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
Xx2 vssd2 x2/Y vccd2 x6/Y vccd2 vssd2 sky130_fd_sc_hd__inv_1
XFILLER_3_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_x6_B1 vssd2 vccd2 vccd2 vssd2 clk sky130_fd_sc_hd__diode_2
XFILLER_12_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_x9_B1 vssd2 vccd2 vccd2 vssd2 clk sky130_fd_sc_hd__diode_2
XFILLER_3_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
Xx3 vssd2 x3/Y vccd2 x9/Y vccd2 vssd2 sky130_fd_sc_hd__inv_1
XFILLER_23_12 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_36 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_0 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_38 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_12_49 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_8
Xx6 vssd2 x6/Y x9/Y clk vccd2 x9/B2 x7/A2 x7/A2 vccd2 vssd2 sky130_fd_sc_hd__o221ai_1
XFILLER_9_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_15_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_49 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_8
XPHY_1 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
Xx7 vssd2 x7/Y x8/Y x8/B1 vccd2 x8/B2 x7/A2 x7/A2 vccd2 vssd2 sky130_fd_sc_hd__a221oi_1
XFILLER_15_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XPHY_2 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_7_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_4_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
Xx8 vssd2 x8/Y x7/Y x8/B1 vccd2 x8/B2 x9/A2 x9/A2 vccd2 vssd2 sky130_fd_sc_hd__a221oi_1
Xx9 vssd2 x9/Y x6/Y clk vccd2 x9/B2 x9/A2 x9/A2 vccd2 vssd2 sky130_fd_sc_hd__o221ai_1
XPHY_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_4_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_21_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XPHY_4 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_4_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input4_A vssd2 vccd2 vccd2 vssd2 VSS sky130_fd_sc_hd__diode_2
XFILLER_19_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_18_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_5 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_6 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
Xinput1 vssd2 x9/A2 vccd2 INN vccd2 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_10_55 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XPHY_7 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
Xinput2 vssd2 x7/A2 vccd2 INP vccd2 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input2_A vssd2 vccd2 vccd2 vssd2 INP sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_8 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
Xinput3 vssd2 x8/B2 vccd2 VDD vccd2 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_1_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_35 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XPHY_9 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_4_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
Xinput4 vssd2 x9/B2 vccd2 VSS vccd2 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_6 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_49 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_5_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_2_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_8_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_8_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_40 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_11_53 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_55 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_12_6 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_41 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
Xx10 vssd2 x11/A vccd2 x3/Y vccd2 x7/Y vssd2 x11/Y sky130_fd_sc_hd__nor3_1
XFILLER_22_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XPHY_31 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_20 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
Xx11 vssd2 x11/Y vccd2 x11/A vccd2 x2/Y vssd2 x8/Y sky130_fd_sc_hd__nor3_1
XFILLER_22_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_43 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_32 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_21 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_10 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_33 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_44 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_22 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_46 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_11_35 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XPHY_11 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_2_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_35 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_14_46 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XPHY_12 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_45 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_34 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_23 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_8_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_24 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_35 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_46 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_13 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
Xx15 vssd2 x8/B1 vccd2 clk vccd2 vssd2 sky130_fd_sc_hd__inv_1
XFILLER_24_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XPHY_25 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_47 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_36 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA_input3_A vssd2 vccd2 vccd2 vssd2 VDD sky130_fd_sc_hd__diode_2
XPHY_14 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_17_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_37 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_26 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_48 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_15 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_0_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_x15_A vssd2 vccd2 vccd2 vssd2 clk sky130_fd_sc_hd__diode_2
XPHY_27 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_49 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_38 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_16 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_51 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_0_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_39 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XPHY_28 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_22_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_17 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA_input1_A vssd2 vccd2 vccd2 vssd2 INN sky130_fd_sc_hd__diode_2
XFILLER_0_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_29 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_6_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_18 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XPHY_19 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_6_54 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_4
Xoutput5 vssd2 Q vccd2 x11/A vccd2 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_5_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_30 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_42 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd2 vccd2 vccd2 vssd2 sky130_fd_sc_hd__decap_12
.ends

.subckt INV w_n6_n456# w_0_0# a_160_n242# a_n88_n102#
X0 a_160_n242# a_n88_n102# w_n6_n456# w_n6_n456# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=610000u l=150000u
X1 a_160_n242# a_n88_n102# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=150000u
.ends

.subckt switch_layout vout gnd vdd dinb din inp1 inp2 dd
XINV_1 gnd vdd dd dinb INV
XINV_0 gnd vdd dinb din INV
X0 inp1 dd vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1 inp2 dd vout inp2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=150000u
X2 vout dinb inp1 inp1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.21e+06u l=150000u
X3 vout dinb inp2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
.ends

.subckt res250_layout a_238_n246# a_410_n248# w_202_n310#
X0 a_238_n246# a_410_n248# w_202_n310# sky130_fd_pr__res_generic_nd w=295000u l=650000u
.ends

.subckt res500_layout a_238_n246# a_528_n240# w_202_n310#
X0 a_238_n246# a_528_n240# w_202_n310# sky130_fd_pr__res_generic_nd w=270000u l=1.24e+06u
.ends

.subckt x2bitdac_layout out_v x2_vout x1_vout d1 d0 vref5 x2_inp1 x1_inp2 x1_inp1
+ vref1 gnd switch_layout_2/vdd
Xswitch_layout_0 x1_vout gnd switch_layout_2/vdd switch_layout_0/dinb d0 x1_inp1 x1_inp2
+ switch_layout_0/dd switch_layout
Xswitch_layout_1 x2_vout gnd switch_layout_2/vdd switch_layout_1/dinb d0 x2_inp1 vref5
+ switch_layout_1/dd switch_layout
Xswitch_layout_2 out_v gnd switch_layout_2/vdd switch_layout_2/dinb d1 x1_vout x2_vout
+ switch_layout_2/dd switch_layout
Xres500_layout_0 x1_inp1 x1_inp2 gnd res500_layout
Xres500_layout_1 x1_inp2 x2_inp1 gnd res500_layout
Xres500_layout_2 vref1 x1_inp1 gnd res500_layout
Xres250_layout_0 x2_inp1 vref5 gnd res250_layout
.ends

.subckt x3bitdac_layout out_v x2_out_v x1_out_v d2 d1 d0 x2_vref1 x1_vref5 inp1 inp2
+ gnd switch_layout_0/vdd
Xswitch_layout_0 out_v gnd switch_layout_0/vdd switch_layout_0/dinb d2 x1_out_v x2_out_v
+ switch_layout_0/dd switch_layout
X2bitdac_layout_0 x1_out_v 2bitdac_layout_0/x2_vout 2bitdac_layout_0/x1_vout d1 d0
+ x1_vref5 2bitdac_layout_0/x2_inp1 2bitdac_layout_0/x1_inp2 2bitdac_layout_0/x1_inp1
+ inp1 gnd switch_layout_0/vdd x2bitdac_layout
X2bitdac_layout_1 x2_out_v 2bitdac_layout_1/x2_vout 2bitdac_layout_1/x1_vout d1 d0
+ inp2 2bitdac_layout_1/x2_inp1 2bitdac_layout_1/x1_inp2 2bitdac_layout_1/x1_inp1
+ x2_vref1 gnd switch_layout_0/vdd x2bitdac_layout
Xres250_layout_0 x1_vref5 x2_vref1 gnd res250_layout
.ends

.subckt x4bitdac_layout x1_out_v x2_out_v inp1 inp2 x1_vref5 x2_vref1 d0 d1 d2 d3
+ out_v gnd vdd
Xswitch_layout_0 out_v gnd vdd switch_layout_0/dinb d3 x1_out_v x2_out_v switch_layout_0/dd
+ switch_layout
X3bitdac_layout_0 x1_out_v 3bitdac_layout_0/x2_out_v 3bitdac_layout_0/x1_out_v d2
+ d1 d0 3bitdac_layout_0/x2_vref1 3bitdac_layout_0/x1_vref5 inp1 x1_vref5 gnd vdd
+ x3bitdac_layout
X3bitdac_layout_1 x2_out_v 3bitdac_layout_1/x2_out_v 3bitdac_layout_1/x1_out_v d2
+ d1 d0 3bitdac_layout_1/x2_vref1 3bitdac_layout_1/x1_vref5 x2_vref1 inp2 gnd vdd
+ x3bitdac_layout
Xres250_layout_0 x2_vref1 x1_vref5 gnd res250_layout
.ends

.subckt x5bitdac_layout inp2 inp1 x1_out_v x2_out_v out_v d4 d3 d2 d1 d0 x2_vref1
+ x1_vref5 gnd vdd
Xswitch_layout_0 out_v gnd vdd switch_layout_0/dinb d4 x1_out_v x2_out_v switch_layout_0/dd
+ switch_layout
Xres250_layout_0 x1_vref5 x2_vref1 gnd res250_layout
X4bitdac_layout_0 4bitdac_layout_0/x1_out_v 4bitdac_layout_0/x2_out_v inp1 x1_vref5
+ 4bitdac_layout_0/x1_vref5 4bitdac_layout_0/x2_vref1 d0 d1 d2 d3 x1_out_v gnd vdd
+ x4bitdac_layout
X4bitdac_layout_1 4bitdac_layout_1/x1_out_v 4bitdac_layout_1/x2_out_v x2_vref1 inp2
+ 4bitdac_layout_1/x1_vref5 4bitdac_layout_1/x2_vref1 d0 d1 d2 d3 x2_out_v gnd vdd
+ x4bitdac_layout
.ends

.subckt x6bitdac_layout d4 d3 d2 d1 d0 inp1 inp2 x2_vref1 x1_vref5 x2_out_v x1_out_v
+ d5 out_v gnd vdd
Xswitch_layout_0 out_v gnd vdd switch_layout_0/dinb d5 x1_out_v x2_out_v switch_layout_0/dd
+ switch_layout
Xres250_layout_0 x1_vref5 x2_vref1 gnd res250_layout
X5bitdac_layout_0 x1_vref5 inp1 5bitdac_layout_0/x1_out_v 5bitdac_layout_0/x2_out_v
+ x1_out_v d4 d3 d2 d1 d0 5bitdac_layout_0/x2_vref1 5bitdac_layout_0/x1_vref5 gnd
+ vdd x5bitdac_layout
X5bitdac_layout_1 inp2 x2_vref1 5bitdac_layout_1/x1_out_v 5bitdac_layout_1/x2_out_v
+ x2_out_v d4 d3 d2 d1 d0 5bitdac_layout_1/x2_vref1 5bitdac_layout_1/x1_vref5 gnd
+ vdd x5bitdac_layout
.ends

.subckt x7bitdac_layout d2 d5 d4 d3 d1 d0 x1_out_v x2_out_v out_v d6 inp1 inp2 x2_vref1
+ x1_vref5 gnd vdd
Xswitch_layout_0 out_v gnd vdd switch_layout_0/dinb d6 x1_out_v x2_out_v switch_layout_0/dd
+ switch_layout
X6bitdac_layout_0 d4 d3 d2 d1 d0 x2_vref1 inp2 6bitdac_layout_0/x2_vref1 6bitdac_layout_0/x1_vref5
+ 6bitdac_layout_0/x2_out_v 6bitdac_layout_0/x1_out_v d5 x2_out_v gnd vdd x6bitdac_layout
X6bitdac_layout_1 d4 d3 d2 d1 d0 inp1 x1_vref5 6bitdac_layout_1/x2_vref1 6bitdac_layout_1/x1_vref5
+ 6bitdac_layout_1/x2_out_v 6bitdac_layout_1/x1_out_v d5 x1_out_v gnd vdd x6bitdac_layout
Xres250_layout_0 x1_vref5 x2_vref1 gnd res250_layout
.ends

.subckt DAC_8BIT d0 d1 d2 d3 d4 d5 d6 x2_out_v x1_out_v out_v d7 inp1 x2_vref1 x1_vref5
+ gnd inp2 vdd
Xswitch_layout_0 out_v gnd vdd switch_layout_0/dinb d7 x1_out_v x2_out_v switch_layout_0/dd
+ switch_layout
X7bitdac_layout_0 d2 d5 d4 d3 d1 d0 7bitdac_layout_0/x1_out_v 7bitdac_layout_0/x2_out_v
+ x2_out_v d6 x2_vref1 inp2 7bitdac_layout_0/x2_vref1 7bitdac_layout_0/x1_vref5 gnd
+ vdd x7bitdac_layout
X7bitdac_layout_1 d2 d5 d4 d3 d1 d0 7bitdac_layout_1/x1_out_v 7bitdac_layout_1/x2_out_v
+ x1_out_v d6 inp1 x1_vref5 7bitdac_layout_1/x2_vref1 7bitdac_layout_1/x1_vref5 gnd
+ vdd x7bitdac_layout
Xres250_layout_0 x1_vref5 x2_vref1 gnd res250_layout
.ends

.subckt adc_wrapper analog_io[10] analog_io[11] analog_io[12] analog_io[8] analog_io[9]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_out[15] io_out[16] io_out[17] io_out[18] analog_io[16] analog_io[13]
+ analog_io[14] analog_io[15] io_oeb[19] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23]
+ io_in[20] io_in[21] io_in[22] io_in[23] io_out[19] io_out[20] io_out[21] io_out[22]
+ io_out[23] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[1] wbs_adr_i[2] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7]
+ wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12]
+ wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[1] wbs_dat_i[2]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[1] wbs_dat_o[2] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_adr_i[18] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_adr_i[19]
+ wbs_dat_i[30] wbs_dat_i[31] la_oenb[0] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] la_oenb[1] wbs_adr_i[30] wbs_adr_i[31] la_oenb[2] wbs_dat_o[17] wbs_dat_o[18]
+ wbs_dat_o[19] la_oenb[3] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23]
+ wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29]
+ la_oenb[4] wbs_dat_o[30] wbs_dat_o[31] la_oenb[5] la_data_in[0] la_data_in[1] la_data_in[2]
+ la_data_in[3] la_data_in[4] la_data_in[5] la_data_out[0] la_data_out[1] la_data_out[2]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] la_data_in[26] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_in[15] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_in[16] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[10] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_data_in[20] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_data_in[21] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_data_in[22] la_data_in[39] la_oenb[45] la_data_in[40] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_in[41] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_in[42] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_oenb[46] la_oenb[38]
+ la_oenb[39] la_oenb[37] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_oenb[44] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_oenb[26]
+ la_oenb[27] la_oenb[28] la_oenb[29] la_data_in[38] la_oenb[30] la_oenb[31] la_oenb[32]
+ la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_out[47] la_data_out[48] la_data_out[49] la_data_in[64]
+ la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_in[65] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_in[66] la_data_in[67] la_data_in[72]
+ la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78]
+ la_data_in[79] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[69] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_data_out[68] la_data_out[69]
+ la_data_in[70] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_in[71] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_in[68] la_oenb[88] la_oenb[89]
+ la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96]
+ la_oenb[97] la_oenb[98] la_oenb[99] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[100] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94]
+ la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[93] la_data_out[106] la_data_out[94] la_data_out[107] la_data_out[95]
+ la_data_out[96] la_data_out[108] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[92] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_data_in[88] la_data_in[89] la_data_out[88]
+ la_data_out[89] la_data_out[90] la_data_out[91] la_data_in[119] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_in[116] la_data_in[117] la_data_out[123]
+ la_data_in[112] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_in[118] la_oenb[109] la_data_in[120] la_oenb[110] la_data_in[121] la_oenb[111]
+ la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_data_in[122] la_data_in[123] la_oenb[120] la_oenb[121] la_oenb[122]
+ la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_out[110] user_clock2 user_irq[0]
+ la_data_in[113] user_irq[1] la_data_in[114] user_irq[2] la_data_out[111] la_data_out[112]
+ la_data_out[109] la_data_in[109] la_data_out[113] la_data_in[110] la_data_out[114]
+ la_oenb[108] la_data_out[115] la_data_out[116] la_data_in[111] la_data_out[117]
+ la_data_in[115] la_data_out[118] la_data_out[119] analog_io[2] analog_io[3] analog_io[4]
+ analog_io[5] analog_io[6] analog_io[7] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[9] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[8] io_oeb[9]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[8] io_out[9] analog_io[22]
+ analog_io[23] analog_io[17] analog_io[18] analog_io[19] io_oeb[24] io_oeb[25] io_oeb[26]
+ io_oeb[27] io_oeb[28] io_oeb[29] analog_io[20] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[30] io_in[30] analog_io[21] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] analog_io[27]
+ analog_io[28] analog_io[24] analog_io[25] analog_io[26] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_oeb[30] io_oeb[31] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_oeb[32] io_oeb[33] io_in[8]
+ analog_io[1] io_oeb[2] io_oeb[0] io_out[1] io_in[2] analog_io[0] io_in[1] io_in[0]
+ io_in[3] io_oeb[1] io_out[2] io_in[4] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_in[5] io_in[6] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[0] io_in[7]
+ vssd2 vccd1 vccd2
XFILLER_23_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1497 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_431 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_639 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_241_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_36 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input127_A vssd2 vccd1 vccd1 vssd2 la_data_in[64] sky130_fd_sc_hd__diode_2
XFILLER_172_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1160 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_35_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_187_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input92_A vssd2 vccd1 vccd1 vssd2 la_data_in[32] sky130_fd_sc_hd__diode_2
XFILLER_35_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_294_ _294_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_220_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_89 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_973 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_240_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput401 vssd2 io_oeb[5] vccd1 _112_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput412 vssd2 io_out[15] vccd1 _132_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput423 vssd2 io_out[25] vccd1 _142_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_218_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput434 vssd2 io_out[35] vccd1 _347_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput445 vssd2 la_data_out[100] vccd1 _244_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput456 vssd2 la_data_out[110] vccd1 _254_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput467 vssd2 la_data_out[120] vccd1 _264_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput478 vssd2 la_data_out[15] vccd1 _159_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_141_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput489 vssd2 la_data_out[25] vccd1 _169_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_60_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_2286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_916 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_927 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_225_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_128_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input244_A vssd2 vccd1 vccd1 vssd2 la_oenb[54] sky130_fd_sc_hd__diode_2
XFILLER_238_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_160_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_61_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_202_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_346_ _346_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _346_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_277_ _277_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_127_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_170_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_696 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_108_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_151_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_386 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1769 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2359 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_25_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1371 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_713 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_724 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_757 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_123_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_200_ _200_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_130_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_131_ _131_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_240_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_201_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input194_A vssd2 vccd1 vccd1 vssd2 la_oenb[124] sky130_fd_sc_hd__diode_2
XFILLER_201_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_062_ vssd2 _351_/D _351_/Q vccd1 _341_/Q _352_/Q _055_/A vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_193_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_611 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_388 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_137_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input361_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[9] sky130_fd_sc_hd__diode_2
XFILLER_180_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_655 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_140_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input55_A vssd2 vccd1 vccd1 vssd2 la_data_in[114] sky130_fd_sc_hd__diode_2
XFILLER_79_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_4_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_329_ vssd2 _329_/X vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2212 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1566 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_162_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_49 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2009 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__351__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_5_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input207_A vssd2 vccd1 vccd1 vssd2 la_oenb[20] sky130_fd_sc_hd__diode_2
XFILLER_245_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_34_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_521 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_160_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_54_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_554 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XPHY_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_587 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_598 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_114_ _114_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_184_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__312__A vssd2 vccd1 vccd1 vssd2 _316_/A sky130_fd_sc_hd__diode_2
XFILLER_226_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_57_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1639 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_183_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1578 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__080__A1 vssd2 vccd1 vccd1 vssd2 _099_/A sky130_fd_sc_hd__diode_2
XFILLER_169_9 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1173 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_198_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_201_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_231_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input157_A vssd2 vccd1 vccd1 vssd2 la_data_in[91] sky130_fd_sc_hd__diode_2
XFILLER_7_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput301 vssd2 input301/X vccd1 wbs_adr_i[13] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput312 vssd2 input312/X vccd1 wbs_adr_i[23] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput323 vssd2 input323/X vccd1 wbs_adr_i[4] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_7_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput334 vssd2 input334/X vccd1 wbs_dat_i[13] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput345 vssd2 input345/X vccd1 wbs_dat_i[23] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_102_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput356 vssd2 input356/X vccd1 wbs_dat_i[4] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput367 vssd2 input367/X vccd1 wbs_we_i vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_152_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input324_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[5] sky130_fd_sc_hd__diode_2
XFILLER_229_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input18_A vssd2 vccd1 vccd1 vssd2 io_in[25] sky130_fd_sc_hd__diode_2
XFILLER_57_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1285 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_362 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_373 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_395 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1948 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_54_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__062__A1 vssd2 vccd1 vccd1 vssd2 _352_/Q sky130_fd_sc_hd__diode_2
XFILLER_228_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__062__B2 vssd2 vccd1 vccd1 vssd2 _341_/Q sky130_fd_sc_hd__diode_2
XFILLER_184_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_91_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_223_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_668 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_2_2104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_213_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2054 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1375 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1160 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input274_A vssd2 vccd1 vccd1 vssd2 la_oenb[81] sky130_fd_sc_hd__diode_2
XFILLER_5_558 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_181_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput120 vssd2 input120/X vccd1 la_data_in[58] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_209_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput131 vssd2 input131/X vccd1 la_data_in[68] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_7_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput142 vssd2 input142/X vccd1 la_data_in[78] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput153 vssd2 input153/X vccd1 la_data_in[88] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_79_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput164 vssd2 input164/X vccd1 la_data_in[98] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_64_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput175 vssd2 input175/X vccd1 la_oenb[107] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput186 vssd2 input186/X vccd1 la_oenb[117] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_1900 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput197 vssd2 input197/X vccd1 la_oenb[127] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_5_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1944 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_18_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput605 vssd2 wbs_dat_o[7] vccd1 _283_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_161_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_172_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_131_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_165_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_161_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_293_ _293_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_220_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input85_A vssd2 vccd1 vccd1 vssd2 la_data_in[26] sky130_fd_sc_hd__diode_2
XFILLER_127_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_81_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_174_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_133_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1741 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_17_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput402 vssd2 io_oeb[6] vccd1 _113_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_145_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput413 vssd2 io_out[16] vccd1 _133_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput424 vssd2 io_out[26] vccd1 _336_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput435 vssd2 io_out[36] vccd1 _348_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_216_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput446 vssd2 la_data_out[101] vccd1 _245_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput457 vssd2 la_data_out[111] vccd1 _255_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput468 vssd2 la_data_out[121] vccd1 _265_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput479 vssd2 la_data_out[16] vccd1 _160_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_60_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__320__A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_214_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_362 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_671 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_23_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_928 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input237_A vssd2 vccd1 vccd1 vssd2 la_oenb[48] sky130_fd_sc_hd__diode_2
XFILLER_58_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_186_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_345_ _345_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _345_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_159_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_276_ _276_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_195_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_110_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_68 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_231_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1748 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__315__A vssd2 vccd1 vccd1 vssd2 _316_/A sky130_fd_sc_hd__diode_2
XFILLER_222_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_116_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_151_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_55_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1383 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_725 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_736 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_758 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_123_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_769 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_130_ _130_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_32_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_061_ vssd2 _352_/D _352_/Q vccd1 _056_/X _353_/Q _055_/A vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_109_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input187_A vssd2 vccd1 vccd1 vssd2 la_oenb[118] sky130_fd_sc_hd__diode_2
XFILLER_192_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_180_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input354_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[31] sky130_fd_sc_hd__diode_2
XFILLER_2_133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_667 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_156_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input48_A vssd2 vccd1 vccd1 vssd2 la_data_in[108] sky130_fd_sc_hd__diode_2
XFILLER_120_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_43_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_4_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_328_ vssd2 _328_/X vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_259_ _259_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_7_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1545 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1388 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_178_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_216_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_2135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1401 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_500 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_31_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input102_A vssd2 vccd1 vccd1 vssd2 la_data_in[41] sky130_fd_sc_hd__diode_2
XPHY_511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_34_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_533 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_54_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_566 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_141_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_599 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_113_ _113_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_156_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_976 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_124_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_228_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_201_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_116_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_113_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_96_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_38_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2021 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_65_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__080__A2 vssd2 vccd1 vccd1 vssd2 _099_/B sky130_fd_sc_hd__diode_2
XFILLER_181_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1342 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_153_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_530 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput302 vssd2 input302/X vccd1 wbs_adr_i[14] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_7_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput313 vssd2 input313/X vccd1 wbs_adr_i[24] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput324 vssd2 input324/X vccd1 wbs_adr_i[5] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput335 vssd2 input335/X vccd1 wbs_dat_i[14] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_195_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_489 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_29_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput346 vssd2 input346/X vccd1 wbs_dat_i[24] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput357 vssd2 input357/X vccd1 wbs_dat_i[5] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_102_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input317_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[28] sky130_fd_sc_hd__diode_2
XFILLER_229_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_72_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_186_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_330 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_213_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_374 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_201_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_201_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA__062__A2 vssd2 vccd1 vccd1 vssd2 _055_/A sky130_fd_sc_hd__diode_2
XFILLER_169_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_195_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__341__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_191_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__323__A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_239_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_2341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1415 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_54_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_1387 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_109_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_202_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input267_A vssd2 vccd1 vccd1 vssd2 la_oenb[75] sky130_fd_sc_hd__diode_2
XFILLER_235_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_231_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput110 vssd2 input110/X vccd1 la_data_in[49] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput121 vssd2 input121/X vccd1 la_data_in[59] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_44_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input30_A vssd2 vccd1 vccd1 vssd2 io_in[36] sky130_fd_sc_hd__diode_2
XFILLER_76_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput132 vssd2 input132/X vccd1 la_data_in[69] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput143 vssd2 input143/X vccd1 la_data_in[79] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput154 vssd2 input154/X vccd1 la_data_in[89] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput165 vssd2 input165/X vccd1 la_data_in[99] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_79_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput176 vssd2 input176/X vccd1 la_oenb[108] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_36_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput187 vssd2 input187/X vccd1 la_oenb[118] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_63_205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput198 vssd2 input198/X vccd1 la_oenb[12] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_91_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1960 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_160 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_171 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_18_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output486_A vssd2 vccd1 vccd1 vssd2 _166_/LO sky130_fd_sc_hd__diode_2
XPHY_193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_195_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput606 vssd2 wbs_dat_o[8] vccd1 _284_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_113_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_98_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_141_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA__318__A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_62_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__053__A vssd2 vccd1 vccd1 vssd2 _075_/A sky130_fd_sc_hd__diode_2
XFILLER_163_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_77_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_374 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_1184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_227_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1256 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_54_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_159_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_292_ _292_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_139_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input78_A vssd2 vccd1 vccd1 vssd2 la_data_in[1] sky130_fd_sc_hd__diode_2
XFILLER_13_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_170_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_123_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_36 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_90 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_224_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_140_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput403 vssd2 io_oeb[7] vccd1 _308_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_145_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput414 vssd2 io_out[17] vccd1 _134_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput425 vssd2 io_out[27] vccd1 _337_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput436 vssd2 io_out[37] vccd1 _349_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput447 vssd2 la_data_out[102] vccd1 _246_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_216_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput458 vssd2 la_data_out[112] vccd1 _256_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput469 vssd2 la_data_out[122] vccd1 _266_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_214_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_234_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_374 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_171 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_97_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_907 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_929 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_184_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_274 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input132_A vssd2 vccd1 vccd1 vssd2 la_data_in[69] sky130_fd_sc_hd__diode_2
XFILLER_246_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_54_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_204_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_344_ _344_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _344_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_275_ _275_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_139_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_127_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_366 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_1550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1414 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_166_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_530 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__331__A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_99_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_59_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1395 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_704 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_715 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_737 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_748 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_060_ vssd2 _353_/D _353_/Q vccd1 _056_/X _354_/Q _055_/A vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_99_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_195_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_82_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_234_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_79_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input347_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[25] sky130_fd_sc_hd__diode_2
XFILLER_120_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_327_ vssd2 _327_/X vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_258_ _258_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_10_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_116_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_189_ _189_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_48_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_390 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_217_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_168_2002 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__092__B1 vssd2 vccd1 vccd1 vssd2 _343_/Q sky130_fd_sc_hd__diode_2
XFILLER_0_2225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_65_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1557 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__326__A vssd2 vccd1 vccd1 vssd2 _326_/A sky130_fd_sc_hd__diode_2
XFILLER_222_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2147 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_85_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__083__B1 vssd2 vccd1 vccd1 vssd2 _346_/Q sky130_fd_sc_hd__diode_2
XFILLER_18_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_501 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_545 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_140_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_34_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_578 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_141_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input297_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[0] sky130_fd_sc_hd__diode_2
X_112_ _112_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_123_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input60_A vssd2 vccd1 vccd1 vssd2 la_data_in[119] sky130_fd_sc_hd__diode_2
XFILLER_193_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_175_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_235_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_75_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1899 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_203_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_188_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2204 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_96_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__080__A3 vssd2 vccd1 vccd1 vssd2 _356_/Q sky130_fd_sc_hd__diode_2
XFILLER_52_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_228_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__056__A vssd2 vccd1 vccd1 vssd2 _341_/Q sky130_fd_sc_hd__diode_2
XFILLER_178_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput303 vssd2 input303/X vccd1 wbs_adr_i[15] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput314 vssd2 input314/X vccd1 wbs_adr_i[25] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_0_468 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput325 vssd2 input325/X vccd1 wbs_adr_i[6] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput336 vssd2 input336/X vccd1 wbs_dat_i[15] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput347 vssd2 input347/X vccd1 wbs_dat_i[25] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput358 vssd2 input358/X vccd1 wbs_dat_i[6] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_378 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input212_A vssd2 vccd1 vccd1 vssd2 la_oenb[25] sky130_fd_sc_hd__diode_2
XFILLER_45_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_331 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_342 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_213_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_375 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_386 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_113_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output431_A vssd2 vccd1 vccd1 vssd2 _344_/Q sky130_fd_sc_hd__diode_2
XFILLER_239_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_182_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_2001 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1300 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_131_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_107_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input162_A vssd2 vccd1 vccd1 vssd2 la_data_in[96] sky130_fd_sc_hd__diode_2
XFILLER_235_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput100 vssd2 input100/X vccd1 la_data_in[3] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput111 vssd2 input111/X vccd1 la_data_in[4] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput122 vssd2 input122/X vccd1 la_data_in[5] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_672 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput133 vssd2 input133/X vccd1 la_data_in[6] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput144 vssd2 input144/X vccd1 la_data_in[7] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput155 vssd2 input155/X vccd1 la_data_in[8] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput166 vssd2 input166/X vccd1 la_data_in[9] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_5_1040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput177 vssd2 input177/X vccd1 la_oenb[109] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input23_A vssd2 vccd1 vccd1 vssd2 io_in[2] sky130_fd_sc_hd__diode_2
XFILLER_79_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput188 vssd2 input188/X vccd1 la_oenb[119] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput199 vssd2 input199/X vccd1 la_oenb[13] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_17_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_103_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_220_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_138_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput607 vssd2 wbs_dat_o[9] vccd1 _285_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_36 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_51_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_489 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_31_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_175_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__334__A vssd2 vccd1 vccd1 vssd2 _335_/A sky130_fd_sc_hd__diode_2
XFILLER_219_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_386 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_199_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_202_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_291_ _291_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_139_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_530 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2357 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_3_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_95_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_378 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput404 vssd2 io_oeb[8] vccd1 _309_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput415 vssd2 io_out[18] vccd1 _135_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput426 vssd2 io_out[28] vccd1 _143_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput437 vssd2 io_out[3] vccd1 _120_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput448 vssd2 la_data_out[103] vccd1 _247_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_160_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput459 vssd2 la_data_out[113] vccd1 _257_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_153_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_228_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_386 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__329__A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_227_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_908 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_919 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_221_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__064__A vssd2 vccd1 vccd1 vssd2 _357_/Q sky130_fd_sc_hd__diode_2
XFILLER_164_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_704 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__354__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_144_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1028 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input125_A vssd2 vccd1 vccd1 vssd2 la_data_in[62] sky130_fd_sc_hd__diode_2
XFILLER_170_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_343_ _343_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _343_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_186_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_202_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input90_A vssd2 vccd1 vccd1 vssd2 la_data_in[30] sky130_fd_sc_hd__diode_2
X_274_ _274_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_10_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_139_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_143 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_142_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_142_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2217 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_65_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_221_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2042 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_55_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_716 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_162_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XPHY_749 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_117_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_215_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input242_A vssd2 vccd1 vccd1 vssd2 la_oenb[52] sky130_fd_sc_hd__diode_2
XFILLER_120_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_38 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_326_ vssd2 _326_/X vccd1 _326_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_257_ _257_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_31_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_188_ _188_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_7_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_174_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_680 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_69_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2204 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA__092__A1 vssd2 vccd1 vccd1 vssd2 _075_/A sky130_fd_sc_hd__diode_2
XFILLER_59_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__083__A1 vssd2 vccd1 vccd1 vssd2 _099_/A sky130_fd_sc_hd__diode_2
XFILLER_18_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_502 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_513 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_546 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_34_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_557 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_34_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_111_ _111_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_138_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input192_A vssd2 vccd1 vccd1 vssd2 la_oenb[122] sky130_fd_sc_hd__diode_2
XFILLER_138_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input53_A vssd2 vccd1 vccd1 vssd2 la_data_in[112] sky130_fd_sc_hd__diode_2
XFILLER_175_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_78_234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_132_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_169_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1834 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_228_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_186 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_1856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_235_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_309_ vssd2 _309_/X vccd1 _316_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_131_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2216 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2001 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_38_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_92 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__337__A vssd2 vccd1 vccd1 vssd2 _337_/A sky130_fd_sc_hd__diode_2
XFILLER_224_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_193_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__072__A vssd2 vccd1 vccd1 vssd2 _072_/A sky130_fd_sc_hd__diode_2
XFILLER_146_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_161_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput304 vssd2 input304/X vccd1 wbs_adr_i[16] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput315 vssd2 input315/X vccd1 wbs_adr_i[26] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput326 vssd2 input326/X vccd1 wbs_adr_i[7] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_357 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput337 vssd2 input337/X vccd1 wbs_dat_i[16] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput348 vssd2 input348/X vccd1 wbs_dat_i[26] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput359 vssd2 input359/X vccd1 wbs_dat_i[7] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_84_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input205_A vssd2 vccd1 vccd1 vssd2 la_oenb[19] sky130_fd_sc_hd__diode_2
XFILLER_72_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_101_60 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_213_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_387 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output424_A vssd2 vccd1 vccd1 vssd2 _336_/X sky130_fd_sc_hd__diode_2
XFILLER_239_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_187_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_74_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_34_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_476 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2013 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_701 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_123_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input155_A vssd2 vccd1 vccd1 vssd2 la_data_in[8] sky130_fd_sc_hd__diode_2
XFILLER_103_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput101 vssd2 input101/X vccd1 la_data_in[40] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput112 vssd2 input112/X vccd1 la_data_in[50] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_44_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput123 vssd2 input123/X vccd1 la_data_in[60] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput134 vssd2 input134/X vccd1 la_data_in[70] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput145 vssd2 input145/X vccd1 la_data_in[80] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput156 vssd2 input156/X vccd1 la_data_in[90] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput167 vssd2 input167/X vccd1 la_oenb[0] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input322_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[3] sky130_fd_sc_hd__diode_2
Xinput178 vssd2 input178/X vccd1 la_oenb[10] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_166_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput189 vssd2 input189/X vccd1 la_oenb[11] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_56_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input16_A vssd2 vccd1 vccd1 vssd2 io_in[23] sky130_fd_sc_hd__diode_2
XFILLER_63_218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1085 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_31_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_173 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_822 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_402 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_35_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_88 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_117_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_8_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input8_A vssd2 vccd1 vccd1 vssd2 io_in[16] sky130_fd_sc_hd__diode_2
XFILLER_230_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_85_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1131 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_73_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_187_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_476 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_290_ _290_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_186_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input272_A vssd2 vccd1 vccd1 vssd2 la_oenb[7] sky130_fd_sc_hd__diode_2
XFILLER_170_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_135_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_542 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_172_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_229_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_17_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput405 vssd2 io_oeb[9] vccd1 _310_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput416 vssd2 io_out[19] vccd1 _136_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_138_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput427 vssd2 io_out[29] vccd1 _338_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput438 vssd2 io_out[4] vccd1 _121_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput449 vssd2 la_data_out[104] vccd1 _248_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_67_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_28_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_97_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_149_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_407 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_232_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1000 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input118_A vssd2 vccd1 vccd1 vssd2 la_data_in[56] sky130_fd_sc_hd__diode_2
XFILLER_163_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_21 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_342_ _342_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _342_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_186_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_941 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_273_ _273_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_10_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input83_A vssd2 vccd1 vccd1 vssd2 la_data_in[24] sky130_fd_sc_hd__diode_2
XFILLER_10_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_155 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_178_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_177_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_102_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_247_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_717 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_728 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_204 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__075__A vssd2 vccd1 vccd1 vssd2 _075_/A sky130_fd_sc_hd__diode_2
XFILLER_225_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input235_A vssd2 vccd1 vccd1 vssd2 la_oenb[46] sky130_fd_sc_hd__diode_2
XFILLER_120_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_17 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_100_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_62_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_64 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_325_ vssd2 _325_/X vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_256_ _256_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_431 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_187_ _187_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_49_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_77_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__092__A2 vssd2 vccd1 vccd1 vssd2 _076_/A sky130_fd_sc_hd__diode_2
XFILLER_59_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2072 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__344__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_222_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__083__A2 vssd2 vccd1 vccd1 vssd2 _099_/B sky130_fd_sc_hd__diode_2
XFILLER_217_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_525 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_558 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_34_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_110_ _110_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_211_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input185_A vssd2 vccd1 vccd1 vssd2 la_oenb[116] sky130_fd_sc_hd__diode_2
XFILLER_138_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_88 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_166_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input352_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[2] sky130_fd_sc_hd__diode_2
XFILLER_106_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_64 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_105_395 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input46_A vssd2 vccd1 vccd1 vssd2 la_data_in[106] sky130_fd_sc_hd__diode_2
XFILLER_132_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_15_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_308_ vssd2 _308_/X vccd1 _316_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_175_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_239_ _239_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_152_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_58_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_113_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_228_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput305 vssd2 input305/X vccd1 wbs_adr_i[17] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput316 vssd2 input316/X vccd1 wbs_adr_i[27] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_48_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput327 vssd2 input327/X vccd1 wbs_adr_i[8] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput338 vssd2 input338/X vccd1 wbs_dat_i[17] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput349 vssd2 input349/X vccd1 wbs_dat_i[27] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input100_A vssd2 vccd1 vccd1 vssd2 la_data_in[3] sky130_fd_sc_hd__diode_2
XPHY_300 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_366 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_388 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_8_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_193_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1643 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_207_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_639 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_374 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_98_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_131_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_111_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1131 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_54_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_179_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_139_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput102 vssd2 input102/X vccd1 la_data_in[41] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput113 vssd2 input113/X vccd1 la_data_in[51] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput124 vssd2 input124/X vccd1 la_data_in[61] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput135 vssd2 input135/X vccd1 la_data_in[71] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input148_A vssd2 vccd1 vccd1 vssd2 la_data_in[83] sky130_fd_sc_hd__diode_2
XFILLER_236_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput146 vssd2 input146/X vccd1 la_data_in[81] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput157 vssd2 input157/X vccd1 la_data_in[91] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput168 vssd2 input168/X vccd1 la_oenb[100] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput179 vssd2 input179/X vccd1 la_oenb[110] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_166_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_56_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1915 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input315_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[26] sky130_fd_sc_hd__diode_2
XFILLER_2_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_56_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_56_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_214_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_374 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_834 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_411 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_246_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1143 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_139_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1857 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input265_A vssd2 vccd1 vccd1 vssd2 la_oenb[73] sky130_fd_sc_hd__diode_2
XFILLER_122_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_194_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_114_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_190_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1712 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_411 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1756 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1793 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_103_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput406 vssd2 io_out[0] vccd1 _117_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput417 vssd2 io_out[1] vccd1 _118_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_138_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput428 vssd2 io_out[2] vccd1 _119_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput439 vssd2 io_out[5] vccd1 _122_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_218_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_110_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1502 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1546 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_419 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_132_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1045 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_341_ _105_/A _341_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _341_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_241_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_33 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_272_ _272_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_953 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA_input76_A vssd2 vccd1 vccd1 vssd2 la_data_in[18] sky130_fd_sc_hd__diode_2
XFILLER_13_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_182_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2200 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1590 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_221_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_440 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_99_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__095__B1 vssd2 vccd1 vccd1 vssd2 _342_/Q sky130_fd_sc_hd__diode_2
XFILLER_190_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_63_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_729 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_216 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_32_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__091__A vssd2 vccd1 vccd1 vssd2 _351_/Q sky130_fd_sc_hd__diode_2
XFILLER_136_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__086__B1 vssd2 vccd1 vccd1 vssd2 _345_/Q sky130_fd_sc_hd__diode_2
XFILLER_232_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_48_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input130_A vssd2 vccd1 vccd1 vssd2 la_data_in[67] sky130_fd_sc_hd__diode_2
XFILLER_169_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input228_A vssd2 vccd1 vccd1 vssd2 la_oenb[3] sky130_fd_sc_hd__diode_2
XFILLER_100_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_76 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_324_ vssd2 _324_/X vccd1 _326_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_243_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_255_ _255_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_186_ _186_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_443 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_48_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_111_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__077__B1 vssd2 vccd1 vccd1 vssd2 _348_/Q sky130_fd_sc_hd__diode_2
XFILLER_96_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_2342 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__092__A3 vssd2 vccd1 vccd1 vssd2 _352_/Q sky130_fd_sc_hd__diode_2
XFILLER_231_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1359 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_659 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_228_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_160 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA__083__A3 vssd2 vccd1 vccd1 vssd2 _355_/Q sky130_fd_sc_hd__diode_2
XFILLER_84_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1871 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_515 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_245_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_180_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_559 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_36_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1760 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_166_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input178_A vssd2 vccd1 vccd1 vssd2 la_oenb[10] sky130_fd_sc_hd__diode_2
XFILLER_4_969 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input345_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[23] sky130_fd_sc_hd__diode_2
XFILLER_78_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_121_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__059__B1 vssd2 vccd1 vccd1 vssd2 _354_/Q sky130_fd_sc_hd__diode_2
XFILLER_94_707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input39_A vssd2 vccd1 vccd1 vssd2 la_data_in[0] sky130_fd_sc_hd__diode_2
XFILLER_219_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_187_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
X_307_ _307_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_147_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_238_ _238_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_183_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_169_ _169_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_109_680 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1313 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_161_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_416 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_103_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput306 vssd2 input306/X vccd1 wbs_adr_i[18] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput317 vssd2 input317/X vccd1 wbs_adr_i[28] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_46 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput328 vssd2 input328/X vccd1 wbs_adr_i[9] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_29_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput339 vssd2 input339/X vccd1 wbs_dat_i[18] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_5_1235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_229_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_246_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_80_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_378 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input295_A vssd2 vccd1 vccd1 vssd2 user_clock2 sky130_fd_sc_hd__diode_2
XFILLER_8_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1888 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_871 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_187_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2059 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_66_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_187_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__357__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_172_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput103 vssd2 input103/X vccd1 la_data_in[42] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_235_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput114 vssd2 input114/X vccd1 la_data_in[52] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput125 vssd2 input125/X vccd1 la_data_in[62] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput136 vssd2 input136/X vccd1 la_data_in[72] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput147 vssd2 input147/X vccd1 la_data_in[82] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput158 vssd2 input158/X vccd1 la_data_in[92] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput169 vssd2 input169/X vccd1 la_oenb[101] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1927 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_5_1098 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input210_A vssd2 vccd1 vccd1 vssd2 la_oenb[23] sky130_fd_sc_hd__diode_2
XFILLER_44_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input308_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[1] sky130_fd_sc_hd__diode_2
XFILLER_71_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_131 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_246_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_142 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_188_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_186 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_140_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_386 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_846 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_2197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_0 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_108_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_1155 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_213_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_26_456 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_166_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_235_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input160_A vssd2 vccd1 vccd1 vssd2 la_data_in[94] sky130_fd_sc_hd__diode_2
XFILLER_122_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_89_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input258_A vssd2 vccd1 vccd1 vssd2 la_oenb[67] sky130_fd_sc_hd__diode_2
XFILLER_122_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input21_A vssd2 vccd1 vccd1 vssd2 io_in[28] sky130_fd_sc_hd__diode_2
XFILLER_188_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1724 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput407 vssd2 io_out[10] vccd1 _127_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput418 vssd2 io_out[20] vccd1 _137_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput429 vssd2 io_out[30] vccd1 _342_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_110_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_3_1514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_82_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1558 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_210_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_340_ _098_/X _340_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _340_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_243_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_45 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_271_ _271_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_52_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_204_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input69_A vssd2 vccd1 vccd1 vssd2 la_data_in[127] sky130_fd_sc_hd__diode_2
XFILLER_162_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2200 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1521 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2212 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_220_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__095__A1 vssd2 vccd1 vccd1 vssd2 _075_/A sky130_fd_sc_hd__diode_2
XFILLER_231_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_2056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__086__A1 vssd2 vccd1 vccd1 vssd2 _099_/A sky130_fd_sc_hd__diode_2
XFILLER_150_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input123_A vssd2 vccd1 vccd1 vssd2 la_data_in[60] sky130_fd_sc_hd__diode_2
XFILLER_62_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_323_ vssd2 _323_/X vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_254_ _254_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_243_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_411 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_185_ _185_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_87_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_136_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_383 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_375 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_96_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__077__A1 vssd2 vccd1 vccd1 vssd2 _099_/A sky130_fd_sc_hd__diode_2
XFILLER_215_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_237_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_153_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_52_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1772 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput590 vssd2 wbs_dat_o[22] vccd1 _298_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__059__A1 vssd2 vccd1 vccd1 vssd2 _355_/Q sky130_fd_sc_hd__diode_2
XANTENNA__059__B2 vssd2 vccd1 vccd1 vssd2 _056_/X sky130_fd_sc_hd__diode_2
XANTENNA_input240_A vssd2 vccd1 vccd1 vssd2 la_oenb[50] sky130_fd_sc_hd__diode_2
XFILLER_121_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input338_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[17] sky130_fd_sc_hd__diode_2
XFILLER_47_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_306_ _306_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_15_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_237_ _237_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_15_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_168_ _168_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_217_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_099_ vssd2 _338_/A vccd1 _099_/A vccd1 _099_/B vssd2 sky130_fd_sc_hd__nor2_4
XFILLER_108_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_78_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_81_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2059 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_439 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_216_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput307 vssd2 input307/X vccd1 wbs_adr_i[19] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput318 vssd2 input318/X vccd1 wbs_adr_i[29] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_233_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput329 vssd2 input329/X vccd1 wbs_cyc_i vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_60_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__097__A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_244_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_302 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_313 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_52_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_357 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_101_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input190_A vssd2 vccd1 vccd1 vssd2 la_oenb[120] sky130_fd_sc_hd__diode_2
XFILLER_201_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input288_A vssd2 vccd1 vccd1 vssd2 la_oenb[94] sky130_fd_sc_hd__diode_2
XFILLER_101_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input51_A vssd2 vccd1 vccd1 vssd2 la_data_in[110] sky130_fd_sc_hd__diode_2
XFILLER_10_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2313 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1667 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_891 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_37 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
Xinput104 vssd2 input104/X vccd1 la_data_in[43] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_163_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput115 vssd2 input115/X vccd1 la_data_in[53] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
Xinput126 vssd2 input126/X vccd1 la_data_in[63] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
Xinput137 vssd2 input137/X vccd1 la_data_in[73] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput148 vssd2 input148/X vccd1 la_data_in[83] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput159 vssd2 input159/X vccd1 la_data_in[93] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_233_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input203_A vssd2 vccd1 vccd1 vssd2 la_oenb[17] sky130_fd_sc_hd__diode_2
XFILLER_147_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_143 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input99_A vssd2 vccd1 vccd1 vssd2 la_data_in[39] sky130_fd_sc_hd__diode_2
XPHY_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_680 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_2132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_35_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_147_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1464 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_1 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_63_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_108_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_176_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_22_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_390 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_468 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_194_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_89_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input153_A vssd2 vccd1 vccd1 vssd2 la_data_in[88] sky130_fd_sc_hd__diode_2
XFILLER_150_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_578 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_89_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input320_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[30] sky130_fd_sc_hd__diode_2
XFILLER_190_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input14_A vssd2 vccd1 vccd1 vssd2 io_in[21] sky130_fd_sc_hd__diode_2
XFILLER_248_1736 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_1379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput408 vssd2 io_out[11] vccd1 _128_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput419 vssd2 io_out[21] vccd1 _138_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2216 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1261 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_184_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__347__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_50_257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_204_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input6_A vssd2 vccd1 vccd1 vssd2 io_in[14] sky130_fd_sc_hd__diode_2
XFILLER_59_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_219_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_74_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_37_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_900 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_270_ _270_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_243_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input270_A vssd2 vccd1 vccd1 vssd2 la_oenb[78] sky130_fd_sc_hd__diode_2
XFILLER_13_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1509 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1533 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_233_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_141_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__095__A2 vssd2 vccd1 vccd1 vssd2 _076_/A sky130_fd_sc_hd__diode_2
XFILLER_229_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_225_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_144_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__086__A2 vssd2 vccd1 vccd1 vssd2 _099_/B sky130_fd_sc_hd__diode_2
XFILLER_210_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_406 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_74_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input116_A vssd2 vccd1 vccd1 vssd2 la_data_in[54] sky130_fd_sc_hd__diode_2
XFILLER_161_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_322_ vssd2 _322_/X vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_187_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
X_253_ _253_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input81_A vssd2 vccd1 vccd1 vssd2 la_data_in[22] sky130_fd_sc_hd__diode_2
XFILLER_80_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_184_ _184_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_183_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1009 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_123_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_151_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_673 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_123_387 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_78_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__077__A2 vssd2 vccd1 vccd1 vssd2 _099_/B sky130_fd_sc_hd__diode_2
XFILLER_96_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_111_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1330 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_146_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2090 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_94_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_186_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_56_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1142 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_517 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_109_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_105_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput580 vssd2 wbs_dat_o[13] vccd1 _289_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput591 vssd2 wbs_dat_o[23] vccd1 _299_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_82_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__059__A2 vssd2 vccd1 vccd1 vssd2 _055_/X sky130_fd_sc_hd__diode_2
XFILLER_169_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_210_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input233_A vssd2 vccd1 vccd1 vssd2 la_oenb[44] sky130_fd_sc_hd__diode_2
XFILLER_169_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1952 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_47_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1827 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_305_ _305_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_230_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_236_ _236_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_167_ _167_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_155_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_098_ vssd2 _098_/X vccd1 _105_/A vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_108_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_41 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_93_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1103 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_2038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput308 vssd2 input308/X vccd1 wbs_adr_i[1] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_29_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
Xinput319 vssd2 input319/X vccd1 wbs_adr_i[2] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_233_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_68_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_56_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_246_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_314 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_101_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input183_A vssd2 vccd1 vccd1 vssd2 la_oenb[114] sky130_fd_sc_hd__diode_2
XFILLER_177_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input350_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[28] sky130_fd_sc_hd__diode_2
XFILLER_79_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input44_A vssd2 vccd1 vccd1 vssd2 la_data_in[104] sky130_fd_sc_hd__diode_2
XFILLER_133_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_86_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_19_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1602 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1782 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_63_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_204_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_870 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_32_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_390 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_219_ _219_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_237_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_57_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_49 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput105 vssd2 input105/X vccd1 la_data_in[44] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_130_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput116 vssd2 input116/X vccd1 la_data_in[54] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
Xinput127 vssd2 input127/X vccd1 la_data_in[64] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_170_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput138 vssd2 input138/X vccd1 la_data_in[74] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_29_411 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput149 vssd2 input149/X vccd1 la_data_in[84] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_243_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1078 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_29_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1988 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_155 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_40_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_692 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_2 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_245_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_176_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_176_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_28_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1102 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_27_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_208_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_239_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input146_A vssd2 vccd1 vccd1 vssd2 la_data_in[81] sky130_fd_sc_hd__diode_2
XFILLER_130_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_218_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input313_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[24] sky130_fd_sc_hd__diode_2
XFILLER_85_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_60 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1473 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput409 vssd2 io_out[12] vccd1 _129_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_94_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_58_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_82_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_225_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_176_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_195_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1059 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_57_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_912 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_108_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input263_A vssd2 vccd1 vccd1 vssd2 la_oenb[71] sky130_fd_sc_hd__diode_2
XFILLER_137_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__089__B1 vssd2 vccd1 vccd1 vssd2 _344_/Q sky130_fd_sc_hd__diode_2
XFILLER_172_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_45_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_57_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__095__A3 vssd2 vccd1 vccd1 vssd2 _351_/Q sky130_fd_sc_hd__diode_2
XFILLER_122_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_133_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_60 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__086__A3 vssd2 vccd1 vccd1 vssd2 _354_/Q sky130_fd_sc_hd__diode_2
XFILLER_86_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_58_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_230_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input109_A vssd2 vccd1 vccd1 vssd2 la_data_in[48] sky130_fd_sc_hd__diode_2
XFILLER_120_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_321_ vssd2 _321_/X vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_230_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_252_ _252_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_17_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_183_ _183_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input74_A vssd2 vccd1 vccd1 vssd2 la_data_in[16] sky130_fd_sc_hd__diode_2
XFILLER_155_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__077__A3 vssd2 vccd1 vccd1 vssd2 _357_/Q sky130_fd_sc_hd__diode_2
XFILLER_78_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_150_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1318 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_31_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_119_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_529 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_137_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_427 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_105_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput570 vssd2 la_data_out[99] vccd1 _243_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput581 vssd2 wbs_dat_o[14] vccd1 _290_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1021 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput592 vssd2 wbs_dat_o[24] vccd1 _300_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input226_A vssd2 vccd1 vccd1 vssd2 la_oenb[38] sky130_fd_sc_hd__diode_2
XFILLER_86_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_304_ _304_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_30_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_235_ _235_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_129_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_166_ _166_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_097_ vssd2 _105_/A vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_170_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_460 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_238_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_81_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_130_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput309 vssd2 input309/X vccd1 wbs_adr_i[20] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_170_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_9_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_83_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_216_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_326 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_359 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_119_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input176_A vssd2 vccd1 vccd1 vssd2 la_oenb[108] sky130_fd_sc_hd__diode_2
XFILLER_238_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input343_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[21] sky130_fd_sc_hd__diode_2
XFILLER_105_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input37_A vssd2 vccd1 vccd1 vssd2 io_in[8] sky130_fd_sc_hd__diode_2
XFILLER_216_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_86_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_896 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_871 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_218_ _218_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_129_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_149_ _149_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_201_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_repeater608_A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_10_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1102 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_0_1179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput106 vssd2 input106/X vccd1 la_data_in[45] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_102_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput117 vssd2 input117/X vccd1 la_data_in[55] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_130_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput128 vssd2 input128/X vccd1 la_data_in[65] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput139 vssd2 input139/X vccd1 la_data_in[75] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_130_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1901 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_22_1851 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1945 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_53_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_198_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_181_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input293_A vssd2 vccd1 vccd1 vssd2 la_oenb[99] sky130_fd_sc_hd__diode_2
XFILLER_166_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_188_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_90_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_212 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_75_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_407 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_17_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_19_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_191_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_15_1176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1114 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_238_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_165_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_941 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_133_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_235_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input139_A vssd2 vccd1 vccd1 vssd2 la_data_in[75] sky130_fd_sc_hd__diode_2
XFILLER_22_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_57_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1720 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_72_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_245_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input306_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[18] sky130_fd_sc_hd__diode_2
XFILLER_72_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1786 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_9_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1485 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_138_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_48_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_204 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_119_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_924 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_180_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__089__A1 vssd2 vccd1 vccd1 vssd2 _075_/A sky130_fd_sc_hd__diode_2
XFILLER_151_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input256_A vssd2 vccd1 vccd1 vssd2 la_oenb[65] sky130_fd_sc_hd__diode_2
XFILLER_172_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1502 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_94_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_100_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_92 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_145_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_145_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_320_ vssd2 _320_/X vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_204_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_251_ _251_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_167_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_182_ _182_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_127_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_155_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input67_A vssd2 vccd1 vccd1 vssd2 la_data_in[125] sky130_fd_sc_hd__diode_2
XFILLER_191_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_631 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_123_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_151_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_402 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_20_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__100__A vssd2 vccd1 vccd1 vssd2 _351_/Q sky130_fd_sc_hd__diode_2
XFILLER_248_2055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_671 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_981 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_142 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_190_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_170_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1886 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XPHY_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_127_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_30_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_406 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_180_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_47_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput560 vssd2 la_data_out[8] vccd1 _152_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xoutput571 vssd2 la_data_out[9] vccd1 _153_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput582 vssd2 wbs_dat_o[15] vccd1 _291_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_120_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput593 vssd2 wbs_dat_o[25] vccd1 _301_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_182_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1033 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input121_A vssd2 vccd1 vccd1 vssd2 la_data_in[59] sky130_fd_sc_hd__diode_2
XFILLER_216_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input219_A vssd2 vccd1 vccd1 vssd2 la_oenb[31] sky130_fd_sc_hd__diode_2
XFILLER_234_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_303_ _303_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_223_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_234_ _234_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_221_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_165_ _165_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_109_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_096_ vssd2 _342_/D _074_/A _095_/X vccd1 _100_/B _339_/X _104_/A vccd1 vssd2 sky130_fd_sc_hd__o311a_1
XFILLER_170_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_984 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_472 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_69_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_65 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_65_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_243 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_53_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1173 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_119_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_220_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_130_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_774 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_240_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input169_A vssd2 vccd1 vccd1 vssd2 la_oenb[101] sky130_fd_sc_hd__diode_2
XFILLER_126_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput390 vssd2 io_oeb[2] vccd1 _109_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_842 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input336_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[15] sky130_fd_sc_hd__diode_2
XFILLER_120_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_235_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_1762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_850 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_872 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_883 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_128_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_217_ _217_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_156_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_148_ _148_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_116_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_079_ vssd2 _079_/Y vccd1 _355_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_217_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_187_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_162_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput107 vssd2 input107/X vccd1 la_data_in[46] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput118 vssd2 input118/X vccd1 la_data_in[56] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_102_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput129 vssd2 input129/X vccd1 la_data_in[66] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_69_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_102 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_112_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_53_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_138_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input286_A vssd2 vccd1 vccd1 vssd2 la_oenb[92] sky130_fd_sc_hd__diode_2
XFILLER_181_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_5_1570 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_147_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_4 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_147_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_419 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_231_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_680 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_195_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_171_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_953 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_195_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_174_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_515 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_27_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_559 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input201_A vssd2 vccd1 vccd1 vssd2 la_oenb[15] sky130_fd_sc_hd__diode_2
XFILLER_32_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input97_A vssd2 vccd1 vccd1 vssd2 la_data_in[37] sky130_fd_sc_hd__diode_2
XFILLER_16_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_201_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_141_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_94_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_500 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_48_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_216 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_32_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_227_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_180_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_958 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__089__A2 vssd2 vccd1 vccd1 vssd2 _076_/A sky130_fd_sc_hd__diode_2
XFILLER_235_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input151_A vssd2 vccd1 vccd1 vssd2 la_data_in[86] sky130_fd_sc_hd__diode_2
XFILLER_231_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input249_A vssd2 vccd1 vccd1 vssd2 la_oenb[59] sky130_fd_sc_hd__diode_2
XFILLER_131_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input12_A vssd2 vccd1 vccd1 vssd2 io_in[1] sky130_fd_sc_hd__diode_2
XFILLER_217_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_232_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_96_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_159_60 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_155_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_673 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_175_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput290 vssd2 input290/X vccd1 la_oenb[96] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1359 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_51_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_36_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input4_A vssd2 vccd1 vccd1 vssd2 io_in[12] sky130_fd_sc_hd__diode_2
XFILLER_101_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_58_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_250_ _250_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_120_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_181_ _181_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_210_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input199_A vssd2 vccd1 vccd1 vssd2 la_oenb[13] sky130_fd_sc_hd__diode_2
XFILLER_182_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input366_A vssd2 vccd1 vccd1 vssd2 wbs_stb_i sky130_fd_sc_hd__diode_2
XFILLER_135_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_414 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__100__B vssd2 vccd1 vccd1 vssd2 _100_/B sky130_fd_sc_hd__diode_2
XFILLER_234_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1388 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_115_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_83_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_221_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_227_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_509 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput550 vssd2 la_data_out[80] vccd1 _224_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput561 vssd2 la_data_out[90] vccd1 _234_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput572 vssd2 user_irq[0] vccd1 _272_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_216_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_59_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput583 vssd2 wbs_dat_o[16] vccd1 _292_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput594 vssd2 wbs_dat_o[26] vccd1 _302_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1900 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_1999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input114_A vssd2 vccd1 vccd1 vssd2 la_data_in[52] sky130_fd_sc_hd__diode_2
XFILLER_93_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_302_ _302_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_19_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_233_ _233_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_15_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_156_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_164_ _164_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_095_ vssd2 _095_/X _342_/Q vccd1 _075_/A _076_/A _351_/Q vccd1 vssd2 sky130_fd_sc_hd__a31o_1
XFILLER_124_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_440 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_9_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_786 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_10_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput380 vssd2 io_oeb[20] vccd1 _318_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput391 vssd2 io_oeb[30] vccd1 _328_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_160_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input231_A vssd2 vccd1 vccd1 vssd2 la_oenb[42] sky130_fd_sc_hd__diode_2
XFILLER_21_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_87_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input329_A vssd2 vccd1 vccd1 vssd2 wbs_cyc_i sky130_fd_sc_hd__diode_2
XFILLER_142_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1774 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_406 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_90_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_210_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__070__B1 vssd2 vccd1 vccd1 vssd2 _069_/Y sky130_fd_sc_hd__diode_2
XFILLER_182_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_851 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_862 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_884 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_895 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_216_ _216_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_147_ _147_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_184_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_078_ vssd2 _348_/D _074_/X _077_/X vccd1 _071_/Y _104_/A _073_/X vccd1 vssd2 sky130_fd_sc_hd__o311a_1
XFILLER_217_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__061__B1 vssd2 vccd1 vccd1 vssd2 _352_/Q sky130_fd_sc_hd__diode_2
XFILLER_221_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput108 vssd2 input108/X vccd1 la_data_in[47] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_9_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput119 vssd2 input119/X vccd1 la_data_in[57] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_213_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_5_1004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_57_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2171 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_186_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_103 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_114 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_112_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_686 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_205_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_147 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input181_A vssd2 vccd1 vccd1 vssd2 la_oenb[112] sky130_fd_sc_hd__diode_2
XFILLER_153_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input279_A vssd2 vccd1 vccd1 vssd2 la_oenb[86] sky130_fd_sc_hd__diode_2
XFILLER_193_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input42_A vssd2 vccd1 vccd1 vssd2 la_data_in[102] sky130_fd_sc_hd__diode_2
XFILLER_212_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_248_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_2283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_130_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_28_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_210_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_5 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_175_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_692 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_50_1036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_30_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_repeater613_A vssd2 vccd1 vccd1 vssd2 input16/X sky130_fd_sc_hd__diode_2
XFILLER_176_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2357 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_135_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput90 vssd2 input90/X vccd1 la_data_in[30] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_123_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_131_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_177_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_1232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_177_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_58_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_187_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1029 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_66_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_120_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__089__A3 vssd2 vccd1 vccd1 vssd2 _353_/Q sky130_fd_sc_hd__diode_2
XFILLER_116_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input144_A vssd2 vccd1 vccd1 vssd2 la_data_in[7] sky130_fd_sc_hd__diode_2
XFILLER_58_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_248_2216 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_2170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_91_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input311_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[22] sky130_fd_sc_hd__diode_2
XFILLER_185_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_91_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_232_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1103 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_173 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_116_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_2006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_228_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput280 vssd2 input280/X vccd1 la_oenb[87] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_184_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput291 vssd2 input291/X vccd1 la_oenb[97] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_180_ _180_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_10_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_167_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input261_A vssd2 vccd1 vccd1 vssd2 la_oenb[6] sky130_fd_sc_hd__diode_2
XFILLER_150_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input359_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[7] sky130_fd_sc_hd__diode_2
XFILLER_215_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_143 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_238_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2002 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_248_1301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_234_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_234_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_142_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_460 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_55_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_815 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput540 vssd2 la_data_out[71] vccd1 _215_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput551 vssd2 la_data_out[81] vccd1 _225_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput562 vssd2 la_data_out[91] vccd1 _235_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput573 vssd2 user_irq[1] vccd1 _273_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1002 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xoutput584 vssd2 wbs_dat_o[17] vccd1 _293_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_232_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput595 vssd2 wbs_dat_o[27] vccd1 _303_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1912 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_515 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_145_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input107_A vssd2 vccd1 vccd1 vssd2 la_data_in[46] sky130_fd_sc_hd__diode_2
XFILLER_106_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_301_ _301_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_24_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_232_ _232_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_163_ _163_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_210_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input72_A vssd2 vccd1 vccd1 vssd2 la_data_in[14] sky130_fd_sc_hd__diode_2
X_094_ vssd2 _100_/B vccd1 _350_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_30_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_34 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2009 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__350__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_225_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_11_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_318 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput370 vssd2 io_oeb[11] vccd1 _312_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput381 vssd2 io_oeb[21] vccd1 _319_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput392 vssd2 io_oeb[31] vccd1 _329_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_248_822 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_888 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input224_A vssd2 vccd1 vccd1 vssd2 la_oenb[36] sky130_fd_sc_hd__diode_2
XFILLER_19_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_62_418 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__070__A1 vssd2 vccd1 vccd1 vssd2 _349_/Q sky130_fd_sc_hd__diode_2
XFILLER_37_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_35_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_245_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_830 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_863 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_204_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_874 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_896 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_204_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_215_ _215_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_146_ _146_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_077_ vssd2 _077_/X _348_/Q vccd1 _099_/A _099_/B _357_/Q vccd1 vssd2 sky130_fd_sc_hd__a31o_1
XFILLER_124_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_692 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__061__A1 vssd2 vccd1 vccd1 vssd2 _353_/Q sky130_fd_sc_hd__diode_2
XFILLER_37_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__061__B2 vssd2 vccd1 vccd1 vssd2 _056_/X sky130_fd_sc_hd__diode_2
XFILLER_76_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_83_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput109 vssd2 input109/X vccd1 la_data_in[48] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_129 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1810 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_65_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_209_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_80_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_241_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_159 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input174_A vssd2 vccd1 vccd1 vssd2 la_oenb[106] sky130_fd_sc_hd__diode_2
XFILLER_106_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input341_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[1] sky130_fd_sc_hd__diode_2
XFILLER_23_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input35_A vssd2 vccd1 vccd1 vssd2 io_in[6] sky130_fd_sc_hd__diode_2
XFILLER_5_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_521 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_2104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_2295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_247_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_660 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_671 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_31_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_178_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_129_ _129_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_176_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_900 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1945 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput80 vssd2 input80/X vccd1 la_data_in[21] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_163_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput91 vssd2 input91/X vccd1 la_data_in[31] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_66_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1712 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_83_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_197_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input291_A vssd2 vccd1 vccd1 vssd2 la_oenb[97] sky130_fd_sc_hd__diode_2
XFILLER_220_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_106_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_34_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_195_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__310__A vssd2 vccd1 vccd1 vssd2 _316_/A sky130_fd_sc_hd__diode_2
XFILLER_39_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_671 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_81_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_175_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_200_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_150_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_2228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input137_A vssd2 vccd1 vccd1 vssd2 la_data_in[73] sky130_fd_sc_hd__diode_2
XFILLER_58_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2243 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input304_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[16] sky130_fd_sc_hd__diode_2
XFILLER_2_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_232_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_159_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_159_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_114_518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_218_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput270 vssd2 input270/X vccd1 la_oenb[78] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput281 vssd2 input281/X vccd1 la_oenb[88] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_3_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput292 vssd2 input292/X vccd1 la_oenb[98] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_162_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_87_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_178_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_109_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_623 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input254_A vssd2 vccd1 vccd1 vssd2 la_oenb[63] sky130_fd_sc_hd__diode_2
XFILLER_150_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_8_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_58_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_166_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_472 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_175_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
Xoutput530 vssd2 la_data_out[62] vccd1 _206_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput541 vssd2 la_data_out[72] vccd1 _216_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput552 vssd2 la_data_out[82] vccd1 _226_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput563 vssd2 la_data_out[92] vccd1 _236_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput574 vssd2 user_irq[2] vccd1 _274_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput585 vssd2 wbs_dat_o[18] vccd1 _294_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput596 vssd2 wbs_dat_o[28] vccd1 _304_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_232_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_228_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_228_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_210_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_300_ _300_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_106_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_231_ _231_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_50_390 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_896 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
X_162_ _162_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_093_ vssd2 _343_/D _074_/A _092_/X vccd1 _091_/Y _072_/A _339_/X vccd1 vssd2 sky130_fd_sc_hd__o311a_1
XFILLER_174_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input65_A vssd2 vccd1 vccd1 vssd2 la_data_in[123] sky130_fd_sc_hd__diode_2
XFILLER_124_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_120_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_45_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_73_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput1 vssd2 input1/X vccd1 io_in[0] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_232_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_45_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_80_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_101_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_138_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput371 vssd2 io_oeb[12] vccd1 _313_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput382 vssd2 io_oeb[22] vccd1 _320_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput393 vssd2 io_oeb[32] vccd1 _330_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_834 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_126_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_5_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_59_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input217_A vssd2 vccd1 vccd1 vssd2 la_oenb[2] sky130_fd_sc_hd__diode_2
XFILLER_243_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_55_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__070__A2 vssd2 vccd1 vccd1 vssd2 _066_/X sky130_fd_sc_hd__diode_2
XFILLER_27_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_19_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_187_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_831 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_842 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_875 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_886 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_214_ _214_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XPHY_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_373 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_204_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_145_ _145_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_167_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_7_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_076_ vssd2 _099_/B vccd1 _076_/A vccd1 vssd2 sky130_fd_sc_hd__buf_4
XFILLER_136_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output436_A vssd2 vccd1 vccd1 vssd2 _349_/Q sky130_fd_sc_hd__diode_2
XFILLER_234_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_228_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__061__A2 vssd2 vccd1 vccd1 vssd2 _055_/A sky130_fd_sc_hd__diode_2
XFILLER_37_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_186_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__313__A vssd2 vccd1 vccd1 vssd2 _316_/A sky130_fd_sc_hd__diode_2
XFILLER_235_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_135_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1028 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1822 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1916 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_44_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_2341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_112_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_116 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_0_1673 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_80_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__340__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_181_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input167_A vssd2 vccd1 vccd1 vssd2 la_oenb[0] sky130_fd_sc_hd__diode_2
XFILLER_97_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input334_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[13] sky130_fd_sc_hd__diode_2
XFILLER_102_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input28_A vssd2 vccd1 vccd1 vssd2 io_in[34] sky130_fd_sc_hd__diode_2
XFILLER_247_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_31_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_672 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_1016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_128_ _128_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_176_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_197_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_059_ vssd2 _354_/D _354_/Q vccd1 _056_/X _355_/Q _055_/X vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_171_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_818 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_912 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__308__A vssd2 vccd1 vccd1 vssd2 _316_/A sky130_fd_sc_hd__diode_2
XFILLER_210_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1957 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput70 vssd2 input70/X vccd1 la_data_in[12] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_200_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput81 vssd2 input81/X vccd1 la_data_in[22] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_172_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput92 vssd2 input92/X vccd1 la_data_in[32] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_239_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_235_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_232_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1757 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1401 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input284_A vssd2 vccd1 vccd1 vssd2 la_oenb[90] sky130_fd_sc_hd__diode_2
XFILLER_165_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_121_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_57_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_189_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_12_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_113_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_65 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_411 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_150_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_183_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input95_A vssd2 vccd1 vccd1 vssd2 la_data_in[35] sky130_fd_sc_hd__diode_2
XFILLER_13_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_99_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput260 vssd2 input260/X vccd1 la_oenb[69] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_236_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput271 vssd2 input271/X vccd1 la_oenb[79] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput282 vssd2 input282/X vccd1 la_oenb[89] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_236_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput293 vssd2 input293/X vccd1 la_oenb[99] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_63_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_162_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1086 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_162_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__321__A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_59_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_602 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_117_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_145_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input247_A vssd2 vccd1 vccd1 vssd2 la_oenb[57] sky130_fd_sc_hd__diode_2
XFILLER_49_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input10_A vssd2 vccd1 vccd1 vssd2 io_in[18] sky130_fd_sc_hd__diode_2
XFILLER_246_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_182_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_484 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_69_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_127_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_63_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_211_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__316__A vssd2 vccd1 vccd1 vssd2 _316_/A sky130_fd_sc_hd__diode_2
XFILLER_242_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput520 vssd2 la_data_out[53] vccd1 _197_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_172_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput531 vssd2 la_data_out[63] vccd1 _207_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput542 vssd2 la_data_out[73] vccd1 _217_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput553 vssd2 la_data_out[83] vccd1 _227_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput564 vssd2 la_data_out[93] vccd1 _237_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput575 vssd2 wbs_ack_o vccd1 _275_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_232_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput586 vssd2 wbs_dat_o[19] vccd1 _295_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput597 vssd2 wbs_dat_o[29] vccd1 _305_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input2_A vssd2 vccd1 vccd1 vssd2 io_in[10] sky130_fd_sc_hd__diode_2
XFILLER_214_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_186_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_180_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_230_ _230_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_243_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_161_ _161_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input197_A vssd2 vccd1 vccd1 vssd2 la_oenb[127] sky130_fd_sc_hd__diode_2
XFILLER_221_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_092_ vssd2 _092_/X _343_/Q vccd1 _075_/A _076_/A _352_/Q vccd1 vssd2 sky130_fd_sc_hd__a31o_1
XFILLER_171_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input364_A vssd2 vccd1 vccd1 vssd2 wbs_sel_i[2] sky130_fd_sc_hd__diode_2
XFILLER_124_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_2315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input58_A vssd2 vccd1 vccd1 vssd2 la_data_in[117] sky130_fd_sc_hd__diode_2
XFILLER_124_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_977 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_172_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_14 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_46_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_185_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output583_A vssd2 vccd1 vccd1 vssd2 _292_/LO sky130_fd_sc_hd__diode_2
XFILLER_204_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput2 vssd2 input2/X vccd1 io_in[10] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_168_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_110_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_146_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_195_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput372 vssd2 io_oeb[13] vccd1 _114_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput383 vssd2 io_oeb[23] vccd1 _321_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_813 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xoutput394 vssd2 io_oeb[33] vccd1 _331_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_28_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input112_A vssd2 vccd1 vccd1 vssd2 la_data_in[50] sky130_fd_sc_hd__diode_2
XFILLER_243_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_810 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_215_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_843 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_145_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_180_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_213_ _213_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XPHY_887 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_144_ _144_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_075_ vssd2 _099_/A vccd1 _075_/A vccd1 vssd2 sky130_fd_sc_hd__buf_4
XFILLER_100_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_215_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_output429_A vssd2 vccd1 vccd1 vssd2 _342_/Q sky130_fd_sc_hd__diode_2
XFILLER_215_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_672 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_187_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_128_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_179_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_590 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_143_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_80_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_700 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_106_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_610 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input327_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[8] sky130_fd_sc_hd__diode_2
XFILLER_75_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_46_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_8 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_189_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_673 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_684 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_1028 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_127_ _127_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_183_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_058_ vssd2 _355_/D _355_/Q vccd1 _056_/X _356_/Q _055_/X vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_113_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_375 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_81_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1972 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_146_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_924 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_228_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1969 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_147_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__324__A vssd2 vccd1 vccd1 vssd2 _326_/A sky130_fd_sc_hd__diode_2
XFILLER_190_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput60 vssd2 input60/X vccd1 la_data_in[119] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput71 vssd2 input71/X vccd1 la_data_in[13] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_200_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput82 vssd2 input82/X vccd1 la_data_in[23] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_128_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput93 vssd2 input93/X vccd1 la_data_in[33] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_239_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_66_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_107_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_153_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input277_A vssd2 vccd1 vccd1 vssd2 la_oenb[84] sky130_fd_sc_hd__diode_2
XFILLER_165_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input40_A vssd2 vccd1 vccd1 vssd2 la_data_in[100] sky130_fd_sc_hd__diode_2
XFILLER_27_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_103_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_180_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_208_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_125_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_157_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_repeater611_A vssd2 vccd1 vccd1 vssd2 _335_/A sky130_fd_sc_hd__diode_2
XFILLER_12_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_342 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__319__A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_187_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_77 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_929 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__054__A vssd2 vccd1 vccd1 vssd2 _065_/A sky130_fd_sc_hd__diode_2
XFILLER_147_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_416 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_159_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_199_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input88_A vssd2 vccd1 vccd1 vssd2 la_data_in[29] sky130_fd_sc_hd__diode_2
XFILLER_182_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_655 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_142_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_688 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_190_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_150_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_110_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__353__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_95_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput250 vssd2 input250/X vccd1 la_oenb[5] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput261 vssd2 input261/X vccd1 la_oenb[6] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput272 vssd2 input272/X vccd1 la_oenb[7] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_231_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput283 vssd2 input283/X vccd1 la_oenb[8] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput294 vssd2 input294/X vccd1 la_oenb[9] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_236_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1021 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_225_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_129_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_89_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input142_A vssd2 vccd1 vccd1 vssd2 la_data_in[78] sky130_fd_sc_hd__diode_2
XFILLER_237_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_54_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_496 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2171 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_32_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__332__A vssd2 vccd1 vccd1 vssd2 _335_/A sky130_fd_sc_hd__diode_2
Xoutput510 vssd2 la_data_out[44] vccd1 _188_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput521 vssd2 la_data_out[54] vccd1 _198_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput532 vssd2 la_data_out[64] vccd1 _208_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_246_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput543 vssd2 la_data_out[74] vccd1 _218_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput554 vssd2 la_data_out[84] vccd1 _228_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput565 vssd2 la_data_out[94] vccd1 _238_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput576 vssd2 wbs_dat_o[0] vccd1 _276_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput587 vssd2 wbs_dat_o[1] vccd1 _277_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput598 vssd2 wbs_dat_o[2] vccd1 _278_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_243_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2072 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_160_ _160_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_24_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_091_ vssd2 _091_/Y vccd1 _351_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_108_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_151_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input357_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[5] sky130_fd_sc_hd__diode_2
XFILLER_215_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_8_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_26 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_232_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_185_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_289_ _289_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput3 vssd2 input3/X vccd1 io_in[11] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_77_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__327__A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_221_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput373 vssd2 io_oeb[14] vccd1 _115_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput384 vssd2 io_oeb[24] vccd1 _322_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput395 vssd2 io_oeb[34] vccd1 _332_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_3_2170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_800 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input105_A vssd2 vccd1 vccd1 vssd2 la_data_in[44] sky130_fd_sc_hd__diode_2
XFILLER_163_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_215_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_822 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_43_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_844 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_855 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_212_ _212_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XPHY_877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_888 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_11_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_899 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_143_ _143_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_183_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input70_A vssd2 vccd1 vccd1 vssd2 la_data_in[12] sky130_fd_sc_hd__diode_2
X_074_ vssd2 _074_/X vccd1 _074_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_4
XFILLER_125_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_136_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_124_478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_111_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2142 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_246_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_55_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_52_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_129 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_224_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_546 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input222_A vssd2 vccd1 vccd1 vssd2 la_oenb[34] sky130_fd_sc_hd__diode_2
XFILLER_186_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1406 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_112_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1428 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_9 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_178_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_696 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_36 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_126_ _126_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_193_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
X_057_ vssd2 _356_/D _356_/Q vccd1 _056_/X _357_/Q _055_/X vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_178_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_206_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_958 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput50 vssd2 input50/X vccd1 la_data_in[10] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_162_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput61 vssd2 input61/X vccd1 la_data_in[11] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput72 vssd2 input72/X vccd1 la_data_in[14] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_238_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput83 vssd2 input83/X vccd1 la_data_in[24] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput94 vssd2 input94/X vccd1 la_data_in[34] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_115_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_37 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_218_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_183_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input172_A vssd2 vccd1 vccd1 vssd2 la_oenb[104] sky130_fd_sc_hd__diode_2
XFILLER_194_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_7_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_164_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_164_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input33_A vssd2 vccd1 vccd1 vssd2 io_in[4] sky130_fd_sc_hd__diode_2
XFILLER_212_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_75_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_1350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_186_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_73_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_71_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_460 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_176_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_193_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_109_ _109_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_172_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__335__A vssd2 vccd1 vccd1 vssd2 _335_/A sky130_fd_sc_hd__diode_2
XFILLER_17_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1501 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_6_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_233_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_428 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput240 vssd2 input240/X vccd1 la_oenb[50] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput251 vssd2 input251/X vccd1 la_oenb[60] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput262 vssd2 input262/X vccd1 la_oenb[70] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput273 vssd2 input273/X vccd1 la_oenb[80] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_208_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput284 vssd2 input284/X vccd1 la_oenb[90] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_36_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput295 vssd2 input295/X vccd1 user_clock2 vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1000 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1066 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_204_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_973 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__065__A vssd2 vccd1 vccd1 vssd2 _065_/A sky130_fd_sc_hd__diode_2
XFILLER_225_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_108_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_215_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_659 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_132_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_427 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_24_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input135_A vssd2 vccd1 vccd1 vssd2 la_data_in[71] sky130_fd_sc_hd__diode_2
XFILLER_2_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2054 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_57_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_183_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2098 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input302_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[14] sky130_fd_sc_hd__diode_2
XFILLER_183_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_1962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1859 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_188_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1748 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput500 vssd2 la_data_out[35] vccd1 _179_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_146_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput511 vssd2 la_data_out[45] vccd1 _189_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput522 vssd2 la_data_out[55] vccd1 _199_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_246_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput533 vssd2 la_data_out[65] vccd1 _209_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput544 vssd2 la_data_out[75] vccd1 _219_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_246_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput555 vssd2 la_data_out[85] vccd1 _229_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput566 vssd2 la_data_out[95] vccd1 _239_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput577 vssd2 wbs_dat_o[10] vccd1 _286_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput588 vssd2 wbs_dat_o[20] vccd1 _296_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput599 vssd2 wbs_dat_o[30] vccd1 _306_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_67_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_36 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_19_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__343__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_183_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_090_ vssd2 _344_/D _074_/A _089_/X vccd1 _088_/Y _072_/A _073_/X vccd1 vssd2 sky130_fd_sc_hd__o311a_1
XFILLER_155_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_668 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_40_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input252_A vssd2 vccd1 vccd1 vssd2 la_oenb[61] sky130_fd_sc_hd__diode_2
XFILLER_191_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_78_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_46_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_18_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
X_357_ _357_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _357_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_18_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_288_ _288_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_204_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput4 vssd2 input4/X vccd1 io_in[12] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_209_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_52_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_133_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_121_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput374 vssd2 io_oeb[15] vccd1 _116_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput385 vssd2 io_oeb[25] vccd1 _323_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput396 vssd2 io_oeb[35] vccd1 _333_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_82_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_801 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_215_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_42_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_834 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_143_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_211_ _211_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_867 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_221_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_11_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_142_ _142_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_195_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_073_ vssd2 _073_/X vccd1 _339_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_4
XFILLER_183_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input63_A vssd2 vccd1 vccd1 vssd2 la_data_in[121] sky130_fd_sc_hd__diode_2
XFILLER_174_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_570 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_115_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_111_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__338__A vssd2 vccd1 vccd1 vssd2 _338_/A sky130_fd_sc_hd__diode_2
XFILLER_168_1475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_40_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__073__A vssd2 vccd1 vccd1 vssd2 _339_/X sky130_fd_sc_hd__diode_2
XFILLER_179_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_43_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_558 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input215_A vssd2 vccd1 vccd1 vssd2 la_oenb[28] sky130_fd_sc_hd__diode_2
XFILLER_56_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XPHY_620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_62_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_631 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_686 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_125_ _125_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_11_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_056_ vssd2 _056_/X vccd1 _341_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_125_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output434_A vssd2 vccd1 vccd1 vssd2 _347_/Q sky130_fd_sc_hd__diode_2
XFILLER_238_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput40 vssd2 input40/X vccd1 la_data_in[100] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_147_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput51 vssd2 input51/X vccd1 la_data_in[110] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_190_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput62 vssd2 input62/X vccd1 la_data_in[120] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_162_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput73 vssd2 input73/X vccd1 la_data_in[15] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput84 vssd2 input84/X vccd1 la_data_in[25] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_196_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput95 vssd2 input95/X vccd1 la_data_in[35] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_190_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_49 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_187_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__068__A vssd2 vccd1 vccd1 vssd2 _341_/Q sky130_fd_sc_hd__diode_2
XFILLER_53_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_198_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_146_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_179_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input165_A vssd2 vccd1 vccd1 vssd2 la_data_in[99] sky130_fd_sc_hd__diode_2
XFILLER_0_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_79_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_431 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2030 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input332_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[11] sky130_fd_sc_hd__diode_2
XFILLER_103_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input26_A vssd2 vccd1 vccd1 vssd2 io_in[32] sky130_fd_sc_hd__diode_2
XFILLER_188_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2085 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_180_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_472 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_144_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_108_ _108_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_193_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_236_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_366 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_208_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1509 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1546 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_183_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_5 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_181_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input282_A vssd2 vccd1 vccd1 vssd2 la_oenb[89] sky130_fd_sc_hd__diode_2
XFILLER_5_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput230 vssd2 input230/X vccd1 la_oenb[41] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput241 vssd2 input241/X vccd1 la_oenb[51] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput252 vssd2 input252/X vccd1 la_oenb[61] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput263 vssd2 input263/X vccd1 la_oenb[71] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput274 vssd2 input274/X vccd1 la_oenb[81] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_229_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput285 vssd2 input285/X vccd1 la_oenb[91] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput296 vssd2 _335_/A vccd1 wb_rst_i vccd1 vssd2 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_223_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_216_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1078 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_44_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_985 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_236_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_104_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_11_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_159 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input128_A vssd2 vccd1 vccd1 vssd2 la_data_in[65] sky130_fd_sc_hd__diode_2
XFILLER_6_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.DAC_d0 vssd2 vccd1 vccd1 vssd2 adc.DAC/d0 sky130_fd_sc_hd__diode_2
XFILLER_205_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1387 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_148_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input93_A vssd2 vccd1 vccd1 vssd2 la_data_in[33] sky130_fd_sc_hd__diode_2
XFILLER_158_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_204_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_973 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_1974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_988 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_126_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_81_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_158_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput501 vssd2 la_data_out[36] vccd1 _180_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput512 vssd2 la_data_out[46] vccd1 _190_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput523 vssd2 la_data_out[56] vccd1 _200_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_246_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput534 vssd2 la_data_out[66] vccd1 _210_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput545 vssd2 la_data_out[76] vccd1 _220_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput556 vssd2 la_data_out[86] vccd1 _230_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_214_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput567 vssd2 la_data_out[96] vccd1 _240_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput578 vssd2 wbs_dat_o[11] vccd1 _287_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput589 vssd2 wbs_dat_o[21] vccd1 _297_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_214_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_242_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__076__A vssd2 vccd1 vccd1 vssd2 _076_/A sky130_fd_sc_hd__diode_2
XFILLER_223_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_145_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input245_A vssd2 vccd1 vccd1 vssd2 la_oenb[55] sky130_fd_sc_hd__diode_2
XFILLER_133_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__058__B1 vssd2 vccd1 vccd1 vssd2 _355_/Q sky130_fd_sc_hd__diode_2
XFILLER_232_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1103 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_356_ _356_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _356_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_35_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_287_ _287_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_155_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_217 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput5 vssd2 input5/X vccd1 io_in[13] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_211_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput375 vssd2 io_oeb[16] vccd1 _314_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput386 vssd2 io_oeb[26] vccd1 _324_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput397 vssd2 io_oeb[36] vccd1 _334_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_60_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_21_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_802 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_58_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_813 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_846 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_210_ _210_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XPHY_857 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_879 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_136_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_141_ _141_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_195_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input195_A vssd2 vccd1 vccd1 vssd2 la_oenb[125] sky130_fd_sc_hd__diode_2
XFILLER_137_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_072_ vssd2 _104_/A vccd1 _072_/A vccd1 vssd2 sky130_fd_sc_hd__buf_4
XFILLER_125_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input362_A vssd2 vccd1 vccd1 vssd2 wbs_sel_i[0] sky130_fd_sc_hd__diode_2
XFILLER_10_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input56_A vssd2 vccd1 vccd1 vssd2 la_data_in[115] sky130_fd_sc_hd__diode_2
XFILLER_133_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_222_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_339_ _339_/S vssd2 _339_/X _337_/A vccd1 _339_/A1 vccd1 vssd2 sky130_fd_sc_hd__mux2_8
XFILLER_187_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_582 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_2312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_20_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1644 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_16_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_240_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_668 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input110_A vssd2 vccd1 vccd1 vssd2 la_data_in[49] sky130_fd_sc_hd__diode_2
XANTENNA_input208_A vssd2 vccd1 vccd1 vssd2 la_oenb[21] sky130_fd_sc_hd__diode_2
XFILLER_204_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_610 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_643 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_62_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_124_ _124_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_200_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_193_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_055_ vssd2 _055_/X vccd1 _055_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_4
XFILLER_137_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__356__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_87_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_43_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput30 vssd2 input30/X vccd1 io_in[36] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput41 vssd2 input41/X vccd1 la_data_in[101] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_162_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput52 vssd2 input52/X vccd1 la_data_in[111] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_11_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput63 vssd2 input63/X vccd1 la_data_in[121] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_190_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput74 vssd2 input74/X vccd1 la_data_in[16] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_162_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput85 vssd2 input85/X vccd1 la_data_in[26] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput96 vssd2 input96/X vccd1 la_data_in[36] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_155_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__068__B vssd2 vccd1 vccd1 vssd2 _076_/A sky130_fd_sc_hd__diode_2
XFILLER_241_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_53_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_445 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input158_A vssd2 vccd1 vccd1 vssd2 la_data_in[92] sky130_fd_sc_hd__diode_2
XFILLER_153_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_48_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input325_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[6] sky130_fd_sc_hd__diode_2
XFILLER_235_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_75_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input19_A vssd2 vccd1 vccd1 vssd2 io_in[26] sky130_fd_sc_hd__diode_2
XFILLER_180_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_231_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_188_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_440 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_160_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_473 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_484 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_156_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_107_ _107_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_201_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_144_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_140_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_91_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_176_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_269 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__079__A vssd2 vccd1 vccd1 vssd2 _355_/Q sky130_fd_sc_hd__diode_2
XFILLER_187_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_57_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1558 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input275_A vssd2 vccd1 vccd1 vssd2 la_oenb[82] sky130_fd_sc_hd__diode_2
XFILLER_119_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_190_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_122_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput220 vssd2 input220/X vccd1 la_oenb[32] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput231 vssd2 input231/X vccd1 la_oenb[42] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_237_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput242 vssd2 input242/X vccd1 la_oenb[52] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput253 vssd2 input253/X vccd1 la_oenb[62] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput264 vssd2 input264/X vccd1 la_oenb[72] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput275 vssd2 input275/X vccd1 la_oenb[82] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_84_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput286 vssd2 input286/X vccd1 la_oenb[92] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_229_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput297 vssd2 input297/X vccd1 wbs_adr_i[0] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1057 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_90_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_997 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA_adc.DAC_out_v vssd2 vccd1 vccd1 vssd2 analog_io[3] sky130_fd_sc_hd__diode_2
XFILLER_152_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1521 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_184_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_11_1176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_100_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1318 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.DAC_d1 vssd2 vccd1 vccd1 vssd2 adc.DAC/d1 sky130_fd_sc_hd__diode_2
XFILLER_72_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_161_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input86_A vssd2 vccd1 vccd1 vssd2 la_data_in[27] sky130_fd_sc_hd__diode_2
XFILLER_70_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_1003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_7_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_237_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_240_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput502 vssd2 la_data_out[37] vccd1 _181_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput513 vssd2 la_data_out[47] vccd1 _191_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput524 vssd2 la_data_out[57] vccd1 _201_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput535 vssd2 la_data_out[67] vccd1 _211_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput546 vssd2 la_data_out[77] vccd1 _221_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput557 vssd2 la_data_out[87] vccd1 _231_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput568 vssd2 la_data_out[97] vccd1 _241_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_141_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_93 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput579 vssd2 wbs_dat_o[12] vccd1 _288_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_171_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_94_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1631 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1686 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_221_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_373 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_195_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_414 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_123_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_78_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__058__A1 vssd2 vccd1 vccd1 vssd2 _356_/Q sky130_fd_sc_hd__diode_2
XANTENNA_input140_A vssd2 vccd1 vccd1 vssd2 la_data_in[76] sky130_fd_sc_hd__diode_2
XFILLER_172_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__058__B2 vssd2 vccd1 vccd1 vssd2 _056_/X sky130_fd_sc_hd__diode_2
XFILLER_219_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input238_A vssd2 vccd1 vccd1 vssd2 la_oenb[49] sky130_fd_sc_hd__diode_2
XFILLER_115_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_86_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_74_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_60 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_355_ _355_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _355_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_126_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_286_ _286_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_127_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput6 vssd2 input6/X vccd1 io_in[14] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_83_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_168_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_37_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_145_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput376 vssd2 io_oeb[17] vccd1 _315_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput387 vssd2 io_oeb[27] vccd1 _325_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput398 vssd2 io_oeb[37] vccd1 _335_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_814 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_32_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_858 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_32_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_140_ _140_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_378 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_071_ vssd2 _071_/Y vccd1 _356_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_137_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input188_A vssd2 vccd1 vccd1 vssd2 la_oenb[119] sky130_fd_sc_hd__diode_2
XFILLER_191_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_701 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input355_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[3] sky130_fd_sc_hd__diode_2
XFILLER_105_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input49_A vssd2 vccd1 vccd1 vssd2 la_data_in[109] sky130_fd_sc_hd__diode_2
XFILLER_232_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_90 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_159_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_338_ vssd2 _338_/X vccd1 _338_/A vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_239_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_269_ _269_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_127_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_142_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_168_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_61 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_1827 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2357 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_37_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_87_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_5_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_188_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input103_A vssd2 vccd1 vccd1 vssd2 la_data_in[42] sky130_fd_sc_hd__diode_2
XPHY_611 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_644 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_62_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_655 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_688 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_156_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_123_ _123_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_205_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_054_ vssd2 _055_/A vccd1 _065_/A vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_124_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_152_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1000 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_78_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_1_1943 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_34_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1965 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput20 vssd2 input20/X vccd1 io_in[27] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput31 vssd2 input31/X vccd1 io_in[37] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_11_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput42 vssd2 input42/X vccd1 la_data_in[102] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput53 vssd2 input53/X vccd1 la_data_in[112] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_11_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput64 vssd2 input64/X vccd1 la_data_in[122] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_239_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput75 vssd2 input75/X vccd1 la_data_in[17] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_196_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput86 vssd2 input86/X vccd1 la_data_in[27] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput97 vssd2 input97/X vccd1 la_data_in[37] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_196_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xrepeater610 vssd2 _314_/A vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__buf_8
XFILLER_6_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1729 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_390 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_122_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA__103__B1 vssd2 vccd1 vccd1 vssd2 _103_/B1 sky130_fd_sc_hd__diode_2
XFILLER_115_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_153_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_170_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input220_A vssd2 vccd1 vccd1 vssd2 la_oenb[32] sky130_fd_sc_hd__diode_2
XFILLER_5_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input318_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[29] sky130_fd_sc_hd__diode_2
XFILLER_75_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1217 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_186_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_430 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_160_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_452 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_485 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_496 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_11_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_184_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_106_ vssd2 _357_/D _074_/X vccd1 _066_/A _055_/X vccd1 vssd2 sky130_fd_sc_hd__o21ai_1
XFILLER_7_166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_171_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_247_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_223_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_2100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_183_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__346__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_16_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input170_A vssd2 vccd1 vccd1 vssd2 la_oenb[102] sky130_fd_sc_hd__diode_2
XANTENNA_input268_A vssd2 vccd1 vccd1 vssd2 la_oenb[76] sky130_fd_sc_hd__diode_2
XFILLER_11_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput210 vssd2 input210/X vccd1 la_oenb[23] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput221 vssd2 input221/X vccd1 la_oenb[33] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input31_A vssd2 vccd1 vccd1 vssd2 io_in[37] sky130_fd_sc_hd__diode_2
XFILLER_7_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput232 vssd2 input232/X vccd1 la_oenb[43] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_102_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput243 vssd2 input243/X vccd1 la_oenb[53] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_237_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput254 vssd2 input254/X vccd1 la_oenb[63] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_274 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput265 vssd2 input265/X vccd1 la_oenb[73] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_229_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput276 vssd2 input276/X vccd1 la_oenb[83] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput287 vssd2 input287/X vccd1 la_oenb[93] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput298 vssd2 input298/X vccd1 wbs_adr_i[10] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_64_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_57_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_90_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_86_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1802 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1533 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_188_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_191_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_131_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2046 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_adc.DAC_d2 vssd2 vccd1 vccd1 vssd2 input15/X sky130_fd_sc_hd__diode_2
XFILLER_72_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input79_A vssd2 vccd1 vccd1 vssd2 la_data_in[20] sky130_fd_sc_hd__diode_2
XFILLER_202_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_42_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_221_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput503 vssd2 la_data_out[38] vccd1 _182_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput514 vssd2 la_data_out[48] vccd1 _192_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput525 vssd2 la_data_out[58] vccd1 _202_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput536 vssd2 la_data_out[68] vccd1 _212_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput547 vssd2 la_data_out[78] vccd1 _222_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput558 vssd2 la_data_out[88] vccd1 _232_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput569 vssd2 la_data_out[98] vccd1 _242_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1009 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__058__A2 vssd2 vccd1 vccd1 vssd2 _055_/X sky130_fd_sc_hd__diode_2
XFILLER_93_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_189_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input133_A vssd2 vccd1 vccd1 vssd2 la_data_in[6] sky130_fd_sc_hd__diode_2
XFILLER_73_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input300_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[12] sky130_fd_sc_hd__diode_2
XFILLER_2_1175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_61_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_121_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_354_ _354_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _354_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_41_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_285_ _285_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_224_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_123_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_993 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_111_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_49_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput7 vssd2 input7/X vccd1 io_in[15] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_64_422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_76_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1827 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_36_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_181_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_140_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_145_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
Xoutput377 vssd2 io_oeb[18] vccd1 _316_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_151_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput388 vssd2 io_oeb[28] vccd1 _326_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_233_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput399 vssd2 io_oeb[3] vccd1 _110_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_815 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_826 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_859 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_32_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_184_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_070_ vssd2 _349_/D _069_/Y vccd1 _349_/Q _066_/X vccd1 vssd2 sky130_fd_sc_hd__a21o_1
XFILLER_109_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_105_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input250_A vssd2 vccd1 vccd1 vssd2 la_oenb[5] sky130_fd_sc_hd__diode_2
XFILLER_120_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input348_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[26] sky130_fd_sc_hd__diode_2
XFILLER_238_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_80 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_91 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_337_ vssd2 _337_/X vccd1 _337_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_268_ _268_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_199_ _199_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_1839 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_95 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_65_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_53_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_701 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_178_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_153_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_87_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1546 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_623 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_656 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_239_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_667 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input298_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[10] sky130_fd_sc_hd__diode_2
XFILLER_156_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_122_ _122_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_158_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_053_ vssd2 _065_/A vccd1 _075_/A vccd1 _340_/Q vssd2 sky130_fd_sc_hd__nand2_2
XFILLER_109_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input61_A vssd2 vccd1 vccd1 vssd2 la_data_in[11] sky130_fd_sc_hd__diode_2
XFILLER_3_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_587 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_815 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_8_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_165_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_61_211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_35_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_929 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_672 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_206_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput10 vssd2 input10/X vccd1 io_in[18] vccd1 vssd2 sky130_fd_sc_hd__clkbuf_4
XFILLER_174_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput21 vssd2 _103_/B1 vccd1 io_in[28] vccd1 vssd2 sky130_fd_sc_hd__clkbuf_4
Xinput32 vssd2 input32/X vccd1 io_in[3] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput43 vssd2 input43/X vccd1 la_data_in[103] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_11_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput54 vssd2 input54/X vccd1 la_data_in[113] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_15_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput65 vssd2 input65/X vccd1 la_data_in[123] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput76 vssd2 input76/X vccd1 la_data_in[18] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput87 vssd2 input87/X vccd1 la_data_in[28] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput98 vssd2 input98/X vccd1 la_data_in[38] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_104_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xrepeater611 vssd2 _331_/A vccd1 _335_/A vccd1 vssd2 sky130_fd_sc_hd__buf_8
XFILLER_245_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_181_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1418 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__103__A1 vssd2 vccd1 vccd1 vssd2 _055_/X sky130_fd_sc_hd__diode_2
XANTENNA__103__B2 vssd2 vccd1 vccd1 vssd2 _069_/Y sky130_fd_sc_hd__diode_2
XFILLER_88_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_87_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_489 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input213_A vssd2 vccd1 vccd1 vssd2 la_oenb[26] sky130_fd_sc_hd__diode_2
XFILLER_90_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_188_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_431 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_464 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_40_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_497 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1941 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_105_ vssd2 _326_/A vccd1 _105_/A vccd1 vssd2 sky130_fd_sc_hd__buf_6
XFILLER_156_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output432_A vssd2 vccd1 vccd1 vssd2 _345_/Q sky130_fd_sc_hd__diode_2
XFILLER_234_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_213_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_113_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_38_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_241_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_178_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_159 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_134_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input163_A vssd2 vccd1 vccd1 vssd2 la_data_in[97] sky130_fd_sc_hd__diode_2
XFILLER_134_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput200 vssd2 input200/X vccd1 la_oenb[14] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput211 vssd2 input211/X vccd1 la_oenb[24] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput222 vssd2 input222/X vccd1 la_oenb[34] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input330_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[0] sky130_fd_sc_hd__diode_2
XFILLER_68_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput233 vssd2 input233/X vccd1 la_oenb[44] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_7_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput244 vssd2 input244/X vccd1 la_oenb[54] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_102_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput255 vssd2 input255/X vccd1 la_oenb[64] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_130_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput266 vssd2 input266/X vccd1 la_oenb[74] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput277 vssd2 input277/X vccd1 la_oenb[84] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_5_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input24_A vssd2 vccd1 vccd1 vssd2 io_in[30] sky130_fd_sc_hd__diode_2
Xinput288 vssd2 input288/X vccd1 la_oenb[94] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput299 vssd2 input299/X vccd1 wbs_adr_i[11] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_217_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_261 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_98_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_200_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_129 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_116_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1230 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_adc.DAC_d3 vssd2 vccd1 vccd1 vssd2 input14/X sky130_fd_sc_hd__diode_2
XFILLER_227_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_659 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1357 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_159_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input280_A vssd2 vccd1 vccd1 vssd2 la_oenb[87] sky130_fd_sc_hd__diode_2
XFILLER_202_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_969 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_194_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_231_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_135_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput504 vssd2 la_data_out[39] vccd1 _183_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_145_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput515 vssd2 la_data_out[49] vccd1 _193_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput526 vssd2 la_data_out[59] vccd1 _203_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput537 vssd2 la_data_out[69] vccd1 _213_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput548 vssd2 la_data_out[79] vccd1 _223_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_216_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput559 vssd2 la_data_out[89] vccd1 _233_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_73 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_113_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_19_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_145_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input126_A vssd2 vccd1 vccd1 vssd2 la_data_in[63] sky130_fd_sc_hd__diode_2
XFILLER_171_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_353_ _353_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _353_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_230_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input91_A vssd2 vccd1 vccd1 vssd2 la_data_in[31] sky130_fd_sc_hd__diode_2
X_284_ _284_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_139_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_49_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput8 vssd2 input8/X vccd1 io_in[16] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_49_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1806 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_181_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_20_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput378 vssd2 io_oeb[19] vccd1 _317_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_151_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput389 vssd2 io_oeb[29] vccd1 _327_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_805 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_827 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_838 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_212_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input243_A vssd2 vccd1 vccd1 vssd2 la_oenb[53] sky130_fd_sc_hd__diode_2
XFILLER_8_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_81 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_186_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_92 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_336_ vssd2 _336_/X vccd1 _336_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_4
XFILLER_186_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_267_ _267_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_239_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_198_ _198_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_109_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2147 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1603 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_53_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_217_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_214_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1558 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_602 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_635 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_123_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_162_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_668 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_121_ _121_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_184_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_240_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input193_A vssd2 vccd1 vccd1 vssd2 la_oenb[123] sky130_fd_sc_hd__diode_2
XFILLER_158_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_052_ vssd2 _075_/A vccd1 _341_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_158_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input360_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[8] sky130_fd_sc_hd__diode_2
XFILLER_152_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input54_A vssd2 vccd1 vccd1 vssd2 la_data_in[113] sky130_fd_sc_hd__diode_2
XFILLER_238_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_599 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_82_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_188_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_206_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_319_ vssd2 _319_/X vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput11 vssd2 input11/X vccd1 io_in[19] vccd1 vssd2 sky130_fd_sc_hd__buf_4
XFILLER_223_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput22 vssd2 input22/X vccd1 io_in[29] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_156_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput33 vssd2 input33/X vccd1 io_in[4] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput44 vssd2 input44/X vccd1 la_data_in[104] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput55 vssd2 input55/X vccd1 la_data_in[114] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput66 vssd2 input66/X vccd1 la_data_in[124] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput77 vssd2 input77/X vccd1 la_data_in[19] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_116_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput88 vssd2 input88/X vccd1 la_data_in[29] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_182_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput99 vssd2 input99/X vccd1 la_data_in[39] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_174_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_269 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xrepeater612 vssd2 adc.DAC/d0 vccd1 input17/X vccd1 vssd2 sky130_fd_sc_hd__buf_8
XFILLER_84_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_245_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1243 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_52_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_213_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_402 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input206_A vssd2 vccd1 vccd1 vssd2 la_oenb[1] sky130_fd_sc_hd__diode_2
XFILLER_16_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_443 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_476 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_106_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_40_974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_104_ vssd2 _341_/D vccd1 _104_/A vccd1 _104_/B vssd2 sky130_fd_sc_hd__nor2_1
XFILLER_10_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_120_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_993 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_241_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1517 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1445 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_96_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input156_A vssd2 vccd1 vccd1 vssd2 la_data_in[90] sky130_fd_sc_hd__diode_2
Xinput201 vssd2 input201/X vccd1 la_oenb[15] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_68_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput212 vssd2 input212/X vccd1 la_oenb[25] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput223 vssd2 input223/X vccd1 la_oenb[35] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput234 vssd2 input234/X vccd1 la_oenb[45] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput245 vssd2 input245/X vccd1 la_oenb[55] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput256 vssd2 input256/X vccd1 la_oenb[65] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input323_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[4] sky130_fd_sc_hd__diode_2
Xinput267 vssd2 input267/X vccd1 la_oenb[75] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput278 vssd2 input278/X vccd1 la_oenb[85] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_64_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput289 vssd2 input289/X vccd1 la_oenb[95] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input17_A vssd2 vccd1 vccd1 vssd2 io_in[24] sky130_fd_sc_hd__diode_2
XFILLER_245_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_220_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_273 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_145_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output375_A vssd2 vccd1 vccd1 vssd2 _314_/X sky130_fd_sc_hd__diode_2
XFILLER_69_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_138_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_160 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_98_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1572 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_62_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_395 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_50_535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_135_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_239_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input9_A vssd2 vccd1 vccd1 vssd2 io_in[17] sky130_fd_sc_hd__diode_2
XFILLER_58_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1314 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_227_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_adc.DAC_d4 vssd2 vccd1 vccd1 vssd2 input13/X sky130_fd_sc_hd__diode_2
XFILLER_214_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_660 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_199_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_220_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_414 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_148_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input273_A vssd2 vccd1 vccd1 vssd2 la_oenb[80] sky130_fd_sc_hd__diode_2
XFILLER_135_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_235_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1888 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_220_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_199_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_47_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput505 vssd2 la_data_out[3] vccd1 _147_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput516 vssd2 la_data_out[4] vccd1 _148_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput527 vssd2 la_data_out[5] vccd1 _149_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput538 vssd2 la_data_out[6] vccd1 _150_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_181_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput549 vssd2 la_data_out[7] vccd1 _151_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_125_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2313 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_117_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_219_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input119_A vssd2 vccd1 vccd1 vssd2 la_data_in[57] sky130_fd_sc_hd__diode_2
XFILLER_226_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_352_ _352_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _352_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_121_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_283_ _283_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_139_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input84_A vssd2 vccd1 vccd1 vssd2 la_data_in[25] sky130_fd_sc_hd__diode_2
XFILLER_154_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_110_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
Xinput9 vssd2 input9/X vccd1 io_in[17] vccd1 vssd2 sky130_fd_sc_hd__buf_6
XFILLER_49_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1818 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput368 vssd2 io_oeb[0] vccd1 _107_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput379 vssd2 io_oeb[1] vccd1 _108_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_206_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_806 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_817 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_839 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_117_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input236_A vssd2 vccd1 vccd1 vssd2 la_oenb[47] sky130_fd_sc_hd__diode_2
XFILLER_76_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_60 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_92_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_186_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_93 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_335_ vssd2 _335_/X vccd1 _335_/A vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_202_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_186_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_871 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_266_ _266_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_41_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_197_ _197_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_237_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_75 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_65_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2159 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1615 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_61_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_639 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_203_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_603 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA__349__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XPHY_614 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_227_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_647 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_123_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_162_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_196_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_120_ _120_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_221_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input186_A vssd2 vccd1 vccd1 vssd2 la_oenb[117] sky130_fd_sc_hd__diode_2
XFILLER_193_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_164_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__106__B1 vssd2 vccd1 vccd1 vssd2 _074_/X sky130_fd_sc_hd__diode_2
XFILLER_238_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_3_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input353_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[30] sky130_fd_sc_hd__diode_2
XFILLER_152_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input47_A vssd2 vccd1 vccd1 vssd2 la_data_in[107] sky130_fd_sc_hd__diode_2
XFILLER_43_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_239_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_235_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_318_ vssd2 _318_/X vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput12 vssd2 input12/X vccd1 io_in[1] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_102_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput23 vssd2 input23/X vccd1 io_in[2] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput34 vssd2 input34/X vccd1 io_in[5] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_128_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput45 vssd2 input45/X vccd1 la_data_in[105] vccd1 vssd2 sky130_fd_sc_hd__buf_1
X_249_ _249_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_15_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput56 vssd2 input56/X vccd1 la_data_in[115] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_156_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput67 vssd2 input67/X vccd1 la_data_in[125] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput78 vssd2 input78/X vccd1 la_data_in[1] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_174_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput89 vssd2 input89/X vccd1 la_data_in[2] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_116_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xrepeater613 vssd2 adc.DAC/d1 vccd1 input16/X vccd1 vssd2 sky130_fd_sc_hd__buf_8
XFILLER_69_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_59_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_217_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_31_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input101_A vssd2 vccd1 vccd1 vssd2 la_data_in[40] sky130_fd_sc_hd__diode_2
XPHY_411 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_24_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_488 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_40_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_103_ vssd2 _340_/D _103_/B1 vccd1 _069_/Y _055_/X _104_/B vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_138_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_502 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_138_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_179_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1798 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_22_419 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_175_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_239_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_246_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1074 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_1228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_146_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput202 vssd2 input202/X vccd1 la_oenb[16] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_44_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_131_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput213 vssd2 input213/X vccd1 la_oenb[26] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput224 vssd2 input224/X vccd1 la_oenb[36] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_213_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input149_A vssd2 vccd1 vccd1 vssd2 la_data_in[84] sky130_fd_sc_hd__diode_2
XFILLER_194_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput235 vssd2 input235/X vccd1 la_oenb[46] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_124_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput246 vssd2 input246/X vccd1 la_oenb[56] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput257 vssd2 input257/X vccd1 la_oenb[66] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput268 vssd2 input268/X vccd1 la_oenb[76] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput279 vssd2 input279/X vccd1 la_oenb[86] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA_input316_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[27] sky130_fd_sc_hd__diode_2
XFILLER_91_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1028 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_84_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_217_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_230 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_274 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_285 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_8_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_113_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_84_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_2241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2285 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_8_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.DAC_d5 vssd2 vccd1 vccd1 vssd2 input11/X sky130_fd_sc_hd__diode_2
XFILLER_22_1276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_672 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_107_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input266_A vssd2 vccd1 vccd1 vssd2 la_oenb[74] sky130_fd_sc_hd__diode_2
XFILLER_135_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_62_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_95_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_166_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output485_A vssd2 vccd1 vccd1 vssd2 _165_/LO sky130_fd_sc_hd__diode_2
XFILLER_199_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_200_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput506 vssd2 la_data_out[40] vccd1 _184_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput517 vssd2 la_data_out[50] vccd1 _194_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput528 vssd2 la_data_out[60] vccd1 _204_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_125_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput539 vssd2 la_data_out[70] vccd1 _214_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_125_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1370 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_407 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_132_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_120_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_187_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_351_ _351_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _351_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_242_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_282_ _282_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_202_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input77_A vssd2 vccd1 vccd1 vssd2 la_data_in[19] sky130_fd_sc_hd__diode_2
XFILLER_237_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_190_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_1_462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_172_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_484 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_39_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__101__A vssd2 vccd1 vccd1 vssd2 _357_/Q sky130_fd_sc_hd__diode_2
XFILLER_188_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput369 vssd2 io_oeb[10] vccd1 _311_/X vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_243_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_149_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1476 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_818 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_829 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input131_A vssd2 vccd1 vccd1 vssd2 la_data_in[68] sky130_fd_sc_hd__diode_2
XFILLER_47_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input229_A vssd2 vccd1 vccd1 vssd2 la_oenb[40] sky130_fd_sc_hd__diode_2
XFILLER_132_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_570 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_50 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_61 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_214_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_42_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_334_ vssd2 _334_/X vccd1 _335_/A vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_41_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_265_ _265_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_883 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_196_ _196_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_32 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__060__B1 vssd2 vccd1 vccd1 vssd2 _353_/Q sky130_fd_sc_hd__diode_2
XFILLER_178_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_99_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_29_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_615 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_162_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_659 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_211_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_178_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input179_A vssd2 vccd1 vccd1 vssd2 la_oenb[110] sky130_fd_sc_hd__diode_2
XFILLER_164_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input346_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[24] sky130_fd_sc_hd__diode_2
XFILLER_132_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_130_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1914 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1958 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_226_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_317_ vssd2 _317_/X vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XANTENNA_output398_A vssd2 vccd1 vccd1 vssd2 _335_/X sky130_fd_sc_hd__diode_2
XFILLER_175_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_680 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput13 vssd2 input13/X vccd1 io_in[20] vccd1 vssd2 sky130_fd_sc_hd__buf_6
XFILLER_223_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_248_ _248_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
Xinput24 vssd2 input24/X vccd1 io_in[30] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput35 vssd2 input35/X vccd1 io_in[6] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_239_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput46 vssd2 input46/X vccd1 la_data_in[106] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_128_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput57 vssd2 input57/X vccd1 la_data_in[116] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput68 vssd2 input68/X vccd1 la_data_in[126] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_239_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.DAC_inp1 vssd2 vccd1 vccd1 vssd2 analog_io[2] sky130_fd_sc_hd__diode_2
XFILLER_143_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_179_ _179_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
Xinput79 vssd2 input79/X vccd1 la_data_in[20] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_139_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_228_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_224_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_193_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_401 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_189_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_445 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_456 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_237_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_489 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_185_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input296_A vssd2 vccd1 vccd1 vssd2 wb_rst_i sky130_fd_sc_hd__diode_2
XFILLER_16_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_102_ vssd2 _104_/B vccd1 _353_/Q vccd1 _352_/Q vssd2 _102_/C _102_/D sky130_fd_sc_hd__or4_4
XFILLER_12_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_159 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_125_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_239_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_960 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_659 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1086 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_179_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_139_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput203 vssd2 input203/X vccd1 la_oenb[17] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput214 vssd2 input214/X vccd1 la_oenb[27] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput225 vssd2 input225/X vccd1 la_oenb[37] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput236 vssd2 input236/X vccd1 la_oenb[47] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput247 vssd2 input247/X vccd1 la_oenb[57] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_5_1110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput258 vssd2 input258/X vccd1 la_oenb[67] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_9_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput269 vssd2 input269/X vccd1 la_oenb[77] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_187_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_56_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input211_A vssd2 vccd1 vccd1 vssd2 la_oenb[24] sky130_fd_sc_hd__diode_2
XANTENNA_input309_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[20] sky130_fd_sc_hd__diode_2
XFILLER_140_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_164_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_8_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_3_140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA__104__A vssd2 vccd1 vccd1 vssd2 _104_/A sky130_fd_sc_hd__diode_2
XFILLER_171_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_696 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_106_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output430_A vssd2 vccd1 vccd1 vssd2 _343_/Q sky130_fd_sc_hd__diode_2
XFILLER_121_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_143_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_66_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_adc.DAC_d6 vssd2 vccd1 vccd1 vssd2 input10/X sky130_fd_sc_hd__diode_2
XFILLER_22_1288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_70_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_5_438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_107_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_150_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input161_A vssd2 vccd1 vccd1 vssd2 la_data_in[95] sky130_fd_sc_hd__diode_2
XFILLER_1_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_172_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input259_A vssd2 vccd1 vccd1 vssd2 la_oenb[68] sky130_fd_sc_hd__diode_2
XFILLER_1_644 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_235_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_103_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input22_A vssd2 vccd1 vccd1 vssd2 io_in[29] sky130_fd_sc_hd__diode_2
XFILLER_236_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_151_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_28_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_166_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1857 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1582 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput507 vssd2 la_data_out[41] vccd1 _185_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_138_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput518 vssd2 la_data_out[51] vccd1 _195_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput529 vssd2 la_data_out[61] vccd1 _205_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_99_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_65 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_125_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_231_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_224_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_378 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_121_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1085 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_198_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_350_ _350_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _350_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_198_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_281_ _281_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_14_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_430 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__101__B vssd2 vccd1 vccd1 vssd2 _356_/Q sky130_fd_sc_hd__diode_2
XFILLER_188_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1488 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_221_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input124_A vssd2 vccd1 vccd1 vssd2 la_data_in[61] sky130_fd_sc_hd__diode_2
XFILLER_128_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_40 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_245_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XPHY_62 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_582 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_73 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_333_ vssd2 _333_/X vccd1 _335_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XPHY_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_95 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_42_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_264_ _264_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_52_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_895 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_195_ _195_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_87_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_55 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__060__A1 vssd2 vccd1 vccd1 vssd2 _354_/Q sky130_fd_sc_hd__diode_2
XANTENNA__060__B2 vssd2 vccd1 vccd1 vssd2 _056_/X sky130_fd_sc_hd__diode_2
XFILLER_221_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_102_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_616 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_627 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_141_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__106__A2 vssd2 vccd1 vccd1 vssd2 _055_/X sky130_fd_sc_hd__diode_2
XFILLER_106_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input241_A vssd2 vccd1 vccd1 vssd2 la_oenb[51] sky130_fd_sc_hd__diode_2
XFILLER_132_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input339_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[18] sky130_fd_sc_hd__diode_2
XFILLER_232_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_28_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_316_ vssd2 _316_/X vccd1 _316_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_141_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput14 vssd2 input14/X vccd1 io_in[21] vccd1 vssd2 sky130_fd_sc_hd__buf_6
XFILLER_204_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_247_ _247_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_692 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput25 vssd2 input25/X vccd1 io_in[31] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_128_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput36 vssd2 input36/X vccd1 io_in[7] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_204_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput47 vssd2 input47/X vccd1 la_data_in[107] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_128_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput58 vssd2 input58/X vccd1 la_data_in[117] vccd1 vssd2 sky130_fd_sc_hd__buf_1
X_178_ _178_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
Xinput69 vssd2 input69/X vccd1 la_data_in[127] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_171_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_96_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_211_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_19_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1458 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2015 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_402 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_52_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_5 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_468 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_8_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_101_ vssd2 _102_/D vccd1 _357_/Q vccd1 _356_/Q vssd2 _355_/Q _354_/Q sky130_fd_sc_hd__or4_4
XFILLER_16_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input191_A vssd2 vccd1 vccd1 vssd2 la_oenb[121] sky130_fd_sc_hd__diode_2
XFILLER_165_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input289_A vssd2 vccd1 vccd1 vssd2 la_oenb[95] sky130_fd_sc_hd__diode_2
XFILLER_138_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input52_A vssd2 vccd1 vccd1 vssd2 la_data_in[111] sky130_fd_sc_hd__diode_2
XFILLER_106_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_121_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_78_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_972 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1712 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_147_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_160 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_239_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1509 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_113_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_671 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_168_1098 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_230_64 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_179_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_222_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput204 vssd2 input204/X vccd1 la_oenb[18] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput215 vssd2 input215/X vccd1 la_oenb[28] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput226 vssd2 input226/X vccd1 la_oenb[38] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_248_257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_131_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput237 vssd2 input237/X vccd1 la_oenb[48] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_236_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput248 vssd2 input248/X vccd1 la_oenb[58] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput259 vssd2 input259/X vccd1 la_oenb[68] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_5_1122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_124_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_232_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input204_A vssd2 vccd1 vccd1 vssd2 la_oenb[18] sky130_fd_sc_hd__diode_2
XFILLER_140_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1616 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_243 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_129_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_157_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_10_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1586 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_225_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_53_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.DAC_d7 vssd2 vccd1 vccd1 vssd2 input9/X sky130_fd_sc_hd__diode_2
XFILLER_241_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_198_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_224_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1005 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_222_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_135_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input154_A vssd2 vccd1 vccd1 vssd2 la_data_in[89] sky130_fd_sc_hd__diode_2
XFILLER_77_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_1009 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_103_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input321_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[31] sky130_fd_sc_hd__diode_2
XFILLER_131_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input15_A vssd2 vccd1 vccd1 vssd2 io_in[22] sky130_fd_sc_hd__diode_2
XFILLER_2_1851 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_166_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_204_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2147 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput508 vssd2 la_data_out[42] vccd1 _186_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_99_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput519 vssd2 la_data_out[52] vccd1 _196_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_67_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_243 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input7_A vssd2 vccd1 vccd1 vssd2 io_in[15] sky130_fd_sc_hd__diode_2
XFILLER_100_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_230_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1103 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_280_ _280_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_14_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input271_A vssd2 vccd1 vccd1 vssd2 la_oenb[79] sky130_fd_sc_hd__diode_2
XFILLER_146_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_122_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__101__C vssd2 vccd1 vccd1 vssd2 _355_/Q sky130_fd_sc_hd__diode_2
XFILLER_77_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_218_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_132_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_1_1180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_243_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_50_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_136_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_191_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input117_A vssd2 vccd1 vccd1 vssd2 la_data_in[55] sky130_fd_sc_hd__diode_2
XFILLER_128_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_226_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_41 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_52 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_63 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_74 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_332_ vssd2 _332_/X vccd1 _335_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XPHY_85 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_42_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_263_ _263_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1886 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input82_A vssd2 vccd1 vccd1 vssd2 la_data_in[23] sky130_fd_sc_hd__diode_2
XFILLER_128_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
X_194_ _194_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_100_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_221_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_124_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_237_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_89 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2142 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_168_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_92_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA__060__A2 vssd2 vccd1 vccd1 vssd2 _055_/A sky130_fd_sc_hd__diode_2
XFILLER_233_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1973 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_639 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__339__A0 vssd2 vccd1 vccd1 vssd2 _337_/A sky130_fd_sc_hd__diode_2
XFILLER_180_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_485 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_5 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_106_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_47_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input234_A vssd2 vccd1 vccd1 vssd2 la_oenb[45] sky130_fd_sc_hd__diode_2
XFILLER_247_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_243_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_315_ vssd2 _315_/X vccd1 _316_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_246_ _246_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
Xinput15 vssd2 input15/X vccd1 io_in[22] vccd1 vssd2 sky130_fd_sc_hd__buf_8
XFILLER_204_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput26 vssd2 input26/X vccd1 io_in[32] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_168_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput37 vssd2 input37/X vccd1 io_in[8] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_183_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput48 vssd2 input48/X vccd1 la_data_in[108] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_155_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput59 vssd2 input59/X vccd1 la_data_in[118] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_139_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_177_ _177_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_59_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_98_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_614 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_60_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_161_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_103_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1770 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_403 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_225_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_414 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_52_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_458 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_100_ vssd2 _102_/C vccd1 _351_/Q vccd1 _100_/B vssd2 sky130_fd_sc_hd__or2_1
XFILLER_240_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input184_A vssd2 vccd1 vccd1 vssd2 la_oenb[115] sky130_fd_sc_hd__diode_2
XFILLER_165_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input351_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[29] sky130_fd_sc_hd__diode_2
XFILLER_133_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input45_A vssd2 vccd1 vccd1 vssd2 la_data_in[105] sky130_fd_sc_hd__diode_2
XFILLER_191_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_78_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_47_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_60 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_981 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_229_ _229_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_155_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1416 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_214_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_187_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_179_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_107_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput205 vssd2 input205/X vccd1 la_oenb[19] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput216 vssd2 input216/X vccd1 la_oenb[29] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput227 vssd2 input227/X vccd1 la_oenb[39] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput238 vssd2 input238/X vccd1 la_oenb[49] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_131_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput249 vssd2 input249/X vccd1 la_oenb[59] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_75_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1972 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_56_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_204_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_200 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_140_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_207_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_32_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_175_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_218_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_79_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_181_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_47_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_56_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__311__A vssd2 vccd1 vccd1 vssd2 _314_/A sky130_fd_sc_hd__diode_2
XFILLER_174_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_224_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1017 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_181_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_407 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_119_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_190_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input147_A vssd2 vccd1 vccd1 vssd2 la_data_in[82] sky130_fd_sc_hd__diode_2
XFILLER_95_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input314_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[25] sky130_fd_sc_hd__diode_2
XFILLER_233_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_686 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2159 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xadc.SCOMP wb_clk_i analog_io[5] analog_io[4] _336_/A vccd2 vssd2 ACMP_HVL
XFILLER_71_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_146_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput509 vssd2 la_data_out[43] vccd1 _187_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2030 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2074 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__090__B1 vssd2 vccd1 vccd1 vssd2 _074_/A sky130_fd_sc_hd__diode_2
XFILLER_63_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_100_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__081__B1 vssd2 vccd1 vccd1 vssd2 _074_/X sky130_fd_sc_hd__diode_2
XFILLER_164_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1860 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_172_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input264_A vssd2 vccd1 vccd1 vssd2 la_oenb[72] sky130_fd_sc_hd__diode_2
XFILLER_190_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_89_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__101__D vssd2 vccd1 vccd1 vssd2 _354_/Q sky130_fd_sc_hd__diode_2
XFILLER_77_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_233_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_195_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_190_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2114 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_110_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_212_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_1_1192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_176_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_603 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_151_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_9 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_219_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_20 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_226_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_331_ vssd2 _331_/X vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XPHY_64 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_187_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_75 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_86 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_97 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_842 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_262_ _262_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_208_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_193_ _193_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_155_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input75_A vssd2 vccd1 vccd1 vssd2 la_data_in[17] sky130_fd_sc_hd__diode_2
XFILLER_87_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_215_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_68 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_2176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_179_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1085 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_31_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1985 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_52_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_629 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_720 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_121_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input227_A vssd2 vccd1 vccd1 vssd2 la_oenb[39] sky130_fd_sc_hd__diode_2
XFILLER_74_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_545 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_217 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_314_ vssd2 _314_/X vccd1 _314_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_70_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_245_ _245_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_180_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput16 vssd2 input16/X vccd1 io_in[23] vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput27 vssd2 input27/X vccd1 io_in[33] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_155_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput38 vssd2 input38/X vccd1 io_in[9] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_196_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_176_ _176_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
Xinput49 vssd2 input49/X vccd1 la_data_in[109] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_183_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_98_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_168_1248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_179_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1295 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__314__A vssd2 vccd1 vccd1 vssd2 _314_/A sky130_fd_sc_hd__diode_2
XFILLER_173_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_407 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_42_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_415 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_52_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1972 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input177_A vssd2 vccd1 vccd1 vssd2 la_oenb[109] sky130_fd_sc_hd__diode_2
XFILLER_118_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_133_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input344_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[22] sky130_fd_sc_hd__diode_2
XFILLER_248_941 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA_input38_A vssd2 vccd1 vccd1 vssd2 io_in[9] sky130_fd_sc_hd__diode_2
XFILLER_121_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_93_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1725 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1769 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_72 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_960 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_54_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_228_ _228_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_10_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_159_ _159_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_217_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_173 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_repeater609_A vssd2 vccd1 vccd1 vssd2 _326_/A sky130_fd_sc_hd__diode_2
XFILLER_217_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2129 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_226_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1045 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__309__A vssd2 vccd1 vccd1 vssd2 _316_/A sky130_fd_sc_hd__diode_2
XFILLER_185_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_194_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_190_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_204 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput206 vssd2 input206/X vccd1 la_oenb[1] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_216_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput217 vssd2 input217/X vccd1 la_oenb[2] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_103_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput228 vssd2 input228/X vccd1 la_oenb[3] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_170_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput239 vssd2 input239/X vccd1 la_oenb[4] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_75_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1984 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_246_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_212 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_140_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_256 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_235_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input294_A vssd2 vccd1 vccd1 vssd2 la_oenb[9] sky130_fd_sc_hd__diode_2
XFILLER_200_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_205_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_140_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_88_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1500 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1566 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_108_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_972 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_144_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__352__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_245_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_26_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1029 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_89_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_85_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1781 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input307_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[19] sky130_fd_sc_hd__diode_2
XFILLER_207_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1541 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_430 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_79 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_79_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_94_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_1_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_223_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_176_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__322__A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_172_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_871 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_11_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input257_A vssd2 vccd1 vccd1 vssd2 la_oenb[66] sky130_fd_sc_hd__diode_2
XFILLER_2_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_215_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input20_A vssd2 vccd1 vccd1 vssd2 io_in[27] sky130_fd_sc_hd__diode_2
XFILLER_64_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1672 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_214_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__063__A1 vssd2 vccd1 vccd1 vssd2 _351_/Q sky130_fd_sc_hd__diode_2
XANTENNA__063__B2 vssd2 vccd1 vccd1 vssd2 _341_/Q sky130_fd_sc_hd__diode_2
XFILLER_222_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__317__A vssd2 vccd1 vccd1 vssd2 _323_/A sky130_fd_sc_hd__diode_2
XFILLER_182_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__052__A vssd2 vccd1 vccd1 vssd2 _341_/Q sky130_fd_sc_hd__diode_2
XFILLER_191_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_10 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_21 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_82_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_32 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_215_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_65 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_330_ vssd2 _330_/X vccd1 _331_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_76 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_98 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_261_ _261_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_243_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_192_ _192_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_183_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input68_A vssd2 vccd1 vccd1 vssd2 la_data_in[126] sky130_fd_sc_hd__diode_2
XFILLER_237_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_692 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_215_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2155 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_209_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_222_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1200 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1997 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_517 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1907 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input122_A vssd2 vccd1 vccd1 vssd2 la_data_in[5] sky130_fd_sc_hd__diode_2
XFILLER_74_557 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_313_ vssd2 _313_/X vccd1 _316_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_230_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_244_ _244_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput17 vssd2 input17/X vccd1 io_in[24] vccd1 vssd2 sky130_fd_sc_hd__buf_2
XFILLER_195_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_167_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput28 vssd2 input28/X vccd1 io_in[34] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_13_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput39 vssd2 input39/X vccd1 la_data_in[0] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_155_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_175_ _175_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_196_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_202_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_139_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__330__A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_244_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_83_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_416 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_427 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput490 vssd2 la_data_out[26] vccd1 _170_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input337_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[16] sky130_fd_sc_hd__diode_2
XFILLER_248_953 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_84 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_30_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_972 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_227_ _227_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_129_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_158_ _158_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_195_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_089_ vssd2 _089_/X _344_/Q vccd1 _075_/A _076_/A _353_/Q vccd1 vssd2 sky130_fd_sc_hd__a31o_1
XFILLER_170_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_26_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1057 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__325__A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_18_1093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_119_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_216 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput207 vssd2 input207/X vccd1 la_oenb[20] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_130_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput218 vssd2 input218/X vccd1 la_oenb[30] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput229 vssd2 input229/X vccd1 la_oenb[40] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_57_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_112_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_44_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_246_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_257 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_199_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input287_A vssd2 vccd1 vccd1 vssd2 la_oenb[93] sky130_fd_sc_hd__diode_2
XFILLER_177_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_152_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A vssd2 vccd1 vccd1 vssd2 la_data_in[10] sky130_fd_sc_hd__diode_2
XFILLER_180_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_50 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_63_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_108_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_80 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_241_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__055__A vssd2 vccd1 vccd1 vssd2 _055_/A sky130_fd_sc_hd__diode_2
XFILLER_166_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_89_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_218_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_611 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_85_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1843 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_246_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1793 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1887 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input202_A vssd2 vccd1 vccd1 vssd2 la_oenb[16] sky130_fd_sc_hd__diode_2
XFILLER_207_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_44_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_53_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input98_A vssd2 vccd1 vccd1 vssd2 la_data_in[38] sky130_fd_sc_hd__diode_2
XFILLER_16_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_976 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_154_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_119_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_692 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_48_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_47_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_47_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_75_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_184_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__090__A2 vssd2 vccd1 vccd1 vssd2 _072_/A sky130_fd_sc_hd__diode_2
XFILLER_188_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_530 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_215_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__081__A2 vssd2 vccd1 vccd1 vssd2 _104_/A sky130_fd_sc_hd__diode_2
XFILLER_215_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_247_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_883 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_172_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input152_A vssd2 vccd1 vccd1 vssd2 la_data_in[87] sky130_fd_sc_hd__diode_2
XFILLER_215_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2330 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input13_A vssd2 vccd1 vccd1 vssd2 io_in[20] sky130_fd_sc_hd__diode_2
XFILLER_57_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_245_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_22_1590 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1684 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_246_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_201_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_185_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__342__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_9_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__063__A2 vssd2 vccd1 vccd1 vssd2 _055_/A sky130_fd_sc_hd__diode_2
XFILLER_225_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__333__A vssd2 vccd1 vccd1 vssd2 _335_/A sky130_fd_sc_hd__diode_2
XFILLER_118_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input5_A vssd2 vccd1 vccd1 vssd2 io_in[13] sky130_fd_sc_hd__diode_2
XFILLER_189_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_11 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_22 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_1993 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_33 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_82_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_44 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_109_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_55 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_77 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_88 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_260_ _260_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_17_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_167_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_680 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_195_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_191_ _191_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_155_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input367_A vssd2 vccd1 vccd1 vssd2 wbs_we_i sky130_fd_sc_hd__diode_2
XFILLER_191_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_237_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_248_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_18_2168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_32_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1212 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__328__A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_212_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_209_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_129 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_180_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input115_A vssd2 vccd1 vccd1 vssd2 la_data_in[53] sky130_fd_sc_hd__diode_2
XFILLER_243_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_312_ vssd2 _312_/X vccd1 _316_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_230_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_243_ _243_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_17_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_167_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput18 vssd2 _339_/A1 vccd1 io_in[25] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input80_A vssd2 vccd1 vccd1 vssd2 la_data_in[21] sky130_fd_sc_hd__diode_2
XFILLER_196_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_174_ _174_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
Xinput29 vssd2 input29/X vccd1 io_in[35] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_167_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_211_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xrepeater608 vssd2 _316_/A vccd1 _323_/A vccd1 vssd2 sky130_fd_sc_hd__buf_8
XFILLER_78_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_37 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_185_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_185_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_58_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_406 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_0_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_428 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_439 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_180_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput480 vssd2 la_data_out[17] vccd1 _161_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput491 vssd2 la_data_out[27] vccd1 _171_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input232_A vssd2 vccd1 vccd1 vssd2 la_oenb[43] sky130_fd_sc_hd__diode_2
XFILLER_208_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_170_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1749 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_103_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_242_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_940 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_973 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_984 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_156_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_460 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_15_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_226_ _226_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_129_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
X_157_ _157_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_144_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_088_ vssd2 _088_/Y vccd1 _352_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_170_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_adc.SCOMP_clk vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_228_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_0_1237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_178_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_120_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_89_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput208 vssd2 input208/X vccd1 la_oenb[21] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput219 vssd2 input219/X vccd1 la_oenb[31] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_130_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_170_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_186_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_231_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_0_1760 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_129_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_269 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input182_A vssd2 vccd1 vccd1 vssd2 la_oenb[113] sky130_fd_sc_hd__diode_2
XFILLER_119_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_3_134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input43_A vssd2 vccd1 vccd1 vssd2 la_data_in[103] sky130_fd_sc_hd__diode_2
XFILLER_216_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1509 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_108_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_770 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_781 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_209_ _209_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_15_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__093__B1 vssd2 vccd1 vccd1 vssd2 _074_/A sky130_fd_sc_hd__diode_2
XFILLER_238_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_916 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_65_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_213_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_adc.COMP_clk vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_80_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__336__A vssd2 vccd1 vccd1 vssd2 _336_/A sky130_fd_sc_hd__diode_2
XFILLER_61_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__071__A vssd2 vccd1 vccd1 vssd2 _356_/Q sky130_fd_sc_hd__diode_2
XFILLER_11_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__084__B1 vssd2 vccd1 vccd1 vssd2 _074_/X sky130_fd_sc_hd__diode_2
XFILLER_211_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1800 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_245_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1822 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_623 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_213_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_138_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_4_454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_671 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_188_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__090__A3 vssd2 vccd1 vccd1 vssd2 _073_/X sky130_fd_sc_hd__diode_2
XFILLER_90_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2019 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_78_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__081__A3 vssd2 vccd1 vccd1 vssd2 _073_/X sky130_fd_sc_hd__diode_2
XFILLER_82_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_165_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_895 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_148_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_102 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input145_A vssd2 vccd1 vccd1 vssd2 la_data_in[80] sky130_fd_sc_hd__diode_2
XFILLER_190_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA__057__B1 vssd2 vccd1 vccd1 vssd2 _356_/Q sky130_fd_sc_hd__diode_2
XFILLER_76_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2342 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input312_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[23] sky130_fd_sc_hd__diode_2
XFILLER_245_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_60_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1173 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_71_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_26_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_199_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_23 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_34 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_45 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_82_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_56 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_109_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_67 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_89 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_692 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
X_190_ _190_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_195_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_174_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input262_A vssd2 vccd1 vccd1 vssd2 la_oenb[70] sky130_fd_sc_hd__diode_2
XFILLER_123_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_213_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1181 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_12_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_141_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_83_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1944 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1991 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_11_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_8_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_42_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input108_A vssd2 vccd1 vccd1 vssd2 la_data_in[47] sky130_fd_sc_hd__diode_2
XFILLER_153_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_243_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_311_ vssd2 _311_/X vccd1 _314_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_204_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_242_ _242_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_22_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput19 vssd2 _339_/S vccd1 io_in[26] vccd1 vssd2 sky130_fd_sc_hd__buf_1
X_173_ _173_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input73_A vssd2 vccd1 vccd1 vssd2 la_data_in[15] sky130_fd_sc_hd__diode_2
XFILLER_170_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_238_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xrepeater609 vssd2 _323_/A vccd1 _326_/A vccd1 vssd2 sky130_fd_sc_hd__buf_8
XFILLER_78_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_20_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_49 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__355__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_87_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_51_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_407 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_418 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__074__A vssd2 vccd1 vccd1 vssd2 _074_/A sky130_fd_sc_hd__diode_2
XFILLER_140_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_20_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_149_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_509 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_164_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput470 vssd2 la_data_out[123] vccd1 _267_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_216_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_900 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput481 vssd2 la_data_out[18] vccd1 _162_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput492 vssd2 la_data_out[28] vccd1 _172_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_87_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input225_A vssd2 vccd1 vccd1 vssd2 la_oenb[37] sky130_fd_sc_hd__diode_2
XFILLER_210_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_179_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_106_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_941 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_952 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_8_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_985 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_30_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_225_ _225_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_15_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_156_ _156_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_087_ vssd2 _345_/D _074_/X _086_/X vccd1 _085_/Y _072_/A _073_/X vccd1 vssd2 sky130_fd_sc_hd__o311a_1
XFILLER_6_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_152_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_80_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_15_1950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput209 vssd2 input209/X vccd1 la_oenb[22] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_69_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1943 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__069__A vssd2 vccd1 vccd1 vssd2 _074_/A sky130_fd_sc_hd__diode_2
XFILLER_186_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_213_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_204 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_224_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_51_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_166_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input175_A vssd2 vccd1 vccd1 vssd2 la_oenb[107] sky130_fd_sc_hd__diode_2
XFILLER_238_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_175_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input342_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[20] sky130_fd_sc_hd__diode_2
XFILLER_160_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input36_A vssd2 vccd1 vccd1 vssd2 io_in[7] sky130_fd_sc_hd__diode_2
XFILLER_94_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2204 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_248_796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_112_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_74_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_186_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_235_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_223_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_760 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_88_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_782 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_793 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_208_ _208_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_139_ _139_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_116_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1002 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_928 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_0_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_148_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_635 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_2270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_668 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_60_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input292_A vssd2 vccd1 vccd1 vssd2 la_oenb[98] sky130_fd_sc_hd__diode_2
XFILLER_60_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_989 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_4_466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_1_2001 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_169_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_188_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_90_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_590 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_156_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_131_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__066__B vssd2 vccd1 vccd1 vssd2 _072_/A sky130_fd_sc_hd__diode_2
XFILLER_224_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__082__A vssd2 vccd1 vccd1 vssd2 _354_/Q sky130_fd_sc_hd__diode_2
XFILLER_135_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_213_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_76_215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__057__A1 vssd2 vccd1 vccd1 vssd2 _357_/Q sky130_fd_sc_hd__diode_2
XFILLER_213_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__057__B2 vssd2 vccd1 vccd1 vssd2 _056_/X sky130_fd_sc_hd__diode_2
XANTENNA_input138_A vssd2 vccd1 vccd1 vssd2 la_data_in[74] sky130_fd_sc_hd__diode_2
XFILLER_162_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_142 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_217_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input305_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[17] sky130_fd_sc_hd__diode_2
XFILLER_144_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1385 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_177_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_390 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1030 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1940 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_26_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_35 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_46 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_202_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_57 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_68 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_79 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_813 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input255_A vssd2 vccd1 vccd1 vssd2 la_oenb[64] sky130_fd_sc_hd__diode_2
XFILLER_235_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2147 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1193 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_108_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_188_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1956 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_310_ vssd2 _310_/X vccd1 _316_/A vccd1 vssd2 sky130_fd_sc_hd__clkbuf_1
XFILLER_242_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_610 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_241_ _241_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_52_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
X_172_ _172_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_52_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_88 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input66_A vssd2 vccd1 vccd1 vssd2 la_data_in[124] sky130_fd_sc_hd__diode_2
XFILLER_219_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_69_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_113_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_1943 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_224_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_419 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_145_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1929 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput460 vssd2 la_data_out[114] vccd1 _258_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
Xoutput471 vssd2 la_data_out[124] vccd1 _268_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput482 vssd2 la_data_out[19] vccd1 _163_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput493 vssd2 la_data_out[29] vccd1 _173_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_160_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_912 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XANTENNA_input120_A vssd2 vccd1 vccd1 vssd2 la_data_in[58] sky130_fd_sc_hd__diode_2
XFILLER_90_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input218_A vssd2 vccd1 vccd1 vssd2 la_oenb[30] sky130_fd_sc_hd__diode_2
XFILLER_216_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2243 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_920 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_931 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_106_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_953 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_964 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_224_ _224_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_7_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_155_ _155_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_144_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_13_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_13_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_086_ vssd2 _086_/X _345_/Q vccd1 _099_/A _099_/B _354_/Q vccd1 vssd2 sky130_fd_sc_hd__a31o_1
XFILLER_124_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_65_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1397 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_213_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_209_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_216 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_213_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__085__A vssd2 vccd1 vccd1 vssd2 _353_/Q sky130_fd_sc_hd__diode_2
XPHY_238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_147 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input168_A vssd2 vccd1 vccd1 vssd2 la_oenb[100] sky130_fd_sc_hd__diode_2
XFILLER_134_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input335_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[14] sky130_fd_sc_hd__diode_2
XFILLER_59_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input29_A vssd2 vccd1 vccd1 vssd2 io_in[35] sky130_fd_sc_hd__diode_2
XFILLER_21_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1673 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1515 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_74_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_75 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1559 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2040 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_188_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_761 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_772 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA__345__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XPHY_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_175_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_794 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_207_ _207_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_209_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_138_ _138_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_7_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_069_ vssd2 _069_/Y vccd1 _074_/A vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_99_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_98_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__093__A2 vssd2 vccd1 vccd1 vssd2 _072_/A sky130_fd_sc_hd__diode_2
XFILLER_130_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_235_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_502 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_116_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_629 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__084__A2 vssd2 vccd1 vccd1 vssd2 _104_/A sky130_fd_sc_hd__diode_2
XFILLER_84_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_647 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_246_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input285_A vssd2 vccd1 vccd1 vssd2 la_oenb[91] sky130_fd_sc_hd__diode_2
XFILLER_138_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_176_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_109_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_68_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_684 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_572 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_48_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_1492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_217_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_189_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_223_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_12_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1015 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_511 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_842 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__066__C vssd2 vccd1 vccd1 vssd2 _339_/X sky130_fd_sc_hd__diode_2
XFILLER_210_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_135_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_235_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__057__A2 vssd2 vccd1 vccd1 vssd2 _055_/X sky130_fd_sc_hd__diode_2
XFILLER_213_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input200_A vssd2 vccd1 vccd1 vssd2 la_oenb[14] sky130_fd_sc_hd__diode_2
XFILLER_44_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input96_A vssd2 vccd1 vccd1 vssd2 la_data_in[36] sky130_fd_sc_hd__diode_2
XFILLER_220_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_7_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_95_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_993 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_121_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput360 vssd2 input360/X vccd1 wbs_dat_i[8] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1407 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_40_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_188_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_91_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1128 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_220_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_167_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_187_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_14 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_1985 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_36 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_26_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_41_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_69 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_210_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input150_A vssd2 vccd1 vccd1 vssd2 la_data_in[85] sky130_fd_sc_hd__diode_2
XFILLER_238_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input248_A vssd2 vccd1 vccd1 vssd2 la_oenb[58] sky130_fd_sc_hd__diode_2
XFILLER_8_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_66_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input11_A vssd2 vccd1 vccd1 vssd2 io_in[19] sky130_fd_sc_hd__diode_2
XFILLER_189_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_2_2185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_61_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_148_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_2105 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_82_53 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_2138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_116_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_231_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_188_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput190 vssd2 input190/X vccd1 la_oenb[120] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_224_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_238_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_736 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_132_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input3_A vssd2 vccd1 vccd1 vssd2 io_in[11] sky130_fd_sc_hd__diode_2
XFILLER_87_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__088__A vssd2 vccd1 vccd1 vssd2 _352_/Q sky130_fd_sc_hd__diode_2
XFILLER_36_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_55_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_93_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_54_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1746 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_240_ _240_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_171_ _171_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_178_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1470 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input198_A vssd2 vccd1 vccd1 vssd2 la_oenb[12] sky130_fd_sc_hd__diode_2
XFILLER_13_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input365_A vssd2 vccd1 vccd1 vssd2 wbs_sel_i[3] sky130_fd_sc_hd__diode_2
XFILLER_109_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_521 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_112_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input59_A vssd2 vccd1 vccd1 vssd2 la_data_in[118] sky130_fd_sc_hd__diode_2
XFILLER_184_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output584_A vssd2 vccd1 vccd1 vssd2 _293_/LO sky130_fd_sc_hd__diode_2
XFILLER_202_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_142_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_95_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_243_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput450 vssd2 la_data_out[105] vccd1 _249_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_138_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput461 vssd2 la_data_out[115] vccd1 _259_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_160_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput472 vssd2 la_data_out[125] vccd1 _269_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput483 vssd2 la_data_out[1] vccd1 _145_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput494 vssd2 la_data_out[2] vccd1 _146_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_232_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_924 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_102_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1844 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1888 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input113_A vssd2 vccd1 vccd1 vssd2 la_data_in[51] sky130_fd_sc_hd__diode_2
XFILLER_19_2211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_2255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_932 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_943 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_106_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_965 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_204_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_976 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_223_ _223_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_223_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_154_ _154_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_7_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_085_ vssd2 _085_/Y vccd1 _353_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_13_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_38_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1028 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1074 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__096__B1 vssd2 vccd1 vccd1 vssd2 _074_/A sky130_fd_sc_hd__diode_2
XFILLER_9_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_168_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_37 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_80_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_217 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_213_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_228 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_205_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1727 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_3_126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_216_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__087__B1 vssd2 vccd1 vccd1 vssd2 _074_/X sky130_fd_sc_hd__diode_2
XFILLER_58_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input230_A vssd2 vccd1 vccd1 vssd2 la_oenb[41] sky130_fd_sc_hd__diode_2
XFILLER_247_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input328_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[9] sky130_fd_sc_hd__diode_2
XFILLER_74_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2052 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_70_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_231_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_773 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_196_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_206_ _206_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_128_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_183_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_137_ _137_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_239_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_7_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_068_ vssd2 _074_/A vccd1 _341_/Q vccd1 _076_/A vssd2 sky130_fd_sc_hd__or2_4
XFILLER_171_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__078__B1 vssd2 vccd1 vccd1 vssd2 _074_/X sky130_fd_sc_hd__diode_2
XFILLER_234_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__093__A3 vssd2 vccd1 vccd1 vssd2 _339_/X sky130_fd_sc_hd__diode_2
XFILLER_120_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1015 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_62 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_94_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__084__A3 vssd2 vccd1 vccd1 vssd2 _073_/X sky130_fd_sc_hd__diode_2
XFILLER_56_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_84_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1858 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_246_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2283 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_225_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1535 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_220_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1568 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input180_A vssd2 vccd1 vccd1 vssd2 la_oenb[111] sky130_fd_sc_hd__diode_2
XFILLER_10_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input278_A vssd2 vccd1 vccd1 vssd2 la_oenb[85] sky130_fd_sc_hd__diode_2
XFILLER_175_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_969 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_181_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input41_A vssd2 vccd1 vccd1 vssd2 la_data_in[101] sky130_fd_sc_hd__diode_2
XFILLER_216_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_570 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_31_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_157_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_repeater612_A vssd2 vccd1 vccd1 vssd2 input17/X sky130_fd_sc_hd__diode_2
XFILLER_12_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_38_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_187_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_214_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_62_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2133 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_416 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_118_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_22_2262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_84_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1655 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_2309 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_144_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_111_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_242_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input89_A vssd2 vccd1 vccd1 vssd2 la_data_in[2] sky130_fd_sc_hd__diode_2
XFILLER_16_1376 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_127_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_460 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_3_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_121_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput350 vssd2 input350/X vccd1 wbs_dat_i[28] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput361 vssd2 input361/X vccd1 wbs_dat_i[9] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_76_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1107 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1953 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_81_242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_765 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_26 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_37 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_35_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_81_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1917 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_13_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_117_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_8_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_686 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_238_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_77_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_62 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input143_A vssd2 vccd1 vccd1 vssd2 la_data_in[79] sky130_fd_sc_hd__diode_2
XFILLER_8_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input310_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[21] sky130_fd_sc_hd__diode_2
XFILLER_66_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1430 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_2117 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_202_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput180 vssd2 input180/X vccd1 la_oenb[111] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_236_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput191 vssd2 input191/X vccd1 la_oenb[121] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_36_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_63_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_24_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_224_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_23_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_99_673 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_629 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_35_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_51_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_170_ _170_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_178_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1482 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_178_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input260_A vssd2 vccd1 vccd1 vssd2 la_oenb[69] sky130_fd_sc_hd__diode_2
XFILLER_123_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input358_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[6] sky130_fd_sc_hd__diode_2
XFILLER_117_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_189_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1547 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output577_A vssd2 vccd1 vccd1 vssd2 _286_/LO sky130_fd_sc_hd__diode_2
XFILLER_174_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_299_ _299_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_139_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_9_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_138_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_2345 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_106_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_105_236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_9 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xoutput440 vssd2 io_out[6] vccd1 _123_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput451 vssd2 la_data_out[106] vccd1 _250_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput462 vssd2 la_data_out[116] vccd1 _260_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput473 vssd2 la_data_out[126] vccd1 _270_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput484 vssd2 la_data_out[20] vccd1 _164_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput495 vssd2 la_data_out[30] vccd1 _174_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_99_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__099__A vssd2 vccd1 vccd1 vssd2 _099_/A sky130_fd_sc_hd__diode_2
XFILLER_5_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_243_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_900 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input106_A vssd2 vccd1 vccd1 vssd2 la_data_in[45] sky130_fd_sc_hd__diode_2
XFILLER_231_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_93_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_145_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2109 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_944 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_106_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_431 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_208_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_51_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_977 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_222_ _222_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_204_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_153_ _153_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_17_1290 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input71_A vssd2 vccd1 vccd1 vssd2 la_data_in[13] sky130_fd_sc_hd__diode_2
X_084_ vssd2 _346_/D _074_/X _083_/X vccd1 _082_/Y _104_/A _073_/X vccd1 vssd2 sky130_fd_sc_hd__o311a_1
XFILLER_13_1176 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_113_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_120_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_228_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_124_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_239_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__096__A1 vssd2 vccd1 vccd1 vssd2 _100_/B sky130_fd_sc_hd__diode_2
XFILLER_233_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_244_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1706 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1739 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_102_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input223_A vssd2 vccd1 vccd1 vssd2 la_oenb[35] sky130_fd_sc_hd__diode_2
XFILLER_247_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_74_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_55 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_227_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_19_2064 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_730 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_741 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_203_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2097 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_774 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_208_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_76 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_785 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_205_ _205_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_7_411 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_23_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_139_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_136_ _136_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_183_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_143_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_394 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
X_067_ vssd2 _076_/A vccd1 _340_/Q vccd1 vssd2 sky130_fd_sc_hd__buf_2
XFILLER_136_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_98_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_193_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_94_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_52 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_169_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_96 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_179_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_62_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_48_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_131_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1815 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2072 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1798 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_197_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_125_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1124 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_109_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_125_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input173_A vssd2 vccd1 vccd1 vssd2 la_oenb[105] sky130_fd_sc_hd__diode_2
XFILLER_10_1157 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_27_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_133_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input340_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[19] sky130_fd_sc_hd__diode_2
XFILLER_23_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_121_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input34_A vssd2 vccd1 vccd1 vssd2 io_in[5] sky130_fd_sc_hd__diode_2
XFILLER_248_552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_76_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2059 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_582 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_145_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_119_ _119_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_125_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_39_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_241_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1812 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_194_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_202_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2145 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2178 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_39_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2274 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_58_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2012 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input290_A vssd2 vccd1 vccd1 vssd2 la_oenb[96] sky130_fd_sc_hd__diode_2
XFILLER_139_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_27_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput340 vssd2 input340/X vccd1 wbs_dat_i[19] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput351 vssd2 input351/X vccd1 wbs_dat_i[29] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput362 vssd2 input362/X vccd1 wbs_sel_i[0] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_236_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1166 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_129 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1119 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_390 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_160_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1000 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_100_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1055 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1965 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_16 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_81_254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_558 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_38 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_49 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_81_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_1620 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1506 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1539 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_190_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_117_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_74 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_8_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input136_A vssd2 vccd1 vccd1 vssd2 la_data_in[72] sky130_fd_sc_hd__diode_2
XFILLER_22_2071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_126 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input303_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[15] sky130_fd_sc_hd__diode_2
XFILLER_73_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_114_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_95_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput170 vssd2 input170/X vccd1 la_oenb[102] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput181 vssd2 input181/X vccd1 la_oenb[112] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1915 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput192 vssd2 input192/X vccd1 la_oenb[122] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_236_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_176_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput600 vssd2 wbs_dat_o[31] vccd1 _307_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_219_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_641 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_236_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_1034 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_160_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_99_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_228_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_51_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_460 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_196_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_668 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1461 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_156_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1347 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1071 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_545 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_117_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input253_A vssd2 vccd1 vccd1 vssd2 la_oenb[62] sky130_fd_sc_hd__diode_2
XFILLER_215_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_120_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1307 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__348__CLK vssd2 vccd1 vccd1 vssd2 wb_clk_i sky130_fd_sc_hd__diode_2
XFILLER_18_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_298_ _298_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_192_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1881 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_122_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1712 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1745 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_33_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_146_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput430 vssd2 io_out[31] vccd1 _343_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_172_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput441 vssd2 io_out[7] vccd1 _124_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput452 vssd2 la_data_out[107] vccd1 _251_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput463 vssd2 la_data_out[117] vccd1 _261_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput474 vssd2 la_data_out[127] vccd1 _271_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput485 vssd2 la_data_out[21] vccd1 _165_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput496 vssd2 la_data_out[31] vccd1 _175_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__099__B vssd2 vccd1 vccd1 vssd2 _099_/B sky130_fd_sc_hd__diode_2
XFILLER_102_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1802 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1570 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2202 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_901 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_912 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_2268 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_934 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_30_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_945 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_956 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_144_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_967 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_221_ _221_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_243_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_168_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_152_ _152_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_183_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_083_ vssd2 _083_/X _346_/Q vccd1 _099_/A _099_/B _355_/Q vccd1 vssd2 sky130_fd_sc_hd__a31o_1
XFILLER_197_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input64_A vssd2 vccd1 vccd1 vssd2 la_data_in[122] sky130_fd_sc_hd__diode_2
XFILLER_136_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_193_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_98_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1087 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_124_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1022 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_15_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA__096__A2 vssd2 vccd1 vccd1 vssd2 _339_/X sky130_fd_sc_hd__diode_2
XFILLER_25_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2333 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1914 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_74 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_20_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1430 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_197_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1798 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_33_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1718 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_149_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_137_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__087__A2 vssd2 vccd1 vccd1 vssd2 _072_/A sky130_fd_sc_hd__diode_2
XFILLER_181_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_229_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_60_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_147_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1529 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input216_A vssd2 vccd1 vccd1 vssd2 la_oenb[29] sky130_fd_sc_hd__diode_2
XFILLER_28_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_720 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_2076 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_753 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_775 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_786 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_204_ _204_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_90_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_135_ _135_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_183_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_066_ vssd2 _066_/X vccd1 _066_/A vccd1 _072_/A vssd2 _339_/X sky130_fd_sc_hd__or3_4
XFILLER_178_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__078__A2 vssd2 vccd1 vccd1 vssd2 _104_/A sky130_fd_sc_hd__diode_2
XFILLER_31_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_151_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output435_A vssd2 vccd1 vccd1 vssd2 _348_/Q sky130_fd_sc_hd__diode_2
XFILLER_78_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_66_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_94_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_207_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_203_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_233_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_111_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_2084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_183_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_55_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_240_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_14_1250 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_822 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1136 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_175_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1169 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input166_A vssd2 vccd1 vccd1 vssd2 la_data_in[9] sky130_fd_sc_hd__diode_2
XFILLER_133_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_62_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_235_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input333_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[12] sky130_fd_sc_hd__diode_2
XFILLER_121_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input27_A vssd2 vccd1 vccd1 vssd2 io_in[33] sky130_fd_sc_hd__diode_2
XFILLER_1_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_5_2185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_76_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1484 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1326 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_182_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_34_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1014 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_572 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_157_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_118_ _118_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_12_1979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_993 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_98_536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_234_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_38_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_34_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1824 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_143_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_58_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_73_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_36 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_2024 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2046 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1063 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_154_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input283_A vssd2 vccd1 vccd1 vssd2 la_oenb[8] sky130_fd_sc_hd__diode_2
XFILLER_139_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1091 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_45_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_150_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput330 vssd2 input330/X vccd1 wbs_dat_i[0] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_96_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput341 vssd2 input341/X vccd1 wbs_dat_i[1] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_88_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput352 vssd2 input352/X vccd1 wbs_dat_i[2] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_29_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput363 vssd2 input363/X vccd1 wbs_sel_i[1] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_222_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_91_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_1873 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_242_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_59_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_167_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_55_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1067 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_55_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1977 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XPHY_17 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_28 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_63_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_81_266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_91_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2073 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1632 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_41_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1665 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_399 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1518 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1698 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1242 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_117_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_217_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input129_A vssd2 vccd1 vccd1 vssd2 la_data_in[66] sky130_fd_sc_hd__diode_2
XFILLER_122_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_138 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2199 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_73_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input94_A vssd2 vccd1 vccd1 vssd2 la_data_in[34] sky130_fd_sc_hd__diode_2
XFILLER_186_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_217_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput160 vssd2 input160/X vccd1 la_data_in[94] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput171 vssd2 input171/X vccd1 la_oenb[103] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput182 vssd2 input182/X vccd1 la_oenb[113] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput193 vssd2 input193/X vccd1 la_oenb[123] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1973 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_108_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput601 vssd2 wbs_dat_o[3] vccd1 _279_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_172_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_100_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_95_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_494 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1050 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1083 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_28_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input246_A vssd2 vccd1 vccd1 vssd2 la_oenb[56] sky130_fd_sc_hd__diode_2
XFILLER_115_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_59_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_92_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1319 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1214 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_18_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1226 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1821 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_1854 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_297_ _297_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_200_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_1893 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_154_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_17 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_77_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1724 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1914 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_20_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1757 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1770 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2060 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput420 vssd2 io_out[22] vccd1 _139_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput431 vssd2 io_out[32] vccd1 _344_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput442 vssd2 io_out[8] vccd1 _125_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput453 vssd2 la_data_out[108] vccd1 _252_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput464 vssd2 la_data_out[118] vccd1 _262_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput475 vssd2 la_data_out[12] vccd1 _156_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput486 vssd2 la_data_out[22] vccd1 _166_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput497 vssd2 la_data_out[32] vccd1 _176_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input1_A vssd2 vccd1 vccd1 vssd2 io_in[0] sky130_fd_sc_hd__diode_2
XFILLER_210_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_102_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_74_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_227_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_43 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_63_47 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_187_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_247_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_924 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_179_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_221_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_11_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_957 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_220_ _220_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XPHY_968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_979 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_151_ _151_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_168_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input196_A vssd2 vccd1 vccd1 vssd2 la_oenb[126] sky130_fd_sc_hd__diode_2
XFILLER_155_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_082_ vssd2 _082_/Y vccd1 _354_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_183_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_178_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input363_A vssd2 vccd1 vccd1 vssd2 wbs_sel_i[1] sky130_fd_sc_hd__diode_2
XFILLER_136_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input57_A vssd2 vccd1 vccd1 vssd2 la_data_in[116] sky130_fd_sc_hd__diode_2
XFILLER_151_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2036 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_59_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_659 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_207_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_209_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1099 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_226_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_124_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_349_ _349_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _349_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_204_1662 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1695 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_239_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_671 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_128_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_103_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__096__A3 vssd2 vccd1 vccd1 vssd2 _104_/A sky130_fd_sc_hd__diode_2
XFILLER_111_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_2200 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_96_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_37_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1521 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_92_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1777 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_244_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1442 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1426 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1421 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1454 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1318 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__087__A3 vssd2 vccd1 vccd1 vssd2 _073_/X sky130_fd_sc_hd__diode_2
XFILLER_88_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1611 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_779 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_182_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input111_A vssd2 vccd1 vccd1 vssd2 la_data_in[4] sky130_fd_sc_hd__diode_2
Xadc.COMP analog_io[1] analog_io[0] _337_/A vccd2 vssd2 wb_clk_i vccd2 vssd2 ACMP
XANTENNA_input209_A vssd2 vccd1 vccd1 vssd2 la_oenb[22] sky130_fd_sc_hd__diode_2
XFILLER_82_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_43_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_732 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_743 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_2088 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_56 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_157_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_765 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_11_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_787 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_180_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_203_ _203_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XPHY_798 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_274 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_998 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_475 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_134_ _134_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_23_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_065_ vssd2 _072_/A vccd1 _065_/A vccd1 vssd2 sky130_fd_sc_hd__buf_2
XFILLER_234_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_151_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_155_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA__078__A3 vssd2 vccd1 vccd1 vssd2 _073_/X sky130_fd_sc_hd__diode_2
XFILLER_78_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_163_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_200_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_115_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_183_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_94_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_556 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_342 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_183_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_212_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_504 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1574 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1267 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1262 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_147_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_834 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1148 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input159_A vssd2 vccd1 vccd1 vssd2 la_data_in[93] sky130_fd_sc_hd__diode_2
XFILLER_0_655 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_88_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_212_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input326_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[7] sky130_fd_sc_hd__diode_2
XFILLER_236_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_2197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_673 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_34_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_19_1140 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1946 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_551 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_573 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_240_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_242_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1026 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_200_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.SCOMP_INN vssd2 vccd1 vccd1 vssd2 analog_io[5] sky130_fd_sc_hd__diode_2
XPHY_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_129_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_117_ _117_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_193_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_10_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_121_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_46_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_241_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_813 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1803 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_2277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_17_1836 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1869 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_2340 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1413 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_537 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_218_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_48 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2008 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1371 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_2003 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_246_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2058 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_179_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1075 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_154_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input276_A vssd2 vccd1 vccd1 vssd2 la_oenb[83] sky130_fd_sc_hd__diode_2
XFILLER_194_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_107_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_150_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_452 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_96_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput320 vssd2 input320/X vccd1 wbs_adr_i[30] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput331 vssd2 input331/X vccd1 wbs_dat_i[10] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_48_423 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput342 vssd2 input342/X vccd1 wbs_dat_i[20] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_96_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput353 vssd2 input353/X vccd1 wbs_dat_i[30] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_75_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput364 vssd2 input364/X vccd1 wbs_sel_i[2] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_29_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_36_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_29_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_90_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_28_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_73_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_370 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_176_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_adc.COMP_INN vssd2 vccd1 vccd1 vssd2 analog_io[1] sky130_fd_sc_hd__diode_2
XFILLER_8_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_repeater610_A vssd2 vccd1 vccd1 vssd2 _331_/A sky130_fd_sc_hd__diode_2
XFILLER_144_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1490 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1079 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_55_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_18 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_29 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_247_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_50_610 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_91_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_104_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_225_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1677 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1221 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_24_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_106_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_8_1889 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_618 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_245_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_2156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_6_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1422 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_233_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_218_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_96_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1488 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_158_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input87_A vssd2 vccd1 vccd1 vssd2 la_data_in[28] sky130_fd_sc_hd__diode_2
XFILLER_194_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_31_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__102__A vssd2 vccd1 vccd1 vssd2 _353_/Q sky130_fd_sc_hd__diode_2
XFILLER_122_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput150 vssd2 input150/X vccd1 la_data_in[85] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput161 vssd2 input161/X vccd1 la_data_in[95] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput172 vssd2 input172/X vccd1 la_oenb[104] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput183 vssd2 input183/X vccd1 la_oenb[114] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput194 vssd2 input194/X vccd1 la_oenb[124] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1952 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1985 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_203_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2231 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_118_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2264 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2297 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput602 vssd2 wbs_dat_o[4] vccd1 _280_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_215_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_36_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_357 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_243_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1170 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1062 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_123_217 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1095 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_232_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input141_A vssd2 vccd1 vccd1 vssd2 la_data_in[77] sky130_fd_sc_hd__diode_2
XFILLER_232_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input239_A vssd2 vccd1 vccd1 vssd2 la_oenb[4] sky130_fd_sc_hd__diode_2
XFILLER_98_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_12 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_459 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_248_1248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_27_971 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1285 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1205 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1238 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1833 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1866 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_296_ _296_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_201_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_157_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_111_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1005 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1736 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_225_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_92_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_248_1782 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1914 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_2191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_165_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1625 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_691 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_118_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_146_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput410 vssd2 io_out[13] vccd1 _130_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput421 vssd2 io_out[23] vccd1 _140_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput432 vssd2 io_out[33] vccd1 _345_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput443 vssd2 io_out[9] vccd1 _126_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput454 vssd2 la_data_out[109] vccd1 _253_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput465 vssd2 la_data_out[119] vccd1 _263_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput476 vssd2 la_data_out[13] vccd1 _157_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput487 vssd2 la_data_out[23] vccd1 _167_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput498 vssd2 la_data_out[33] vccd1 _177_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_214_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1859 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_110_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_903 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_914 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_936 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_70_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_23_451 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_958 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_221_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_969 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_243_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_646 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_150_ _150_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_10_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_489 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_195_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_081_ vssd2 _347_/D _074_/X _080_/X vccd1 _079_/Y _104_/A _073_/X vccd1 vssd2 sky130_fd_sc_hd__o311a_1
XFILLER_148_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input189_A vssd2 vccd1 vccd1 vssd2 la_oenb[11] sky130_fd_sc_hd__diode_2
XFILLER_128_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input356_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[4] sky130_fd_sc_hd__diode_2
XFILLER_191_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_151_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2162 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2195 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_2048 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_649 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_207_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1045 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_1082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_222_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1057 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_348_ _348_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _348_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_180_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1674 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_279_ _279_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_155_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_128_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_183_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_143_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_1938 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_168_2234 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1533 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_209_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1789 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1405 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1438 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1580 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_177_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1433 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_88_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_137_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_14_1466 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_49_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_58_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_25_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_21_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2081 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_56_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_130_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1311 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_700 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XANTENNA_input104_A vssd2 vccd1 vccd1 vssd2 la_data_in[43] sky130_fd_sc_hd__diode_2
XPHY_711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_722 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_744 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_755 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_230_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_777 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_202_ _202_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_32_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_432 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_23_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_157_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
X_133_ _133_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_201_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_11_487 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_139_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_193_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_064_ vssd2 _066_/A vccd1 _357_/Q vccd1 vssd2 sky130_fd_sc_hd__inv_2
XFILLER_165_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1820 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_125_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1853 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_97_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_65_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_565 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_228_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_44 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_88 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_185_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_174_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_31_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_119_139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_239_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_7_992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_127_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_192_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_135_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_130_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1434 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_135_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1467 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2031 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1829 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_244_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1330 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_53_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2254 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_187_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_321 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_64_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_52_354 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_2207 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1586 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_516 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_142_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_139_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1279 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_119_640 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_406 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_147_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_846 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_25 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_107_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_194_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_153_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_197_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input221_A vssd2 vccd1 vccd1 vssd2 la_oenb[33] sky130_fd_sc_hd__diode_2
XFILLER_1_1306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_63_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input319_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[2] sky130_fd_sc_hd__diode_2
XFILLER_244_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_188_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_73_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_71_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_530 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_160_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_541 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1152 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1958 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_563 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_574 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_585 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1185 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_156_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_596 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1038 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1780 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_197_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_200_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_116_ _116_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_197_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1661 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_4_962 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_180_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_80_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_315 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1694 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_234_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_2289 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1848 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_2352 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1425 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_162_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_226_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_549 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_22_2233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1532 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_2_1615 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1626 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_0_2051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_226_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_53_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_198_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1383 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_201 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_481 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input171_A vssd2 vccd1 vccd1 vssd2 la_oenb[103] sky130_fd_sc_hd__diode_2
XFILLER_107_676 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input269_A vssd2 vccd1 vccd1 vssd2 la_oenb[77] sky130_fd_sc_hd__diode_2
XFILLER_136_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1039 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_431 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_122_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_110_819 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_153_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput310 vssd2 input310/X vccd1 wbs_adr_i[21] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_150_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput321 vssd2 input321/X vccd1 wbs_adr_i[31] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_96_78 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input32_A vssd2 vccd1 vccd1 vssd2 io_in[3] sky130_fd_sc_hd__diode_2
XFILLER_216_1194 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput332 vssd2 input332/X vccd1 wbs_dat_i[11] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput343 vssd2 input343/X vccd1 wbs_dat_i[21] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_188_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_1047 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xinput354 vssd2 input354/X vccd1 wbs_dat_i[31] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_0_497 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_48_435 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput365 vssd2 input365/X vccd1 wbs_sel_i[3] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_29_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1261 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_182_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_229_1588 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_164_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_43_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_71_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_125_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_371 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_84_7 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_382 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_242_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_393 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output488_A vssd2 vccd1 vccd1 vssd2 _168_/LO sky130_fd_sc_hd__diode_2
XFILLER_61_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_201_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_84_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_173_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_112_123 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1540 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_156 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_79_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1581 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_67_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_19 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_63_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_63_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1809 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_91_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1341 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_510 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_543 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1227 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_1689 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_429 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_129_790 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_237_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_219_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1266 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_624 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_173_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1312 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_132_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_66_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2030 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_106_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_1401 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_57_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_72_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_630 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_663 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1409 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_198_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_16_1100 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_534 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_154_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_589 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_235_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__102__B vssd2 vccd1 vccd1 vssd2 _352_/Q sky130_fd_sc_hd__diode_2
XFILLER_7_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput140 vssd2 input140/X vccd1 la_data_in[76] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_7_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_171 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
Xinput151 vssd2 input151/X vccd1 la_data_in[86] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput162 vssd2 input162/X vccd1 la_data_in[96] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_237_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput173 vssd2 input173/X vccd1 la_oenb[105] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_64_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput184 vssd2 input184/X vccd1 la_oenb[115] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_229_2020 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput195 vssd2 input195/X vccd1 la_oenb[125] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_40_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_229_2053 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_52_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1964 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1997 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_44_471 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_60_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1910 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_2215 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_2248 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_32_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_852 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_705 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_75_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_738 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2276 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput603 vssd2 wbs_dat_o[5] vccd1 _281_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_82_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_933 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_2322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_966 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_114_999 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_210_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1381 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_208_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_199_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_247_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_23_622 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1485 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_17_2121 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1617 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_196_914 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_223_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_17_2154 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_167_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_17 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_1182 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_351 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_384 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_202_1068 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_237 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_191_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_2_515 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_123_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_270 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_1735 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1768 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_465 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1890 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_77_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1120 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1776 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1153 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input134_A vssd2 vccd1 vccd1 vssd2 la_data_in[70] sky130_fd_sc_hd__diode_2
XFILLER_98_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_24 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_33_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input301_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[13] sky130_fd_sc_hd__diode_2
XFILLER_226_1503 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_27_983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1536 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_35_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1569 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_161_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_243_1861 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_699 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_35_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_243_1894 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1845 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_1113 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_295_ _295_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_155_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_1878 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_166_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_181_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1621 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_771 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1654 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1507 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_81_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1930 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_42_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1963 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_77 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_1816 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_1996 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_211_1849 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_1028 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_7_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1905 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_64_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_24_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_92_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_1877 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_248_1794 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_181_1926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_1609 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2061 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_149_115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1751 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2094 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1923 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1604 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_18_1784 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_203_2089 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1637 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_670 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_145_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_693 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_579 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput400 vssd2 io_oeb[4] vccd1 _111_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput411 vssd2 io_out[14] vccd1 _131_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput422 vssd2 io_out[24] vccd1 _141_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_229 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_86_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_538 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_161_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput433 vssd2 io_out[34] vccd1 _346_/Q vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput444 vssd2 la_data_out[0] vccd1 _144_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput455 vssd2 la_data_out[10] vccd1 _154_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
Xoutput466 vssd2 la_data_out[11] vccd1 _155_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_214_2130 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput477 vssd2 la_data_out[14] vccd1 _158_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_240 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xoutput488 vssd2 la_data_out[24] vccd1 _168_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_234_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xoutput499 vssd2 la_data_out[34] vccd1 _178_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_141_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_929 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2016 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_214_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_1974 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_210_2049 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_86_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1608 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2252 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2274 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_227_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_3_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_242_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_915 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_106_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_926 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_169_925 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_402 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_221_2101 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_225_2281 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_24_986 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_948 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_23_463 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_221_2134 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_221_2167 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_658 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_080_ vssd2 _080_/X _347_/Q vccd1 _099_/A _099_/B _356_/Q vccd1 vssd2 sky130_fd_sc_hd__a31o_1
XFILLER_10_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_192 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_128_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_178_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_13 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_178_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XANTENNA_input251_A vssd2 vccd1 vccd1 vssd2 la_oenb[60] sky130_fd_sc_hd__diode_2
XFILLER_151_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input349_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[27] sky130_fd_sc_hd__diode_2
XFILLER_191_1576 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_8_2174 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_78_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_703 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_93_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_1057 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_74_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_215_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_2310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_159_424 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1377 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_1006 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_457 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1069 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_347_ _347_/Q vssd2 wb_clk_i vccd1 vccd1 vssd2 _347_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_147_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_169_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_1992 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_278_ _278_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_13_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_127_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_651 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_115_505 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_170_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_143_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_172 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_237_1462 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1605 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1495 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_123_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_1007 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_233_1348 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1638 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_111_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_68_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_96_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_111_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_83_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2246 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_37_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_1702 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_2292 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1108 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_374 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1567 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_209_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_248_1591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_181_1723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_212_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1455 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_391 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1417 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_222_1731 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_220_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_2263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_811 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1592 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1764 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_203_1141 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_2247 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_1797 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1478 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1524 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_64_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_39 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_88_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_2275 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_99_2332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1882 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_101_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1657 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_612 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_56_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1449 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_114_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1918 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_2093 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_204_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_56_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_701 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_130_54 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1323 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_712 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_723 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_734 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_212_840 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_733 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_745 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_130_87 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_1356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_2251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_142_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_756 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_767 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
X_201_ _201_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_15_1209 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_169_766 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_32_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_789 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_184_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_619 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1951 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_444 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_169_799 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_132_ _132_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_201_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input299_A vssd2 vccd1 vccd1 vssd2 wbs_adr_i[11] sky130_fd_sc_hd__diode_2
XFILLER_109_310 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_172_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_499 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_343 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
X_063_ vssd2 _350_/D _350_/Q vccd1 _341_/Q _351_/Q _055_/A vccd1 vssd2 sky130_fd_sc_hd__a22o_1
XFILLER_152_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_165_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1832 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_180_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_847 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input62_A vssd2 vccd1 vccd1 vssd2 la_data_in[120] sky130_fd_sc_hd__diode_2
XFILLER_10_1865 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_643 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_155_51 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_234_2358 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_97_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_10_1898 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_3_687 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_105_571 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_2320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_2082 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1911 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_4_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_65_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_228_2118 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_544 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1950 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_577 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_206_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_21_1983 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_46_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_185_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_61_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_2329 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_204_2151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1710 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2203 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_159_298 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_200_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_13_2190 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_127_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_127_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_155_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_492 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_89_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_192_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_103_508 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_379 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_174_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_2122 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1446 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_85_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_6_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1189 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_57_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1479 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_2043 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xadc.DAC adc.DAC/d0 adc.DAC/d1 input15/X input14/X input13/X input11/X input10/X adc.DAC/x2_out_v
+ adc.DAC/x1_out_v analog_io[3] input9/X analog_io[2] adc.DAC/x2_vref1 adc.DAC/x1_vref5
+ vssd2 adc.DAC/inp2 vccd2 DAC_8BIT
XFILLER_20_2150 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1769 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2233 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_226_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_2183 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_168_1364 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_37_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_52_366 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_16_2219 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_40_528 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_244_1263 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_1296 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_1597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1149 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_220_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_652 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_134_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_685 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_147_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_238_1023 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_238_1056 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_69_37 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_613 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_115_880 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1332 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_2111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_9_2280 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_523 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_1365 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_48_606 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_87_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1218 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_0_679 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_216_1398 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_233_1690 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_1980 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_47_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_58 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_420 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_141_31 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_1498 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XANTENNA_input214_A vssd2 vccd1 vccd1 vssd2 la_oenb[27] sky130_fd_sc_hd__diode_2
XFILLER_244_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_186_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_216_453 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_28_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_1759 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_245_1027 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_244_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_486 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_648 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_160_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1450 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_54_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_520 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_71_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1303 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XPHY_531 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_227_1483 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_542 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_160_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_553 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_564 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1164 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_1336 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_681 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_575 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_586 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_19_1197 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_1369 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_597 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_156_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1650 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.SCOMP_INP vssd2 vccd1 vccd1 vssd2 analog_io[4] sky130_fd_sc_hd__diode_2
XFILLER_200_876 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_1792 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_240_1683 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
X_115_ _115_/LO vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__conb_1
XFILLER_197_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_158_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_144_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_109_151 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_83 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_193_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_109_184 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_137_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_236_1719 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1410 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_80_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_171_1711 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_327 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_output433_A vssd2 vccd1 vccd1 vssd2 _346_/Q sky130_fd_sc_hd__diode_2
XFILLER_67_904 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_140_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_71 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_6 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_67_937 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1752 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_78_2235 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_39_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1804 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_93_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_247_1837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_19_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1841 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_21_1791 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_62_653 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_1_1885 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_234_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_50_837 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_206_1512 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_714 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_30_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_136_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_30_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_961 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_11_1404 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_15_1584 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2044 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_176_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_600 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_129_994 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1437 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_239_2077 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_219_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_196_1092 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_828 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_170_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_69_241 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_130_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_84_211 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_2245 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_436 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_29_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1763 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_246_2004 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_469 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_85_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2305 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_1796 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1566 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_2308 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2030 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_246_2037 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2338 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_168_1161 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_412 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__080__B1 vssd2 vccd1 vccd1 vssd2 _347_/Q sky130_fd_sc_hd__diode_2
XFILLER_53_664 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_0_2096 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_198_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2346 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_607 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_53_697 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_71_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_222_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_27 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_138_213 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_119_493 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_218_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_175_1132 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_136_42 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_1788 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1165 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input164_A vssd2 vccd1 vccd1 vssd2 la_data_in[98] sky130_fd_sc_hd__diode_2
XFILLER_231_2317 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1018 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_175_1198 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_248_320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput300 vssd2 input300/X vccd1 wbs_adr_i[12] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput311 vssd2 input311/X vccd1 wbs_adr_i[22] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_7_1527 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput322 vssd2 input322/X vccd1 wbs_adr_i[3] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_0_476 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
Xinput333 vssd2 input333/X vccd1 wbs_dat_i[12] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input331_A vssd2 vccd1 vccd1 vssd2 wbs_dat_i[10] sky130_fd_sc_hd__diode_2
Xinput344 vssd2 input344/X vccd1 wbs_dat_i[22] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_49_959 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_152_30 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput355 vssd2 input355/X vccd1 wbs_dat_i[3] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_48_447 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput366 vssd2 input366/X vccd1 wbs_stb_i vccd1 vssd2 sky130_fd_sc_hd__buf_1
XANTENNA_input25_A vssd2 vccd1 vccd1 vssd2 io_in[31] sky130_fd_sc_hd__diode_2
XFILLER_229_2224 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1548 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_970 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_75_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_5_1273 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1115 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_205_913 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_90_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_44_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_1_1159 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_90_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_216_294 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_1125 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_44_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_94 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_43_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_164_2271 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_188_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_125_2244 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_188_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_1291 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_231_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_350 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_201_2110 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_372 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_383 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_125_2299 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_12_561 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_394 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_223_1177 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1633 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_118_909 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_61_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_594 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1666 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_184_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_240_1491 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_195_1519 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_82 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_adc.COMP_INP vssd2 vccd1 vccd1 vssd2 analog_io[0] sky130_fd_sc_hd__diode_2
XFILLER_184_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1210 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_1975 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_6_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_70 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_180_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_152_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_135 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_234_1251 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_550 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1552 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_112_168 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_140_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_230_1104 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_132_2259 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_234_1284 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_79_583 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_1137 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_227_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1560 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_67_778 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_82_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_1593 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_762 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_184_1902 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_81_236 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_228_1011 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_212_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1645 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_223_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_208_795 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA__062__B1 vssd2 vccd1 vccd1 vssd2 _351_/Q sky130_fd_sc_hd__diode_2
XFILLER_184_1935 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1660 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_212_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2232 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_247_1678 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_182_2360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_184_1968 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_223_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_1_1682 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_17_2325 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_50_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_143_2344 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_6
XFILLER_206_1320 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_91_2287 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_211_949 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_204_990 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_195_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1222 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_2328 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_206_1353 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_225_1987 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_148_522 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_1255 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1206 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_148_555 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_202_1239 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_408 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_163_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_15_1392 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_176_2175 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_116_441 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_151_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_2_708 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_191_1906 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_11_1278 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_219_1747 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_131_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_144_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_191_1939 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_104_636 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2304 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_63_2356 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_104_669 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_132_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_44_1010 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_150_2337 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_232_1947 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_1324 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_97_380 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_230_2361 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_22_2042 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_100_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_187_2260 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_57_277 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_100_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_245_367 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_22_1363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_225 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_187_2293 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_38_480 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2146 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_26_642 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_15 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_66 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_72_258 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_226_1707 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_26_675 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_99 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_183_2179 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_601 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_25_163 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_82_59 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_241_562 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_213_253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_41_634 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2316 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_213_286 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_198_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_241_595 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_70_2349 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_224_2187 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_16_1112 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_448 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_185_127 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_40_188 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_202_1740 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_363 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_194_2220 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XANTENNA_input281_A vssd2 vccd1 vccd1 vssd2 la_oenb[88] sky130_fd_sc_hd__diode_2
XFILLER_68_2223 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_322 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_166_396 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_120_2196 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_108_942 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_194_2253 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_5_546 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_126_249 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_190_2106 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_181_355 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_237_1825 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_190_2139 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_134_282 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_591 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_235_2272 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_96_807 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_122_477 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_231_2158 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_89_892 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_7_1335 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput130 vssd2 input130/X vccd1 la_data_in[67] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput141 vssd2 input141/X vccd1 la_data_in[77] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_237_835 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_209_526 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput152 vssd2 input152/X vccd1 la_data_in[87] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_7_1368 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput163 vssd2 input163/X vccd1 la_data_in[97] vccd1 vssd2 sky130_fd_sc_hd__buf_1
Xinput174 vssd2 input174/X vccd1 la_oenb[106] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_237_868 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput185 vssd2 input185/X vccd1 la_oenb[116] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_64_726 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
Xinput196 vssd2 input196/X vccd1 la_oenb[126] vccd1 vssd2 sky130_fd_sc_hd__buf_1
XFILLER_229_2032 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_229_2065 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_188_1389 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_205_721 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_189_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_162_2208 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_205_754 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_186_1080 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_921 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_45_995 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_60_954 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1922 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_242_2265 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_177_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_18_1955 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_14_1808 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XPHY_180 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XPHY_191 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_3
XFILLER_158_864 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_201_982 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_823 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_145_514 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_158_897 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_199_1474 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_68_3 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_173_856 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_12_2288 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_236_2025 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_133_709 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
Xoutput604 vssd2 wbs_dat_o[6] vccd1 _282_/LO vccd1 vssd2 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_750 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_113_400 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_126_783 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2301 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_193_1051 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_111 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_141_742 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_214_2334 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_193_1084 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_98_144 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_154_1035 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_4
XFILLER_114_978 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_86_306 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_101_628 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
XFILLER_171_1360 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_8
XFILLER_86_339 vssd2 vccd1 vccd1 vssd2 sky130_fd_sc_hd__decap_12
.ends

