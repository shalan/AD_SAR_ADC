magic
tech sky130A
magscale 1 2
timestamp 1626450099
<< checkpaint >>
rect -1520 -25390 20976 25102
<< locali >>
rect 302 23654 358 23734
rect 16410 13092 19408 13156
rect 19358 13050 19408 13092
rect 13744 12924 13862 13024
rect 13744 6592 13790 12924
rect 19358 12682 19412 13050
rect 19358 11948 19420 12682
rect 19358 11592 19424 11948
rect 19358 11198 19416 11592
rect 19358 10832 19420 11198
rect 19358 10068 19416 10832
rect 19358 9674 19412 10068
rect 19358 9330 19424 9674
rect 19358 8946 19416 9330
rect 19358 7038 19412 8946
rect 19366 6664 19420 7038
rect 13728 6575 13810 6592
rect 13728 6541 13754 6575
rect 13788 6541 13810 6575
rect 13728 6522 13810 6541
rect 10752 6176 11058 6318
rect 13738 6190 13820 6208
rect 10752 6172 10932 6176
rect 10752 4848 10844 6172
rect 13738 6156 13759 6190
rect 13793 6156 13820 6190
rect 13738 6138 13820 6156
rect 10770 4804 10844 4848
rect 10770 4018 10848 4804
rect 10770 3984 10805 4018
rect 10839 3984 10848 4018
rect 10770 3946 10848 3984
rect 7328 3404 7468 3486
rect 7330 3272 7460 3404
rect 10776 3312 10854 3374
rect 10776 3278 10787 3312
rect 10821 3278 10854 3312
rect 7326 2298 7464 3272
rect 7326 2264 7374 2298
rect 7408 2264 7464 2298
rect 7326 2226 7464 2264
rect 10776 3004 10854 3278
rect 3862 1257 3936 1772
rect 10776 1562 10848 3004
rect 3862 1223 3883 1257
rect 3917 1223 3936 1257
rect 3862 1194 3936 1223
rect 7348 1450 7464 1544
rect 7348 1416 7388 1450
rect 7422 1416 7464 1450
rect 806 531 864 904
rect 806 497 821 531
rect 855 497 864 531
rect 806 486 864 497
rect 3862 799 3946 828
rect 3862 765 3881 799
rect 3915 765 3946 799
rect 806 327 864 342
rect 806 293 816 327
rect 850 293 864 327
rect 10 -112 80 20
rect -244 -180 80 -112
rect 10 -182 80 -180
rect 806 -174 864 293
rect 806 -208 817 -174
rect 851 -208 864 -174
rect 806 -216 864 -208
rect -70 -450 258 -386
rect 3862 -437 3946 765
rect 804 -494 862 -466
rect 804 -528 817 -494
rect 851 -528 862 -494
rect 3862 -471 3893 -437
rect 3927 -471 3946 -437
rect 3862 -528 3946 -471
rect 7348 -278 7464 1416
rect 10776 696 10854 1562
rect 10776 -14 10856 696
rect 10774 -56 10856 -14
rect 804 -1038 862 -528
rect 3862 -955 3946 -916
rect 3862 -989 3883 -955
rect 3917 -989 3946 -955
rect 3862 -1558 3946 -989
rect 7348 -1044 7486 -278
rect 7348 -1078 7412 -1044
rect 7446 -1078 7486 -1044
rect 7348 -1120 7486 -1078
rect 7368 -1648 7486 -1600
rect 7368 -1682 7414 -1648
rect 7448 -1682 7486 -1648
rect 7368 -2730 7486 -1682
rect 10772 -2194 10856 -56
rect 10772 -2228 10795 -2194
rect 10829 -2228 10856 -2194
rect 10772 -2256 10856 -2228
rect 10780 -2748 10858 -2740
rect 10780 -2816 10864 -2748
rect 10780 -2850 10809 -2816
rect 10843 -2850 10864 -2816
rect 10780 -5774 10864 -2850
rect 13748 -4448 13794 6138
rect 19366 5536 19416 6664
rect 19366 5142 19412 5536
rect 19366 4764 19416 5142
rect 19366 4404 19420 4764
rect 19366 3356 19424 4404
rect 19366 2962 19412 3356
rect 19366 2244 19420 2962
rect 19366 1880 19416 2244
rect 19366 1188 19412 1880
rect 19358 1106 19412 1188
rect 19358 794 19408 1106
rect 19550 506 19716 518
rect 19550 472 19559 506
rect 19593 472 19716 506
rect 19550 456 19716 472
rect 17108 300 17190 392
rect 19422 -20 19532 42
rect 13752 -4700 13792 -4448
rect 13750 -4712 13792 -4700
rect 13750 -4994 13790 -4712
rect 13748 -5006 13790 -4994
rect 13748 -5530 13788 -5006
rect 13734 -5552 13812 -5530
rect 13734 -5586 13758 -5552
rect 13792 -5586 13812 -5552
rect 13734 -5614 13812 -5586
rect 10780 -5850 10888 -5774
rect 13730 -5804 13808 -5776
rect 13730 -5838 13757 -5804
rect 13791 -5838 13808 -5804
rect 13730 -5860 13808 -5838
rect 13748 -6196 13788 -5860
rect 13748 -6212 13792 -6196
rect 13750 -11026 13792 -6212
rect 19472 -10888 19532 -20
rect 16320 -10972 19532 -10888
rect 16320 -10974 19466 -10972
rect 13750 -11034 13828 -11026
rect 13750 -11118 13792 -11034
rect 13750 -11126 13818 -11118
rect -90 -24130 -32 -24014
<< viali >>
rect 13754 6541 13788 6575
rect 13759 6156 13793 6190
rect 10805 3984 10839 4018
rect 10787 3278 10821 3312
rect 7374 2264 7408 2298
rect 3883 1223 3917 1257
rect 7388 1416 7422 1450
rect 821 497 855 531
rect 3881 765 3915 799
rect 816 293 850 327
rect 817 -208 851 -174
rect 817 -528 851 -494
rect 3893 -471 3927 -437
rect 3883 -989 3917 -955
rect 7412 -1078 7446 -1044
rect 7414 -1682 7448 -1648
rect 10795 -2228 10829 -2194
rect 10809 -2850 10843 -2816
rect 19559 472 19593 506
rect 13758 -5586 13792 -5552
rect 13757 -5838 13791 -5804
<< metal1 >>
rect 13728 6575 13810 6592
rect 13728 6541 13754 6575
rect 13788 6541 13810 6575
rect 13728 6522 13810 6541
rect 13750 6208 13790 6522
rect 13738 6190 13820 6208
rect 13738 6156 13759 6190
rect 13793 6156 13820 6190
rect 13738 6138 13820 6156
rect 13750 6132 13790 6138
rect 10770 4018 10848 4098
rect 10770 3984 10805 4018
rect 10839 3984 10848 4018
rect 10770 3418 10848 3984
rect 10776 3406 10848 3418
rect 10776 3312 10854 3406
rect 10776 3278 10787 3312
rect 10821 3278 10854 3312
rect 10776 3026 10854 3278
rect 7326 2298 7464 2376
rect 7326 2264 7374 2298
rect 7408 2264 7464 2298
rect 7326 1450 7464 2264
rect 7326 1416 7388 1450
rect 7422 1416 7464 1450
rect 7326 1330 7464 1416
rect 3862 1257 3936 1290
rect 3862 1223 3883 1257
rect 3917 1223 3936 1257
rect 3862 799 3936 1223
rect 3862 765 3881 799
rect 3915 765 3936 799
rect 3862 712 3936 765
rect 18010 827 18118 840
rect 18010 775 18042 827
rect 18094 775 18118 827
rect 18010 760 18118 775
rect 804 531 868 554
rect 804 497 821 531
rect 855 497 868 531
rect 19590 510 19608 518
rect 804 490 868 497
rect 19558 506 19608 510
rect 808 348 866 490
rect 19558 472 19559 506
rect 19593 472 19608 506
rect 19558 468 19608 472
rect 19590 462 19608 468
rect 806 328 866 348
rect 804 327 866 328
rect 804 293 816 327
rect 850 293 866 327
rect 804 290 866 293
rect 804 286 860 290
rect 806 266 860 286
rect 17252 41 17368 102
rect 17252 -11 17281 41
rect 17333 -11 17368 41
rect 17252 -40 17368 -11
rect 804 -174 866 -160
rect 804 -190 817 -174
rect 806 -208 817 -190
rect 851 -190 866 -174
rect 851 -208 864 -190
rect 806 -494 864 -208
rect 806 -528 817 -494
rect 851 -528 864 -494
rect 806 -554 864 -528
rect 3862 -437 3946 -386
rect 3862 -471 3893 -437
rect 3927 -471 3946 -437
rect 3862 -955 3946 -471
rect 3862 -989 3883 -955
rect 3917 -989 3946 -955
rect 3862 -1028 3946 -989
rect 7358 -1044 7496 -950
rect 7358 -1078 7412 -1044
rect 7446 -1078 7496 -1044
rect 7358 -1648 7496 -1078
rect 7358 -1682 7414 -1648
rect 7448 -1682 7496 -1648
rect 7358 -1792 7496 -1682
rect 10772 -2194 10866 -2116
rect 10772 -2228 10795 -2194
rect 10829 -2228 10866 -2194
rect 10772 -2268 10866 -2228
rect 10770 -2658 10866 -2268
rect 10770 -2748 10858 -2658
rect 10770 -2816 10864 -2748
rect 10770 -2850 10809 -2816
rect 10843 -2850 10864 -2816
rect 10770 -2912 10864 -2850
rect 13734 -5552 13812 -5530
rect 13734 -5586 13758 -5552
rect 13792 -5586 13812 -5552
rect 13734 -5614 13812 -5586
rect 13748 -5776 13788 -5614
rect 13730 -5804 13808 -5776
rect 13730 -5838 13757 -5804
rect 13791 -5838 13808 -5804
rect 13730 -5860 13808 -5838
<< via1 >>
rect 18042 775 18094 827
rect 17281 -11 17333 41
<< metal2 >>
rect 13448 5058 16794 5164
rect 16686 50 16786 5058
rect 18028 911 18120 940
rect 18028 902 18050 911
rect 18030 855 18050 902
rect 18106 855 18120 911
rect 18030 827 18120 855
rect 18030 775 18042 827
rect 18094 775 18120 827
rect 18030 760 18120 775
rect 17272 50 17354 52
rect 16686 41 17354 50
rect 16686 0 17281 41
rect 16686 -4344 16786 0
rect 17272 -11 17281 0
rect 17333 -11 17354 41
rect 17272 -28 17354 -11
rect 16680 -6858 16794 -4344
rect 16680 -6972 16808 -6858
rect 16686 -7334 16808 -6972
rect 13370 -7440 16808 -7334
rect 16686 -7468 16808 -7440
<< via2 >>
rect 18050 855 18106 911
<< metal3 >>
rect 18030 1042 18120 1062
rect 18030 978 18045 1042
rect 18109 978 18120 1042
rect 18030 911 18120 978
rect 18030 855 18050 911
rect 18106 855 18120 911
rect 18030 844 18120 855
<< via3 >>
rect 18045 978 18109 1042
<< metal4 >>
rect 17440 7122 18112 7124
rect 16590 7120 18112 7122
rect 15890 7116 18112 7120
rect 15122 7114 18112 7116
rect 13468 7106 18112 7114
rect 12650 7100 18112 7106
rect 11842 7052 18112 7100
rect 11842 7050 16780 7052
rect 11842 7046 16012 7050
rect 11842 7044 15172 7046
rect 11842 7036 13540 7044
rect 11842 7030 12732 7036
rect 18030 3468 18112 7052
rect 18030 3398 18116 3468
rect 18030 2540 18124 3398
rect 18032 2156 18124 2540
rect 17972 2150 18124 2156
rect 14668 2098 18124 2150
rect 14660 2070 18124 2098
rect 14660 -9234 14766 2070
rect 17972 2068 18124 2070
rect 18032 1822 18124 2068
rect 18030 1806 18124 1822
rect 18030 1076 18122 1806
rect 18030 1042 18120 1076
rect 18030 978 18045 1042
rect 18109 978 18120 1042
rect 18030 962 18120 978
rect 14660 -9304 14784 -9234
rect 14668 -10260 14784 -9304
use switch_layout  switch_layout_0
timestamp 1626450099
transform 1 0 17134 0 1 -222
box 40 154 2460 1180
use res250_layout  res250_layout_0
timestamp 1626450099
transform 1 0 -462 0 1 -66
box 202 -342 510 -90
use 5bitdac_layout  5bitdac_layout_0
timestamp 1626450099
transform 1 0 68 0 1 12070
box -70 -12070 16372 11772
use 5bitdac_layout  5bitdac_layout_1
timestamp 1626450099
transform 1 0 -32 0 1 -11978
box -70 -12070 16372 11772
<< labels >>
rlabel locali s 13766 -734 13766 -734 4 d4
port 1 nsew
rlabel locali s 10798 -618 10798 -618 4 d3
port 2 nsew
rlabel locali s 7406 -58 7406 -58 4 d2
port 3 nsew
rlabel locali s 3912 -58 3912 -58 4 d1
port 4 nsew
rlabel locali s 834 58 834 58 4 d0
port 5 nsew
rlabel locali s 322 23712 322 23712 4 inp1
port 6 nsew
rlabel locali s -66 -24090 -66 -24090 4 inp2
port 7 nsew
rlabel locali s 64 -428 64 -428 4 x2_vref1
port 8 nsew
rlabel locali s -160 -152 -160 -152 4 x1_vref5
port 9 nsew
rlabel locali s 19514 -126 19514 -126 4 x2_out_v
port 10 nsew
rlabel locali s 19384 1048 19384 1048 4 x1_out_v
port 11 nsew
rlabel locali s 17138 330 17138 330 4 d5
port 12 nsew
rlabel locali s 19666 494 19666 494 4 out_v
port 13 nsew
rlabel metal2 s 16740 20 16740 20 4 gnd!
port 14 nsew
rlabel metal4 s 18068 1250 18068 1250 4 vdd!
port 15 nsew
<< properties >>
string GDS_FILE gds/adc_wrapper.gds
string GDS_END 56236
string GDS_START 44146
<< end >>
