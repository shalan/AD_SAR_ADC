magic
tech sky130A
magscale 1 2
timestamp 1626641363
<< checkpaint >>
rect -1284 -2558 7762 2690
<< locali >>
rect 400 1308 2254 1310
rect 2630 1308 3014 1310
rect 400 1270 3014 1308
rect 400 1268 2872 1270
rect 400 1066 442 1268
rect 2252 1266 2632 1268
rect 170 738 220 986
rect 400 864 440 1066
rect 2978 1060 3014 1270
rect 150 438 200 538
rect 402 438 440 864
rect 3424 854 3468 856
rect 3424 816 6160 854
rect 3424 790 3468 816
rect 3132 778 3468 790
rect 3132 744 3145 778
rect 3179 744 3468 778
rect 3132 730 3468 744
rect 3132 728 3464 730
rect 778 658 816 662
rect 150 398 440 438
rect 768 410 816 658
rect 6110 576 6160 816
rect 150 290 200 398
rect 672 170 728 184
rect 390 169 728 170
rect 390 135 682 169
rect 716 135 728 169
rect 768 168 818 410
rect 908 176 964 182
rect 2998 176 3056 306
rect 6272 294 6502 306
rect 6272 260 6281 294
rect 6315 260 6502 294
rect 6272 242 6502 260
rect 908 174 3056 176
rect 390 130 728 135
rect 148 0 204 92
rect 390 0 436 130
rect 672 118 728 130
rect 772 128 818 168
rect 904 165 3056 174
rect 904 131 918 165
rect 952 131 3056 165
rect 904 128 3056 131
rect 772 124 816 128
rect 668 6 722 20
rect 668 4 678 6
rect 148 -42 436 0
rect 546 -28 678 4
rect 712 -28 722 6
rect 546 -40 722 -28
rect 148 -340 204 -42
rect 546 -202 590 -40
rect 668 -46 722 -40
rect 770 12 816 124
rect 908 126 3056 128
rect 908 124 3048 126
rect 908 116 964 124
rect 3832 78 4062 180
rect 894 12 952 22
rect 770 -26 818 12
rect 894 8 3044 12
rect 894 -26 904 8
rect 938 -24 3044 8
rect 938 -26 952 -24
rect 1862 -26 2588 -24
rect 770 -120 816 -26
rect 894 -44 952 -26
rect 696 -164 816 -120
rect 192 -342 204 -340
rect 166 -632 260 -542
rect 200 -712 260 -632
rect 544 -708 590 -202
rect 768 -706 816 -164
rect 3004 -222 3044 -24
rect 6156 -482 6196 -172
rect 4644 -486 4882 -484
rect 5080 -486 5318 -484
rect 5524 -486 5762 -484
rect 5960 -486 6198 -482
rect 4202 -488 6198 -486
rect 3524 -492 3762 -490
rect 3980 -492 6198 -488
rect 3156 -509 6198 -492
rect 3156 -543 3170 -509
rect 3204 -538 6198 -509
rect 3204 -540 5988 -538
rect 3204 -542 4662 -540
rect 4864 -542 5102 -540
rect 5294 -542 5532 -540
rect 5750 -542 5988 -540
rect 3204 -543 4218 -542
rect 3156 -544 4218 -543
rect 3156 -546 3990 -544
rect 3156 -548 3534 -546
rect 3752 -548 3990 -546
rect 3156 -550 3300 -548
rect 358 -712 590 -708
rect 776 -712 816 -706
rect 200 -748 590 -712
rect 200 -750 330 -748
rect 200 -908 260 -750
rect -10 -1140 40 -986
rect 1584 -1098 1952 -1096
rect 3034 -1098 3068 -972
rect 332 -1100 380 -1098
rect 548 -1100 3068 -1098
rect 332 -1132 3068 -1100
rect 332 -1134 2634 -1132
rect 330 -1136 1594 -1134
rect 1904 -1136 2634 -1134
rect 330 -1138 704 -1136
rect 330 -1140 380 -1138
rect -10 -1174 380 -1140
rect -10 -1234 40 -1174
<< viali >>
rect 3145 744 3179 778
rect 682 135 716 169
rect 6281 260 6315 294
rect 918 131 952 165
rect 678 -28 712 6
rect 904 -26 938 8
rect 3170 -543 3204 -509
<< metal1 >>
rect 1602 1126 1622 1200
rect 1602 1124 1682 1126
rect 1602 1106 1694 1124
rect 1602 1054 1630 1106
rect 1682 1054 1694 1106
rect 1602 1036 1694 1054
rect 3144 778 3180 780
rect 3144 744 3145 778
rect 3179 744 3180 778
rect 3144 742 3180 744
rect 4742 620 4864 642
rect 4742 568 4789 620
rect 4841 568 4864 620
rect 4742 548 4864 568
rect 906 327 966 374
rect 906 275 909 327
rect 961 275 966 327
rect 906 230 966 275
rect 6280 294 6316 296
rect 6280 260 6281 294
rect 6315 260 6316 294
rect 6280 258 6316 260
rect 672 169 728 184
rect 908 176 964 182
rect 672 168 682 169
rect 670 135 682 168
rect 716 168 728 169
rect 904 168 966 176
rect 716 165 966 168
rect 716 135 918 165
rect 670 131 918 135
rect 952 131 966 165
rect 670 130 966 131
rect 670 128 964 130
rect 672 118 728 128
rect 908 116 964 128
rect 668 12 722 20
rect 894 12 952 22
rect 668 8 952 12
rect 668 6 904 8
rect 668 -28 678 6
rect 712 -26 904 6
rect 938 -26 952 8
rect 712 -28 722 -26
rect 668 -46 722 -28
rect 894 -44 952 -26
rect 1644 -177 1732 -154
rect 1644 -229 1665 -177
rect 1717 -229 1732 -177
rect 1644 -248 1732 -229
rect 4030 -173 4112 -108
rect 4030 -225 4039 -173
rect 4091 -225 4112 -173
rect 4030 -250 4112 -225
rect 4058 -252 4112 -250
rect 3170 -509 3204 -508
rect 3170 -544 3204 -543
rect 942 -955 1002 -904
rect 942 -1007 943 -955
rect 995 -1007 1002 -955
rect 942 -1048 1002 -1007
<< via1 >>
rect 1630 1054 1682 1106
rect 4789 568 4841 620
rect 909 275 961 327
rect 1665 -229 1717 -177
rect 4039 -225 4091 -173
rect 943 -1007 995 -955
<< metal2 >>
rect 1622 1202 1706 1234
rect 1622 1146 1635 1202
rect 1691 1146 1706 1202
rect 1622 1130 1706 1146
rect 1622 1106 1694 1130
rect 1622 1054 1630 1106
rect 1682 1054 1694 1106
rect 1622 1034 1694 1054
rect 4766 721 4866 752
rect 4766 665 4788 721
rect 4844 665 4866 721
rect 4766 620 4866 665
rect 4766 568 4789 620
rect 4841 568 4866 620
rect 4766 548 4866 568
rect 872 327 968 338
rect 872 275 909 327
rect 961 275 968 327
rect 872 258 968 275
rect 872 -936 910 258
rect 1656 -83 1732 -66
rect 1656 -139 1665 -83
rect 1721 -139 1732 -83
rect 1656 -177 1732 -139
rect 4000 -162 4042 -160
rect 3910 -170 4094 -162
rect 1656 -229 1665 -177
rect 1717 -229 1732 -177
rect 1656 -248 1732 -229
rect 3900 -173 4094 -170
rect 3900 -225 4039 -173
rect 4091 -178 4094 -173
rect 4091 -225 4096 -178
rect 3900 -232 4096 -225
rect 3900 -238 4094 -232
rect 3900 -684 3948 -238
rect 4000 -240 4042 -238
rect 3900 -914 3950 -684
rect 872 -942 922 -936
rect 872 -955 1002 -942
rect 872 -1007 943 -955
rect 995 -1007 1002 -955
rect 872 -1022 1002 -1007
rect 874 -1250 922 -1022
rect 3902 -1250 3950 -914
rect 874 -1284 3950 -1250
rect 874 -1298 3896 -1284
<< via2 >>
rect 1635 1146 1691 1202
rect 4788 665 4844 721
rect 1665 -139 1721 -83
<< metal3 >>
rect 1620 1402 1728 1426
rect 1620 1338 1636 1402
rect 1700 1338 1728 1402
rect 1620 1316 1728 1338
rect 1622 1234 1702 1316
rect 1622 1202 1706 1234
rect 1622 1146 1635 1202
rect 1691 1146 1706 1202
rect 1622 1130 1706 1146
rect 1622 1126 1694 1130
rect 4766 940 4868 956
rect 4766 876 4784 940
rect 4848 876 4868 940
rect 4766 858 4868 876
rect 4766 721 4866 858
rect 4766 665 4788 721
rect 4844 665 4866 721
rect 4766 642 4866 665
rect 1656 89 1746 104
rect 1656 25 1668 89
rect 1732 25 1746 89
rect 1656 18 1746 25
rect 1656 -83 1744 18
rect 1656 -139 1665 -83
rect 1721 -139 1744 -83
rect 1656 -154 1744 -139
<< via3 >>
rect 1636 1338 1700 1402
rect 4784 876 4848 940
rect 1668 25 1732 89
<< metal4 >>
rect 2188 1426 4042 1428
rect 4488 1426 4870 1430
rect 1622 1402 4870 1426
rect 1622 1338 1636 1402
rect 1700 1338 4870 1402
rect 1622 1322 4870 1338
rect 1622 1320 4504 1322
rect 1622 1318 2190 1320
rect 4032 1318 4504 1320
rect 1744 102 1854 1318
rect 4766 956 4864 1322
rect 4766 940 4868 956
rect 4766 876 4784 940
rect 4848 876 4868 940
rect 4766 858 4868 876
rect 1656 89 1854 102
rect 1656 25 1668 89
rect 1732 25 1854 89
rect 1656 22 1854 25
rect 1656 18 1772 22
use switch_layout  switch_layout_0
timestamp 1626641363
transform 1 0 732 0 1 50
box 40 154 2460 1180
use switch_layout  switch_layout_1
timestamp 1626641363
transform 1 0 764 0 1 -1230
box 40 154 2460 1180
use switch_layout  switch_layout_2
timestamp 1626641363
transform 1 0 3868 0 1 -434
box 40 154 2460 1180
use res250_layout  res250_layout_0
timestamp 1626641363
transform 0 1 340 -1 0 -598
box 202 -342 510 -90
use res500_layout  res500_layout_0
timestamp 1626641363
transform 0 1 288 -1 0 598
box 202 -312 622 -90
use res500_layout  res500_layout_1
timestamp 1626641363
transform 0 1 288 -1 0 -34
box 202 -312 622 -90
use res500_layout  res500_layout_2
timestamp 1626641363
transform 0 1 296 -1 0 1046
box 202 -312 622 -90
<< labels >>
rlabel locali s 6396 274 6396 274 4 out_v
port 1 nsew
rlabel locali s 3530 -520 3530 -520 4 x2_vout
port 2 nsew
rlabel locali s 3302 754 3302 754 4 x1_vout
port 3 nsew
rlabel locali s 3868 120 3868 120 4 d1
port 4 nsew
rlabel locali s 780 -162 780 -162 4 d0
port 5 nsew
rlabel locali s 6 -1154 6 -1154 4 vref5
port 6 nsew
rlabel locali s 244 -730 244 -730 4 x2_inp1
port 7 nsew
rlabel locali s 160 -128 160 -128 4 x1_inp2
port 8 nsew
rlabel locali s 196 412 196 412 4 x1_inp1
port 9 nsew
rlabel locali s 200 816 200 816 4 vref1
port 10 nsew
rlabel metal2 s 2062 -1274 2062 -1274 4 gnd!
port 11 nsew
<< properties >>
string GDS_FILE gds/adc_wrapper.gds
string GDS_END 23820
string GDS_START 11688
<< end >>
