magic
tech sky130A
magscale 1 2
timestamp 1626101651
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 1104 2128 48852 47376
<< metal2 >>
rect 12438 0 12494 800
rect 37370 0 37426 800
<< obsm2 >>
rect 1398 856 48190 47569
rect 1398 800 12382 856
rect 12550 800 37314 856
rect 37482 800 48190 856
<< metal3 >>
rect 0 47472 800 47592
rect 0 42440 800 42560
rect 49200 41624 50000 41744
rect 0 37408 800 37528
rect 0 32376 800 32496
rect 0 27480 800 27600
rect 49200 24896 50000 25016
rect 0 22448 800 22568
rect 0 17416 800 17536
rect 0 12384 800 12504
rect 49200 8304 50000 8424
rect 0 7352 800 7472
rect 0 2456 800 2576
<< obsm3 >>
rect 880 47392 49200 47565
rect 800 42640 49200 47392
rect 880 42360 49200 42640
rect 800 41824 49200 42360
rect 800 41544 49120 41824
rect 800 37608 49200 41544
rect 880 37328 49200 37608
rect 800 32576 49200 37328
rect 880 32296 49200 32576
rect 800 27680 49200 32296
rect 880 27400 49200 27680
rect 800 25096 49200 27400
rect 800 24816 49120 25096
rect 800 22648 49200 24816
rect 880 22368 49200 22648
rect 800 17616 49200 22368
rect 880 17336 49200 17616
rect 800 12584 49200 17336
rect 880 12304 49200 12584
rect 800 8504 49200 12304
rect 800 8224 49120 8504
rect 800 7552 49200 8224
rect 880 7272 49200 7552
rect 800 2656 49200 7272
rect 880 2376 49200 2656
rect 800 2000 49200 2376
<< metal4 >>
rect 4208 2128 4528 47376
rect 9208 2128 9528 47376
rect 14208 2128 14528 47376
rect 19208 2176 19528 47376
rect 24208 2176 24528 47376
rect 29208 2176 29528 47376
rect 34208 2176 34528 47376
rect 39208 2128 39528 47376
rect 44208 2128 44528 47376
<< labels >>
rlabel metal3 s 49200 24896 50000 25016 6 INN
port 1 nsew signal input
rlabel metal3 s 49200 8304 50000 8424 6 INP
port 2 nsew signal input
rlabel metal3 s 49200 41624 50000 41744 6 Q
port 3 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 clk
port 4 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 data[0]
port 5 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 data[1]
port 6 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 data[2]
port 7 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 data[3]
port 8 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 data[4]
port 9 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 data[5]
port 10 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 data[6]
port 11 nsew signal output
rlabel metal3 s 0 47472 800 47592 6 data[7]
port 12 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 done
port 13 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 rstn
port 14 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 start
port 15 nsew signal input
rlabel metal4 s 44208 2128 44528 47376 6 VPWR
port 16 nsew power bidirectional
rlabel metal4 s 34208 2176 34528 47376 6 VPWR
port 17 nsew power bidirectional
rlabel metal4 s 24208 2176 24528 47376 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 47376 6 VPWR
port 19 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 47376 6 VPWR
port 20 nsew power bidirectional
rlabel metal4 s 39208 2128 39528 47376 6 VGND
port 21 nsew ground bidirectional
rlabel metal4 s 29208 2176 29528 47376 6 VGND
port 22 nsew ground bidirectional
rlabel metal4 s 19208 2176 19528 47376 6 VGND
port 23 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 47376 6 VGND
port 24 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 50000 50000
string LEFview TRUE
string GDS_FILE /project/openlane/adc/runs/adc/results/magic/adc.gds
string GDS_END 1347906
string GDS_START 368056
<< end >>

