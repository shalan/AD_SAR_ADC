magic
tech sky130A
magscale 1 2
timestamp 1626122247
<< obsli1 >>
rect 1104 969 68971 67473
<< obsm1 >>
rect 14 892 69906 67504
<< metal2 >>
rect 938 69200 994 70000
rect 2870 69200 2926 70000
rect 4802 69200 4858 70000
rect 6734 69200 6790 70000
rect 8666 69200 8722 70000
rect 10598 69200 10654 70000
rect 12530 69200 12586 70000
rect 14462 69200 14518 70000
rect 16486 69200 16542 70000
rect 18418 69200 18474 70000
rect 20350 69200 20406 70000
rect 22282 69200 22338 70000
rect 24214 69200 24270 70000
rect 26146 69200 26202 70000
rect 28078 69200 28134 70000
rect 30102 69200 30158 70000
rect 32034 69200 32090 70000
rect 33966 69200 34022 70000
rect 35898 69200 35954 70000
rect 37830 69200 37886 70000
rect 39762 69200 39818 70000
rect 41694 69200 41750 70000
rect 43718 69200 43774 70000
rect 45650 69200 45706 70000
rect 47582 69200 47638 70000
rect 49514 69200 49570 70000
rect 51446 69200 51502 70000
rect 53378 69200 53434 70000
rect 55310 69200 55366 70000
rect 57334 69200 57390 70000
rect 59266 69200 59322 70000
rect 61198 69200 61254 70000
rect 63130 69200 63186 70000
rect 65062 69200 65118 70000
rect 66994 69200 67050 70000
rect 68926 69200 68982 70000
rect 18 0 74 800
rect 110 0 166 800
rect 294 0 350 800
rect 386 0 442 800
rect 570 0 626 800
rect 662 0 718 800
rect 846 0 902 800
rect 938 0 994 800
rect 1122 0 1178 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 1950 0 2006 800
rect 2134 0 2190 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68098 0 68154 800
rect 68282 0 68338 800
rect 68466 0 68522 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69662 0 69718 800
rect 69846 0 69902 800
<< obsm2 >>
rect 20 69144 882 69329
rect 1050 69144 2814 69329
rect 2982 69144 4746 69329
rect 4914 69144 6678 69329
rect 6846 69144 8610 69329
rect 8778 69144 10542 69329
rect 10710 69144 12474 69329
rect 12642 69144 14406 69329
rect 14574 69144 16430 69329
rect 16598 69144 18362 69329
rect 18530 69144 20294 69329
rect 20462 69144 22226 69329
rect 22394 69144 24158 69329
rect 24326 69144 26090 69329
rect 26258 69144 28022 69329
rect 28190 69144 30046 69329
rect 30214 69144 31978 69329
rect 32146 69144 33910 69329
rect 34078 69144 35842 69329
rect 36010 69144 37774 69329
rect 37942 69144 39706 69329
rect 39874 69144 41638 69329
rect 41806 69144 43662 69329
rect 43830 69144 45594 69329
rect 45762 69144 47526 69329
rect 47694 69144 49458 69329
rect 49626 69144 51390 69329
rect 51558 69144 53322 69329
rect 53490 69144 55254 69329
rect 55422 69144 57278 69329
rect 57446 69144 59210 69329
rect 59378 69144 61142 69329
rect 61310 69144 63074 69329
rect 63242 69144 65006 69329
rect 65174 69144 66938 69329
rect 67106 69144 68870 69329
rect 69038 69144 69900 69329
rect 20 856 69900 69144
rect 222 575 238 856
rect 498 575 514 856
rect 774 575 790 856
rect 1050 575 1066 856
rect 1326 575 1342 856
rect 1602 575 1618 856
rect 1786 575 1802 856
rect 2062 575 2078 856
rect 2338 575 2354 856
rect 2614 575 2630 856
rect 2890 575 2906 856
rect 3166 575 3182 856
rect 3442 575 3458 856
rect 3626 575 3642 856
rect 3902 575 3918 856
rect 4178 575 4194 856
rect 4454 575 4470 856
rect 4730 575 4746 856
rect 5006 575 5022 856
rect 5282 575 5298 856
rect 5466 575 5482 856
rect 5742 575 5758 856
rect 6018 575 6034 856
rect 6294 575 6310 856
rect 6570 575 6586 856
rect 6846 575 6862 856
rect 7030 575 7046 856
rect 7306 575 7322 856
rect 7582 575 7598 856
rect 7858 575 7874 856
rect 8134 575 8150 856
rect 8410 575 8426 856
rect 8686 575 8702 856
rect 8870 575 8886 856
rect 9146 575 9162 856
rect 9422 575 9438 856
rect 9698 575 9714 856
rect 9974 575 9990 856
rect 10250 575 10266 856
rect 10526 575 10542 856
rect 10710 575 10726 856
rect 10986 575 11002 856
rect 11262 575 11278 856
rect 11538 575 11554 856
rect 11814 575 11830 856
rect 12090 575 12106 856
rect 12274 575 12290 856
rect 12550 575 12566 856
rect 12826 575 12842 856
rect 13102 575 13118 856
rect 13378 575 13394 856
rect 13654 575 13670 856
rect 13930 575 13946 856
rect 14114 575 14130 856
rect 14390 575 14406 856
rect 14666 575 14682 856
rect 14942 575 14958 856
rect 15218 575 15234 856
rect 15494 575 15510 856
rect 15770 575 15786 856
rect 15954 575 15970 856
rect 16230 575 16246 856
rect 16506 575 16522 856
rect 16782 575 16798 856
rect 17058 575 17074 856
rect 17334 575 17350 856
rect 17518 575 17534 856
rect 17794 575 17810 856
rect 18070 575 18086 856
rect 18346 575 18362 856
rect 18622 575 18638 856
rect 18898 575 18914 856
rect 19174 575 19190 856
rect 19358 575 19374 856
rect 19634 575 19650 856
rect 19910 575 19926 856
rect 20186 575 20202 856
rect 20462 575 20478 856
rect 20738 575 20754 856
rect 21014 575 21030 856
rect 21198 575 21214 856
rect 21474 575 21490 856
rect 21750 575 21766 856
rect 22026 575 22042 856
rect 22302 575 22318 856
rect 22578 575 22594 856
rect 22762 575 22778 856
rect 23038 575 23054 856
rect 23314 575 23330 856
rect 23590 575 23606 856
rect 23866 575 23882 856
rect 24142 575 24158 856
rect 24418 575 24434 856
rect 24602 575 24618 856
rect 24878 575 24894 856
rect 25154 575 25170 856
rect 25430 575 25446 856
rect 25706 575 25722 856
rect 25982 575 25998 856
rect 26258 575 26274 856
rect 26442 575 26458 856
rect 26718 575 26734 856
rect 26994 575 27010 856
rect 27270 575 27286 856
rect 27546 575 27562 856
rect 27822 575 27838 856
rect 28006 575 28022 856
rect 28282 575 28298 856
rect 28558 575 28574 856
rect 28834 575 28850 856
rect 29110 575 29126 856
rect 29386 575 29402 856
rect 29662 575 29678 856
rect 29846 575 29862 856
rect 30122 575 30138 856
rect 30398 575 30414 856
rect 30674 575 30690 856
rect 30950 575 30966 856
rect 31226 575 31242 856
rect 31502 575 31518 856
rect 31686 575 31702 856
rect 31962 575 31978 856
rect 32238 575 32254 856
rect 32514 575 32530 856
rect 32790 575 32806 856
rect 33066 575 33082 856
rect 33250 575 33266 856
rect 33526 575 33542 856
rect 33802 575 33818 856
rect 34078 575 34094 856
rect 34354 575 34370 856
rect 34630 575 34646 856
rect 34906 575 34922 856
rect 35090 575 35106 856
rect 35366 575 35382 856
rect 35642 575 35658 856
rect 35918 575 35934 856
rect 36194 575 36210 856
rect 36470 575 36486 856
rect 36746 575 36762 856
rect 36930 575 36946 856
rect 37206 575 37222 856
rect 37482 575 37498 856
rect 37758 575 37774 856
rect 38034 575 38050 856
rect 38310 575 38326 856
rect 38494 575 38510 856
rect 38770 575 38786 856
rect 39046 575 39062 856
rect 39322 575 39338 856
rect 39598 575 39614 856
rect 39874 575 39890 856
rect 40150 575 40166 856
rect 40334 575 40350 856
rect 40610 575 40626 856
rect 40886 575 40902 856
rect 41162 575 41178 856
rect 41438 575 41454 856
rect 41714 575 41730 856
rect 41990 575 42006 856
rect 42174 575 42190 856
rect 42450 575 42466 856
rect 42726 575 42742 856
rect 43002 575 43018 856
rect 43278 575 43294 856
rect 43554 575 43570 856
rect 43738 575 43754 856
rect 44014 575 44030 856
rect 44290 575 44306 856
rect 44566 575 44582 856
rect 44842 575 44858 856
rect 45118 575 45134 856
rect 45394 575 45410 856
rect 45578 575 45594 856
rect 45854 575 45870 856
rect 46130 575 46146 856
rect 46406 575 46422 856
rect 46682 575 46698 856
rect 46958 575 46974 856
rect 47234 575 47250 856
rect 47418 575 47434 856
rect 47694 575 47710 856
rect 47970 575 47986 856
rect 48246 575 48262 856
rect 48522 575 48538 856
rect 48798 575 48814 856
rect 48982 575 48998 856
rect 49258 575 49274 856
rect 49534 575 49550 856
rect 49810 575 49826 856
rect 50086 575 50102 856
rect 50362 575 50378 856
rect 50638 575 50654 856
rect 50822 575 50838 856
rect 51098 575 51114 856
rect 51374 575 51390 856
rect 51650 575 51666 856
rect 51926 575 51942 856
rect 52202 575 52218 856
rect 52478 575 52494 856
rect 52662 575 52678 856
rect 52938 575 52954 856
rect 53214 575 53230 856
rect 53490 575 53506 856
rect 53766 575 53782 856
rect 54042 575 54058 856
rect 54226 575 54242 856
rect 54502 575 54518 856
rect 54778 575 54794 856
rect 55054 575 55070 856
rect 55330 575 55346 856
rect 55606 575 55622 856
rect 55882 575 55898 856
rect 56066 575 56082 856
rect 56342 575 56358 856
rect 56618 575 56634 856
rect 56894 575 56910 856
rect 57170 575 57186 856
rect 57446 575 57462 856
rect 57722 575 57738 856
rect 57906 575 57922 856
rect 58182 575 58198 856
rect 58458 575 58474 856
rect 58734 575 58750 856
rect 59010 575 59026 856
rect 59286 575 59302 856
rect 59470 575 59486 856
rect 59746 575 59762 856
rect 60022 575 60038 856
rect 60298 575 60314 856
rect 60574 575 60590 856
rect 60850 575 60866 856
rect 61126 575 61142 856
rect 61310 575 61326 856
rect 61586 575 61602 856
rect 61862 575 61878 856
rect 62138 575 62154 856
rect 62414 575 62430 856
rect 62690 575 62706 856
rect 62966 575 62982 856
rect 63150 575 63166 856
rect 63426 575 63442 856
rect 63702 575 63718 856
rect 63978 575 63994 856
rect 64254 575 64270 856
rect 64530 575 64546 856
rect 64714 575 64730 856
rect 64990 575 65006 856
rect 65266 575 65282 856
rect 65542 575 65558 856
rect 65818 575 65834 856
rect 66094 575 66110 856
rect 66370 575 66386 856
rect 66554 575 66570 856
rect 66830 575 66846 856
rect 67106 575 67122 856
rect 67382 575 67398 856
rect 67658 575 67674 856
rect 67934 575 67950 856
rect 68210 575 68226 856
rect 68394 575 68410 856
rect 68670 575 68686 856
rect 68946 575 68962 856
rect 69222 575 69238 856
rect 69498 575 69514 856
rect 69774 575 69790 856
<< metal3 >>
rect 0 69232 800 69352
rect 69200 69232 70000 69352
rect 0 67872 800 67992
rect 69200 67872 70000 67992
rect 0 66648 800 66768
rect 69200 66512 70000 66632
rect 0 65288 800 65408
rect 69200 65288 70000 65408
rect 0 64064 800 64184
rect 69200 63928 70000 64048
rect 0 62704 800 62824
rect 69200 62568 70000 62688
rect 0 61480 800 61600
rect 69200 61208 70000 61328
rect 0 60120 800 60240
rect 69200 59984 70000 60104
rect 0 58896 800 59016
rect 69200 58624 70000 58744
rect 0 57536 800 57656
rect 69200 57264 70000 57384
rect 0 56312 800 56432
rect 69200 56040 70000 56160
rect 0 54952 800 55072
rect 69200 54680 70000 54800
rect 0 53728 800 53848
rect 69200 53320 70000 53440
rect 0 52368 800 52488
rect 69200 51960 70000 52080
rect 0 51008 800 51128
rect 69200 50736 70000 50856
rect 0 49784 800 49904
rect 69200 49376 70000 49496
rect 0 48424 800 48544
rect 69200 48016 70000 48136
rect 0 47200 800 47320
rect 69200 46792 70000 46912
rect 0 45840 800 45960
rect 69200 45432 70000 45552
rect 0 44616 800 44736
rect 69200 44072 70000 44192
rect 0 43256 800 43376
rect 69200 42712 70000 42832
rect 0 42032 800 42152
rect 69200 41488 70000 41608
rect 0 40672 800 40792
rect 69200 40128 70000 40248
rect 0 39448 800 39568
rect 69200 38768 70000 38888
rect 0 38088 800 38208
rect 69200 37544 70000 37664
rect 0 36864 800 36984
rect 69200 36184 70000 36304
rect 0 35504 800 35624
rect 69200 34824 70000 34944
rect 0 34144 800 34264
rect 69200 33464 70000 33584
rect 0 32920 800 33040
rect 69200 32240 70000 32360
rect 0 31560 800 31680
rect 69200 30880 70000 31000
rect 0 30336 800 30456
rect 69200 29520 70000 29640
rect 0 28976 800 29096
rect 69200 28296 70000 28416
rect 0 27752 800 27872
rect 69200 26936 70000 27056
rect 0 26392 800 26512
rect 69200 25576 70000 25696
rect 0 25168 800 25288
rect 69200 24216 70000 24336
rect 0 23808 800 23928
rect 69200 22992 70000 23112
rect 0 22584 800 22704
rect 69200 21632 70000 21752
rect 0 21224 800 21344
rect 69200 20272 70000 20392
rect 0 20000 800 20120
rect 69200 19048 70000 19168
rect 0 18640 800 18760
rect 69200 17688 70000 17808
rect 0 17280 800 17400
rect 69200 16328 70000 16448
rect 0 16056 800 16176
rect 69200 14968 70000 15088
rect 0 14696 800 14816
rect 69200 13744 70000 13864
rect 0 13472 800 13592
rect 69200 12384 70000 12504
rect 0 12112 800 12232
rect 0 10888 800 11008
rect 69200 11024 70000 11144
rect 69200 9800 70000 9920
rect 0 9528 800 9648
rect 0 8304 800 8424
rect 69200 8440 70000 8560
rect 0 6944 800 7064
rect 69200 7080 70000 7200
rect 0 5720 800 5840
rect 69200 5720 70000 5840
rect 0 4360 800 4480
rect 69200 4496 70000 4616
rect 0 3136 800 3256
rect 69200 3136 70000 3256
rect 0 1776 800 1896
rect 69200 1776 70000 1896
rect 0 552 800 672
rect 69200 552 70000 672
<< obsm3 >>
rect 880 69152 69120 69325
rect 800 68072 69200 69152
rect 880 67792 69120 68072
rect 800 66848 69200 67792
rect 880 66712 69200 66848
rect 880 66568 69120 66712
rect 800 66432 69120 66568
rect 800 65488 69200 66432
rect 880 65208 69120 65488
rect 800 64264 69200 65208
rect 880 64128 69200 64264
rect 880 63984 69120 64128
rect 800 63848 69120 63984
rect 800 62904 69200 63848
rect 880 62768 69200 62904
rect 880 62624 69120 62768
rect 800 62488 69120 62624
rect 800 61680 69200 62488
rect 880 61408 69200 61680
rect 880 61400 69120 61408
rect 800 61128 69120 61400
rect 800 60320 69200 61128
rect 880 60184 69200 60320
rect 880 60040 69120 60184
rect 800 59904 69120 60040
rect 800 59096 69200 59904
rect 880 58824 69200 59096
rect 880 58816 69120 58824
rect 800 58544 69120 58816
rect 800 57736 69200 58544
rect 880 57464 69200 57736
rect 880 57456 69120 57464
rect 800 57184 69120 57456
rect 800 56512 69200 57184
rect 880 56240 69200 56512
rect 880 56232 69120 56240
rect 800 55960 69120 56232
rect 800 55152 69200 55960
rect 880 54880 69200 55152
rect 880 54872 69120 54880
rect 800 54600 69120 54872
rect 800 53928 69200 54600
rect 880 53648 69200 53928
rect 800 53520 69200 53648
rect 800 53240 69120 53520
rect 800 52568 69200 53240
rect 880 52288 69200 52568
rect 800 52160 69200 52288
rect 800 51880 69120 52160
rect 800 51208 69200 51880
rect 880 50936 69200 51208
rect 880 50928 69120 50936
rect 800 50656 69120 50928
rect 800 49984 69200 50656
rect 880 49704 69200 49984
rect 800 49576 69200 49704
rect 800 49296 69120 49576
rect 800 48624 69200 49296
rect 880 48344 69200 48624
rect 800 48216 69200 48344
rect 800 47936 69120 48216
rect 800 47400 69200 47936
rect 880 47120 69200 47400
rect 800 46992 69200 47120
rect 800 46712 69120 46992
rect 800 46040 69200 46712
rect 880 45760 69200 46040
rect 800 45632 69200 45760
rect 800 45352 69120 45632
rect 800 44816 69200 45352
rect 880 44536 69200 44816
rect 800 44272 69200 44536
rect 800 43992 69120 44272
rect 800 43456 69200 43992
rect 880 43176 69200 43456
rect 800 42912 69200 43176
rect 800 42632 69120 42912
rect 800 42232 69200 42632
rect 880 41952 69200 42232
rect 800 41688 69200 41952
rect 800 41408 69120 41688
rect 800 40872 69200 41408
rect 880 40592 69200 40872
rect 800 40328 69200 40592
rect 800 40048 69120 40328
rect 800 39648 69200 40048
rect 880 39368 69200 39648
rect 800 38968 69200 39368
rect 800 38688 69120 38968
rect 800 38288 69200 38688
rect 880 38008 69200 38288
rect 800 37744 69200 38008
rect 800 37464 69120 37744
rect 800 37064 69200 37464
rect 880 36784 69200 37064
rect 800 36384 69200 36784
rect 800 36104 69120 36384
rect 800 35704 69200 36104
rect 880 35424 69200 35704
rect 800 35024 69200 35424
rect 800 34744 69120 35024
rect 800 34344 69200 34744
rect 880 34064 69200 34344
rect 800 33664 69200 34064
rect 800 33384 69120 33664
rect 800 33120 69200 33384
rect 880 32840 69200 33120
rect 800 32440 69200 32840
rect 800 32160 69120 32440
rect 800 31760 69200 32160
rect 880 31480 69200 31760
rect 800 31080 69200 31480
rect 800 30800 69120 31080
rect 800 30536 69200 30800
rect 880 30256 69200 30536
rect 800 29720 69200 30256
rect 800 29440 69120 29720
rect 800 29176 69200 29440
rect 880 28896 69200 29176
rect 800 28496 69200 28896
rect 800 28216 69120 28496
rect 800 27952 69200 28216
rect 880 27672 69200 27952
rect 800 27136 69200 27672
rect 800 26856 69120 27136
rect 800 26592 69200 26856
rect 880 26312 69200 26592
rect 800 25776 69200 26312
rect 800 25496 69120 25776
rect 800 25368 69200 25496
rect 880 25088 69200 25368
rect 800 24416 69200 25088
rect 800 24136 69120 24416
rect 800 24008 69200 24136
rect 880 23728 69200 24008
rect 800 23192 69200 23728
rect 800 22912 69120 23192
rect 800 22784 69200 22912
rect 880 22504 69200 22784
rect 800 21832 69200 22504
rect 800 21552 69120 21832
rect 800 21424 69200 21552
rect 880 21144 69200 21424
rect 800 20472 69200 21144
rect 800 20200 69120 20472
rect 880 20192 69120 20200
rect 880 19920 69200 20192
rect 800 19248 69200 19920
rect 800 18968 69120 19248
rect 800 18840 69200 18968
rect 880 18560 69200 18840
rect 800 17888 69200 18560
rect 800 17608 69120 17888
rect 800 17480 69200 17608
rect 880 17200 69200 17480
rect 800 16528 69200 17200
rect 800 16256 69120 16528
rect 880 16248 69120 16256
rect 880 15976 69200 16248
rect 800 15168 69200 15976
rect 800 14896 69120 15168
rect 880 14888 69120 14896
rect 880 14616 69200 14888
rect 800 13944 69200 14616
rect 800 13672 69120 13944
rect 880 13664 69120 13672
rect 880 13392 69200 13664
rect 800 12584 69200 13392
rect 800 12312 69120 12584
rect 880 12304 69120 12312
rect 880 12032 69200 12304
rect 800 11224 69200 12032
rect 800 11088 69120 11224
rect 880 10944 69120 11088
rect 880 10808 69200 10944
rect 800 10000 69200 10808
rect 800 9728 69120 10000
rect 880 9720 69120 9728
rect 880 9448 69200 9720
rect 800 8640 69200 9448
rect 800 8504 69120 8640
rect 880 8360 69120 8504
rect 880 8224 69200 8360
rect 800 7280 69200 8224
rect 800 7144 69120 7280
rect 880 7000 69120 7144
rect 880 6864 69200 7000
rect 800 5920 69200 6864
rect 880 5640 69120 5920
rect 800 4696 69200 5640
rect 800 4560 69120 4696
rect 880 4416 69120 4560
rect 880 4280 69200 4416
rect 800 3336 69200 4280
rect 880 3056 69120 3336
rect 800 1976 69200 3056
rect 880 1696 69120 1976
rect 800 752 69200 1696
rect 880 579 69120 752
<< metal4 >>
rect 4208 2128 4528 67504
rect 9208 2128 9528 67504
rect 14208 2128 14528 67504
rect 19208 2176 19528 67504
rect 24208 2176 24528 67504
rect 29208 2176 29528 67504
rect 34208 2176 34528 67504
rect 39208 2128 39528 67504
rect 44208 2128 44528 67504
rect 49208 2128 49528 67504
rect 54208 2128 54528 67504
rect 59208 2128 59528 67504
rect 64208 2128 64528 67504
<< obsm4 >>
rect 5395 2048 9128 32469
rect 9608 2048 14128 32469
rect 14608 2096 19128 32469
rect 19608 2096 24128 32469
rect 24608 2096 29128 32469
rect 29608 2096 34128 32469
rect 34608 2096 39128 32469
rect 14608 2048 39128 2096
rect 39608 2048 44128 32469
rect 44608 2048 49128 32469
rect 49608 2048 54128 32469
rect 54608 2048 59128 32469
rect 59608 2048 64128 32469
rect 64608 2048 64709 32469
rect 5395 1123 64709 2048
<< labels >>
rlabel metal3 s 69200 28296 70000 28416 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 53378 69200 53434 70000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 45650 69200 45706 70000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 37830 69200 37886 70000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 30102 69200 30158 70000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 22282 69200 22338 70000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 14462 69200 14518 70000 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 6734 69200 6790 70000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 69232 800 69352 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 64064 800 64184 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 58896 800 59016 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 69200 33464 70000 33584 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 53728 800 53848 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 48424 800 48544 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 43256 800 43376 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 38088 800 38208 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 32920 800 33040 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 27752 800 27872 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 22584 800 22704 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 17280 800 17400 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 12112 800 12232 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 69200 38768 70000 38888 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 69200 44072 70000 44192 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 69200 49376 70000 49496 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 69200 54680 70000 54800 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 69200 59984 70000 60104 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 69200 65288 70000 65408 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 68926 69200 68982 70000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 61198 69200 61254 70000 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 69200 552 70000 672 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 69200 45432 70000 45552 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 69200 50736 70000 50856 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 69200 56040 70000 56160 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 69200 61208 70000 61328 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 69200 66512 70000 66632 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 66994 69200 67050 70000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 59266 69200 59322 70000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 51446 69200 51502 70000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 43718 69200 43774 70000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 35898 69200 35954 70000 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 69200 4496 70000 4616 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 28078 69200 28134 70000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 20350 69200 20406 70000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 12530 69200 12586 70000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 4802 69200 4858 70000 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 69200 8440 70000 8560 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 69200 12384 70000 12504 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 69200 16328 70000 16448 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 69200 20272 70000 20392 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 69200 24216 70000 24336 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 69200 29520 70000 29640 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 69200 34824 70000 34944 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 69200 40128 70000 40248 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 69200 3136 70000 3256 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 69200 48016 70000 48136 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 69200 53320 70000 53440 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 69200 58624 70000 58744 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 69200 63928 70000 64048 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 69200 69232 70000 69352 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 63130 69200 63186 70000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 55310 69200 55366 70000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 47582 69200 47638 70000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 39762 69200 39818 70000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 32034 69200 32090 70000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 69200 7080 70000 7200 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 24214 69200 24270 70000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 16486 69200 16542 70000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 8666 69200 8722 70000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 938 69200 994 70000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 69200 11024 70000 11144 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 28976 800 29096 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 552 800 672 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 69200 14968 70000 15088 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 69200 19048 70000 19168 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 69200 22992 70000 23112 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 69200 26936 70000 27056 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 69200 32240 70000 32360 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 69200 37544 70000 37664 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 69200 42712 70000 42832 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 69200 1776 70000 1896 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 69200 46792 70000 46912 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 69200 51960 70000 52080 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 69200 57264 70000 57384 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 69200 62568 70000 62688 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 69200 67872 70000 67992 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 65062 69200 65118 70000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 57334 69200 57390 70000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 49514 69200 49570 70000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 41694 69200 41750 70000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 33966 69200 34022 70000 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 69200 5720 70000 5840 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 26146 69200 26202 70000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 18418 69200 18474 70000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 10598 69200 10654 70000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 2870 69200 2926 70000 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 69200 9800 70000 9920 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 35504 800 35624 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 69200 13744 70000 13864 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 69200 17688 70000 17808 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 69200 21632 70000 21752 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 69200 25576 70000 25696 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 69200 30880 70000 31000 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 69200 36184 70000 36304 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 69200 41488 70000 41608 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 532 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 294 0 350 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 846 0 902 800 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 386 0 442 800 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 64208 2128 64528 67504 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 67504 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 67504 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 34208 2176 34528 67504 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 24208 2176 24528 67504 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 67504 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 67504 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 59208 2128 59528 67504 6 VGND
port 645 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 67504 6 VGND
port 646 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 67504 6 VGND
port 647 nsew ground bidirectional
rlabel metal4 s 29208 2176 29528 67504 6 VGND
port 648 nsew ground bidirectional
rlabel metal4 s 19208 2176 19528 67504 6 VGND
port 649 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 67504 6 VGND
port 650 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 70000 70000
string LEFview TRUE
string GDS_FILE /project/openlane/adc_wrapper/runs/adc_wrapper/results/magic/adc_wrapper.gds
string GDS_END 4002228
string GDS_START 446762
<< end >>

